* NGSPICE file created from cordic_system.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

.subckt cordic_system VGND VPWR aclk araddr[0] araddr[10] araddr[11] araddr[12] araddr[13]
+ araddr[14] araddr[15] araddr[16] araddr[17] araddr[18] araddr[19] araddr[1] araddr[20]
+ araddr[21] araddr[22] araddr[23] araddr[24] araddr[25] araddr[26] araddr[27] araddr[28]
+ araddr[29] araddr[2] araddr[30] araddr[31] araddr[3] araddr[4] araddr[5] araddr[6]
+ araddr[7] araddr[8] araddr[9] aresetn arready arvalid awaddr[0] awaddr[10] awaddr[11]
+ awaddr[12] awaddr[13] awaddr[14] awaddr[15] awaddr[16] awaddr[17] awaddr[18] awaddr[19]
+ awaddr[1] awaddr[20] awaddr[21] awaddr[22] awaddr[23] awaddr[24] awaddr[25] awaddr[26]
+ awaddr[27] awaddr[28] awaddr[29] awaddr[2] awaddr[30] awaddr[31] awaddr[3] awaddr[4]
+ awaddr[5] awaddr[6] awaddr[7] awaddr[8] awaddr[9] awready awvalid bready bresp[0]
+ bresp[1] bvalid rdata[0] rdata[10] rdata[11] rdata[12] rdata[13] rdata[14] rdata[15]
+ rdata[16] rdata[17] rdata[18] rdata[19] rdata[1] rdata[20] rdata[21] rdata[22] rdata[23]
+ rdata[24] rdata[25] rdata[26] rdata[27] rdata[28] rdata[29] rdata[2] rdata[30] rdata[31]
+ rdata[3] rdata[4] rdata[5] rdata[6] rdata[7] rdata[8] rdata[9] rready rresp[0] rresp[1]
+ rvalid wdata[0] wdata[10] wdata[11] wdata[12] wdata[13] wdata[14] wdata[15] wdata[16]
+ wdata[17] wdata[18] wdata[19] wdata[1] wdata[20] wdata[21] wdata[22] wdata[23] wdata[24]
+ wdata[25] wdata[26] wdata[27] wdata[28] wdata[29] wdata[2] wdata[30] wdata[31] wdata[3]
+ wdata[4] wdata[5] wdata[6] wdata[7] wdata[8] wdata[9] wready wstrb[0] wstrb[1] wstrb[2]
+ wstrb[3] wvalid
XFILLER_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3155_ _1318_ _1441_ _1329_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__o21a_1
X_3086_ _1387_ _1388_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__and2_1
XFILLER_54_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3988_ _1939_ _1941_ _1997_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__or3_1
X_2939_ _1103_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_20_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4609_ net377 _0341_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4960_ net411 _0589_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_1
X_3911_ axi_controller.read_addr_reg\[12\] net5 net195 VGND VGND VPWR VPWR _0278_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4891_ net378 _0044_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3842_ net145 net70 net194 VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__a21oi_1
X_3773_ axi_controller.reg_input_data\[30\] axi_controller.reg_input_data\[29\] _1877_
+ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__nand3_1
XFILLER_8_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2724_ _0925_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__or2_1
X_2655_ cordic_inst.cordic_inst.y\[25\] _0988_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nand2_1
X_4325_ net121 net192 net155 axi_controller.result_out\[18\] VGND VGND VPWR VPWR _0576_
+ sky130_fd_sc_hd__a22o_1
X_2586_ net252 _0770_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__nor2_1
XFILLER_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4256_ net316 _2214_ _2215_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__and3_1
Xfanout149 net150 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3207_ cordic_inst.cordic_inst.y\[26\] cordic_inst.cordic_inst.sin_out\[26\] net207
+ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
X_4187_ cordic_inst.cordic_inst.cos_out\[18\] _2147_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__or2_1
X_3138_ net180 _1421_ _1429_ net160 cordic_inst.cordic_inst.x\[20\] VGND VGND VPWR
+ VPWR _0518_ sky130_fd_sc_hd__a32o_1
XFILLER_67_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3069_ cordic_inst.cordic_inst.x\[23\] _1334_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_53_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2440_ _0719_ _0722_ _0727_ _0720_ net283 net233 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__mux4_1
X_2371_ net242 net314 VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__nand2_1
X_4110_ cordic_inst.cordic_inst.sin_out\[10\] net261 _2086_ VGND VGND VPWR VPWR _2087_
+ sky130_fd_sc_hd__and3_1
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4041_ cordic_inst.cordic_inst.cos_out\[0\] cordic_inst.cordic_inst.sin_out\[0\]
+ net319 VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4943_ net368 _0572_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4874_ net388 axi_controller.reg_input_data\[6\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3825_ cordic_inst.cordic_inst.start cordic_inst.cordic_inst.state\[1\] cordic_inst.cordic_inst.state\[0\]
+ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__o21ba_1
X_3756_ cordic_inst.deg_handler_inst.theta_norm\[29\] cordic_inst.deg_handler_inst.theta_norm\[28\]
+ _1859_ net253 VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__o31a_1
X_2707_ _0854_ _0858_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_30_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3687_ net256 _1819_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__nand2_1
X_2638_ _0869_ _0968_ _0970_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__or3_1
X_2569_ _0889_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nor2_1
X_4308_ axi_controller.state\[0\] axi_controller.state\[1\] _0621_ net144 VGND VGND
+ VPWR VPWR _2255_ sky130_fd_sc_hd__or4b_1
X_4239_ cordic_inst.cordic_inst.sin_out\[25\] net257 _2199_ net228 VGND VGND VPWR
+ VPWR _2201_ sky130_fd_sc_hd__a31o_1
XFILLER_74_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_85_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4590_ net360 _0322_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[23\] sky130_fd_sc_hd__dfxtp_1
X_3610_ cordic_inst.deg_handler_inst.theta_abs\[24\] cordic_inst.deg_handler_inst.theta_abs\[25\]
+ cordic_inst.deg_handler_inst.theta_abs\[26\] cordic_inst.deg_handler_inst.theta_abs\[27\]
+ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__or4_1
X_3541_ net183 _1601_ _1749_ _1750_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a31o_1
X_3472_ cordic_inst.cordic_inst.angle\[21\] net170 net164 cordic_inst.cordic_inst.z\[21\]
+ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__a22o_1
X_2423_ _0684_ _0693_ _0750_ _0756_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__and4_1
XFILLER_69_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2354_ net286 _0685_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__a21o_1
XFILLER_84_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2285_ net350 VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__inv_2
X_4024_ net103 _1963_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__nand2_2
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4926_ net373 _0026_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_4857_ net386 _0066_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[21\] sky130_fd_sc_hd__dfxtp_1
X_3808_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1900_
+ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__and3_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4788_ net397 _0515_ _0210_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[17\] sky130_fd_sc_hd__dfrtp_4
X_3739_ cordic_inst.deg_handler_inst.theta_norm\[23\] cordic_inst.deg_handler_inst.theta_norm\[22\]
+ _1849_ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_7_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2972_ cordic_inst.cordic_inst.x\[3\] _1262_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__or2_1
X_4711_ net403 _0438_ _0133_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_61_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4642_ net394 _0373_ net329 VGND VGND VPWR VPWR axi_controller.result_out\[19\] sky130_fd_sc_hd__dfrtp_1
X_4573_ net370 _0305_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_3524_ net176 _1610_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__or2_1
XFILLER_89_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3455_ _1686_ _1687_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__nor2_1
X_2406_ _0679_ net219 _0739_ net286 VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__a22o_1
X_3386_ _1540_ _1546_ _1621_ _1624_ _1539_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_4_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2337_ net280 _0670_ _0671_ _0631_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o31a_1
X_2268_ cordic_inst.cordic_inst.cos_out\[26\] VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__inv_2
X_4007_ axi_controller.reg_input_data\[24\] _2008_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__or2_1
XFILLER_72_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4909_ net390 _0039_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3240_ net249 cordic_inst.cordic_inst.z\[24\] VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__or2_1
X_3171_ net175 _1452_ _1453_ cordic_inst.cordic_inst.next_state\[1\] cordic_inst.cordic_inst.x\[11\]
+ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__o32a_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2955_ _1257_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__inv_2
X_2886_ _1180_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__or2_1
X_4625_ net412 _0356_ net347 VGND VGND VPWR VPWR axi_controller.result_out\[2\] sky130_fd_sc_hd__dfrtp_1
X_4556_ net359 _0288_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[22\] sky130_fd_sc_hd__dfxtp_1
X_3507_ _1535_ _1625_ _1626_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__and3_1
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4487_ net345 VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__inv_2
X_3438_ _1475_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__xnor2_1
X_3369_ _1568_ _1606_ _1563_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__o21ba_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2740_ cordic_inst.cordic_inst.y\[10\] net161 _1052_ _1053_ VGND VGND VPWR VPWR _0540_
+ sky130_fd_sc_hd__a22o_1
X_2671_ _1004_ _1005_ net264 net158 VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4410_ net339 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__inv_2
X_4341_ net134 net193 net154 axi_controller.result_out\[2\] VGND VGND VPWR VPWR _0592_
+ sky130_fd_sc_hd__a22o_1
X_4272_ axi_controller.result_out\[29\] _2229_ net199 VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__mux2_1
Xfanout309 net310 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_4
X_3223_ cordic_inst.cordic_inst.y\[10\] cordic_inst.cordic_inst.sin_out\[10\] net213
+ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
X_3154_ _1293_ _1323_ _1440_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__or3_1
XFILLER_82_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3085_ cordic_inst.cordic_inst.x\[26\] _1386_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__or2_1
XFILLER_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3987_ net61 net62 net63 VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__or3b_1
X_2938_ _1116_ _1131_ _1178_ net250 VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__a31o_1
X_2869_ net219 _1139_ _1143_ net221 VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__a22o_1
X_4608_ net377 _0340_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[26\] sky130_fd_sc_hd__dfxtp_1
X_4539_ net358 _0271_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3910_ axi_controller.read_addr_reg\[11\] net4 net195 VGND VGND VPWR VPWR _0277_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4890_ net378 _0043_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_3841_ axi_controller.state\[1\] net350 VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__nand2_1
X_3772_ axi_controller.reg_input_data\[28\] axi_controller.reg_input_data\[27\] axi_controller.reg_input_data\[26\]
+ axi_controller.reg_input_data\[25\] VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__and4_1
X_2723_ _0965_ _1041_ _0933_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__a21o_1
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2654_ cordic_inst.cordic_inst.y\[25\] _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__or2_1
XFILLER_8_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2585_ cordic_inst.cordic_inst.y\[15\] _0917_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__xnor2_1
X_4324_ net122 net194 net155 axi_controller.result_out\[19\] VGND VGND VPWR VPWR _0575_
+ sky130_fd_sc_hd__a22o_1
X_4255_ cordic_inst.cordic_inst.sin_out\[27\] net257 _2213_ VGND VGND VPWR VPWR _2215_
+ sky130_fd_sc_hd__nand3_1
X_3206_ cordic_inst.cordic_inst.y\[27\] cordic_inst.cordic_inst.sin_out\[27\] net207
+ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
X_4186_ net228 _2152_ _2153_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__or3_1
XFILLER_67_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3137_ _1343_ _1375_ _1420_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__nand3_1
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3068_ cordic_inst.cordic_inst.x\[23\] _1334_ _1337_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_53_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2370_ net293 net303 VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nor2_1
X_4040_ net100 _2019_ _2027_ net354 VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o211a_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4942_ net393 _0571_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_1
X_4873_ net382 axi_controller.reg_input_data\[5\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3824_ _1874_ _1915_ _1916_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3755_ cordic_inst.deg_handler_inst.theta_norm\[29\] _1862_ VGND VGND VPWR VPWR _0029_
+ sky130_fd_sc_hd__xnor2_1
X_3686_ cordic_inst.deg_handler_inst.theta_norm\[0\] cordic_inst.deg_handler_inst.theta_norm\[1\]
+ cordic_inst.deg_handler_inst.theta_norm\[3\] cordic_inst.deg_handler_inst.theta_norm\[2\]
+ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__or4_1
X_2706_ _0860_ _0861_ _0972_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2637_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2568_ cordic_inst.cordic_inst.y\[3\] _0888_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nor2_1
X_4307_ _1989_ _2253_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__nor2_1
X_2499_ _0793_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4238_ net257 _2199_ cordic_inst.cordic_inst.sin_out\[25\] VGND VGND VPWR VPWR _2200_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_59_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4169_ _2137_ _2138_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__or2_1
XFILLER_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3540_ cordic_inst.cordic_inst.angle\[2\] net172 net165 cordic_inst.cordic_inst.z\[2\]
+ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__a22o_1
X_3471_ _1488_ _1691_ _1486_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__a21o_1
X_2422_ _0750_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and2_1
X_2353_ _0673_ net219 _0687_ net221 net281 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a221o_1
XFILLER_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4023_ net103 _1963_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__and2_1
X_2284_ cordic_inst.state\[1\] VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4925_ net373 _0025_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_4856_ net386 _0065_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[20\] sky130_fd_sc_hd__dfxtp_1
X_3807_ axi_controller.reg_input_data\[26\] _1904_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__xnor2_1
X_4787_ net397 _0514_ _0209_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[16\] sky130_fd_sc_hd__dfrtp_4
X_3738_ cordic_inst.deg_handler_inst.theta_norm\[23\] _1851_ VGND VGND VPWR VPWR _0023_
+ sky130_fd_sc_hd__xnor2_1
X_3669_ _0617_ _1783_ _1808_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__or3_1
XFILLER_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2971_ _1269_ _1272_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__a21o_1
X_4710_ net403 _0437_ _0132_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4641_ net396 _0372_ net332 VGND VGND VPWR VPWR axi_controller.result_out\[18\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4572_ net372 _0304_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[5\] sky130_fd_sc_hd__dfxtp_1
X_3523_ cordic_inst.cordic_inst.angle\[8\] net172 net167 cordic_inst.cordic_inst.z\[8\]
+ _1738_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__a221o_1
X_3454_ _1478_ _1658_ _1659_ net176 VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__a31o_1
X_2405_ _0709_ _0729_ _0731_ _0713_ net282 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__a221o_1
X_3385_ _1538_ _1544_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2336_ net238 _0650_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nor2_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2267_ net270 VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__inv_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4006_ net106 _1963_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__nand2_2
XFILLER_25_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4908_ net390 _0038_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4839_ net391 _0078_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3170_ _1318_ _1321_ _1441_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__and3b_1
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2954_ cordic_inst.cordic_inst.x\[4\] _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__and2_1
X_2885_ _1098_ _1185_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__or3_1
X_4624_ net412 _0355_ net347 VGND VGND VPWR VPWR axi_controller.result_out\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4555_ net356 _0287_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[21\] sky130_fd_sc_hd__dfxtp_1
X_3506_ net183 _1724_ _1725_ _1726_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a31o_1
X_4486_ net340 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__inv_2
X_3437_ net249 cordic_inst.cordic_inst.z\[28\] _1667_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__a21oi_1
X_3368_ _1568_ _1606_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__nor2_1
X_2319_ cordic_inst.cordic_inst.x\[22\] cordic_inst.cordic_inst.x\[23\] cordic_inst.cordic_inst.x\[24\]
+ cordic_inst.cordic_inst.x\[25\] net306 net296 VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux4_1
XFILLER_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3299_ cordic_inst.cordic_inst.z\[11\] _1537_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2670_ _0810_ _1000_ _1003_ net174 VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a31o_1
X_4340_ net137 net193 net154 axi_controller.result_out\[3\] VGND VGND VPWR VPWR _0591_
+ sky130_fd_sc_hd__a22o_1
X_4271_ net316 _2224_ _2225_ _2228_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__a31o_1
X_3222_ cordic_inst.cordic_inst.y\[11\] cordic_inst.cordic_inst.sin_out\[11\] net213
+ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3153_ _1287_ _1290_ _1294_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__and3_1
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3084_ cordic_inst.cordic_inst.x\[26\] _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__nand2_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3986_ net107 net103 _1922_ _1943_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__nand4_1
X_2937_ _1236_ _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__and2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4607_ net377 _0339_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[25\] sky130_fd_sc_hd__dfxtp_1
X_2868_ _1132_ _1140_ net235 VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__mux2_1
X_2799_ net285 _1099_ _1101_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__a21oi_1
X_4538_ net358 _0270_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_4469_ net331 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3840_ net68 net35 axi_controller.state\[0\] net350 VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__and4b_1
X_3771_ axi_controller.reg_input_data\[22\] _1875_ axi_controller.reg_input_data\[23\]
+ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__a21oi_1
X_2722_ _0963_ _1039_ _0930_ _0939_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__o211ai_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2653_ _0802_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__xnor2_1
X_2584_ cordic_inst.cordic_inst.y\[15\] _0917_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__nor2_1
X_4323_ net124 net192 net155 axi_controller.result_out\[20\] VGND VGND VPWR VPWR _0574_
+ sky130_fd_sc_hd__a22o_1
X_4254_ net257 _2213_ cordic_inst.cordic_inst.sin_out\[27\] VGND VGND VPWR VPWR _2214_
+ sky130_fd_sc_hd__a21o_1
X_3205_ cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.sin_out\[28\] net207
+ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
X_4185_ net259 _2151_ cordic_inst.cordic_inst.sin_out\[19\] VGND VGND VPWR VPWR _2153_
+ sky130_fd_sc_hd__a21oi_1
X_3136_ _1427_ _1428_ cordic_inst.cordic_inst.x\[21\] net160 VGND VGND VPWR VPWR _0519_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3067_ _1335_ _1339_ _1346_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__or4_1
XFILLER_55_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3969_ axi_controller.write_addr_reg\[18\] net45 net188 VGND VGND VPWR VPWR _0317_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4941_ net367 _0570_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4872_ net382 axi_controller.reg_input_data\[4\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3823_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1872_
+ _1903_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_22_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3754_ cordic_inst.deg_handler_inst.theta_norm\[28\] _1859_ net253 VGND VGND VPWR
+ VPWR _1862_ sky130_fd_sc_hd__o21ai_1
X_3685_ cordic_inst.deg_handler_inst.theta_norm\[3\] _1818_ VGND VGND VPWR VPWR _0033_
+ sky130_fd_sc_hd__xor2_1
X_2705_ net180 _1021_ _1028_ net160 cordic_inst.cordic_inst.y\[20\] VGND VGND VPWR
+ VPWR _0550_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_30_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2636_ _0968_ _0970_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__nor2_1
X_2567_ _0899_ _0900_ _0892_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a21o_1
X_4306_ _1976_ _2252_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__nand2_1
X_2498_ net268 _0789_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__nand2_1
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4237_ cordic_inst.cordic_inst.sin_out\[24\] _2191_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__or2_1
X_4168_ cordic_inst.cordic_inst.sin_out\[17\] net259 _2136_ net228 VGND VGND VPWR
+ VPWR _2138_ sky130_fd_sc_hd__a31o_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3119_ net179 _1413_ _1416_ net162 cordic_inst.cordic_inst.x\[26\] VGND VGND VPWR
+ VPWR _0524_ sky130_fd_sc_hd__a32o_1
X_4099_ _2076_ _2077_ net203 _2074_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__o211a_1
XFILLER_70_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3470_ _1486_ _1488_ _1691_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__nand3_1
X_2421_ net247 _0755_ _0753_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__o21ai_1
X_2352_ cordic_inst.cordic_inst.x\[6\] cordic_inst.cordic_inst.x\[7\] cordic_inst.cordic_inst.x\[8\]
+ cordic_inst.cordic_inst.x\[9\] net315 net302 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__mux4_1
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2283_ axi_controller.state\[1\] VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__inv_2
X_4022_ net95 _2009_ _2017_ net352 VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_35_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4924_ net373 _0024_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_4855_ net384 _0063_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[19\] sky130_fd_sc_hd__dfxtp_1
X_3806_ _1903_ _1899_ axi_controller.reg_input_data\[25\] VGND VGND VPWR VPWR _1904_
+ sky130_fd_sc_hd__mux2_1
X_4786_ net397 _0513_ _0208_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3737_ cordic_inst.deg_handler_inst.theta_norm\[22\] _1849_ net254 VGND VGND VPWR
+ VPWR _1851_ sky130_fd_sc_hd__o21ai_1
X_3668_ cordic_inst.deg_handler_inst.theta_abs\[21\] net149 net148 _1813_ VGND VGND
+ VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
X_3599_ cordic_inst.deg_handler_inst.theta_abs\[10\] _1766_ VGND VGND VPWR VPWR _1767_
+ sky130_fd_sc_hd__or2_1
X_2619_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__inv_2
XFILLER_87_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout290 cordic_inst.cordic_inst.i\[3\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2970_ cordic_inst.cordic_inst.x\[2\] _1265_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__xnor2_1
X_4640_ net398 _0371_ net332 VGND VGND VPWR VPWR axi_controller.result_out\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4571_ net372 _0303_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_3522_ _1611_ _1618_ _1737_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__o21a_1
X_3453_ _1478_ _1658_ _1659_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__a21oi_1
X_2404_ _0668_ _0681_ net235 VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__mux2_1
X_3384_ _1616_ _1619_ _1620_ _1550_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__o31a_1
X_2335_ net283 _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__nor2_1
X_2266_ cordic_inst.cordic_inst.x\[0\] VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__inv_2
X_4005_ net106 _1963_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__and2_1
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4907_ net390 _0037_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_4838_ net391 _0075_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[2\] sky130_fd_sc_hd__dfxtp_1
X_4769_ net364 _0496_ _0191_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2953_ _1177_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__xnor2_1
X_2884_ cordic_inst.cordic_inst.y\[31\] _1161_ _1162_ _1158_ net245 net241 VGND VGND
+ VPWR VPWR _1187_ sky130_fd_sc_hd__mux4_1
X_4623_ net373 _0354_ net338 VGND VGND VPWR VPWR axi_controller.result_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_4554_ net357 _0286_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[20\] sky130_fd_sc_hd__dfxtp_1
X_3505_ cordic_inst.cordic_inst.angle\[13\] net173 net165 cordic_inst.cordic_inst.z\[13\]
+ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__a22o_1
X_4485_ net327 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__inv_2
X_3436_ cordic_inst.cordic_inst.z\[30\] net157 _1673_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__o21a_1
X_3367_ _1575_ _1605_ _1570_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__a21boi_1
X_2318_ cordic_inst.cordic_inst.x\[18\] cordic_inst.cordic_inst.x\[19\] cordic_inst.cordic_inst.x\[20\]
+ cordic_inst.cordic_inst.x\[21\] net308 net298 VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux4_1
X_3298_ net274 _1504_ _1536_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__mux2_1
XFILLER_72_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput100 wdata[7] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4270_ net316 _2226_ _2227_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__nor3b_1
X_3221_ cordic_inst.cordic_inst.y\[12\] cordic_inst.cordic_inst.sin_out\[12\] net213
+ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
X_3152_ _1287_ _1290_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__nand2_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3083_ _1213_ _1223_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3985_ _0624_ _1994_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__nor2_1
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2936_ cordic_inst.cordic_inst.x\[28\] _1235_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__or2_1
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2867_ _1148_ _1157_ _1164_ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__or4b_2
X_4606_ net376 _0338_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[24\] sky130_fd_sc_hd__dfxtp_1
X_2798_ net219 _1095_ _1100_ net221 net279 VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__a221o_1
X_4537_ net358 _0269_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_4468_ net331 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__inv_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3419_ _1655_ _1657_ _1480_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__a21o_1
X_4399_ net347 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_26_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3770_ axi_controller.reg_input_data\[19\] axi_controller.reg_input_data\[18\] axi_controller.reg_input_data\[21\]
+ axi_controller.reg_input_data\[20\] VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__a211o_1
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2721_ _0963_ _1039_ _0939_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__o21a_1
X_2652_ net169 _0796_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__nor2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2583_ cordic_inst.cordic_inst.y\[15\] _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nand2_1
X_4322_ net125 net192 net155 axi_controller.result_out\[21\] VGND VGND VPWR VPWR _0573_
+ sky130_fd_sc_hd__a22o_1
X_4253_ cordic_inst.cordic_inst.sin_out\[26\] cordic_inst.cordic_inst.sin_out\[25\]
+ _2199_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__or3_1
X_3204_ cordic_inst.cordic_inst.y\[29\] cordic_inst.cordic_inst.sin_out\[29\] net207
+ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux2_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4184_ cordic_inst.cordic_inst.sin_out\[19\] net259 _2151_ VGND VGND VPWR VPWR _2152_
+ sky130_fd_sc_hd__and3_1
X_3135_ _1341_ _1348_ _1421_ net175 VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__a31o_1
X_3066_ _1341_ _1347_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3968_ axi_controller.write_addr_reg\[17\] net44 net188 VGND VGND VPWR VPWR _0316_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2919_ net268 _1211_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__a21o_1
X_3899_ axi_controller.read_addr_reg\[0\] net2 net198 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
XFILLER_18_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4940_ net366 _0569_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_1
XFILLER_91_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4871_ net380 axi_controller.reg_input_data\[3\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3822_ _1880_ _1914_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3753_ cordic_inst.deg_handler_inst.theta_norm\[28\] _1859_ VGND VGND VPWR VPWR _1861_
+ sky130_fd_sc_hd__nor2_1
X_3684_ cordic_inst.deg_handler_inst.theta_norm\[0\] cordic_inst.deg_handler_inst.theta_norm\[1\]
+ cordic_inst.deg_handler_inst.theta_norm\[2\] net255 VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__o31a_1
X_2704_ _0837_ _0864_ _0973_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_30_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2635_ _0860_ _0969_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__nand2_1
X_4305_ axi_controller.read_addr_reg\[5\] _1977_ axi_controller.read_addr_reg\[3\]
+ axi_controller.read_addr_reg\[4\] VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__and4b_1
X_2566_ _0899_ _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__nand2_1
X_2497_ _0825_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nand2_1
X_4236_ net223 _2196_ cordic_inst.cordic_inst.cos_out\[25\] VGND VGND VPWR VPWR _2198_
+ sky130_fd_sc_hd__a21oi_1
X_4167_ net259 _2136_ cordic_inst.cordic_inst.sin_out\[17\] VGND VGND VPWR VPWR _2137_
+ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_27_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3118_ _1390_ _1412_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4098_ cordic_inst.cordic_inst.sin_out\[8\] net261 _2075_ net229 VGND VGND VPWR VPWR
+ _2077_ sky130_fd_sc_hd__a31o_1
X_3049_ _1203_ _1351_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_36_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_45_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2420_ net265 _0722_ _0723_ _0720_ net240 net233 VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__mux4_1
X_2351_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__inv_2
X_2282_ cordic_inst.state\[0\] VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_63_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4021_ axi_controller.reg_input_data\[31\] _2008_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4923_ net373 _0023_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_72_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4854_ net389 _0062_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3805_ _1901_ _1903_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4785_ net397 _0512_ _0207_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[14\] sky130_fd_sc_hd__dfrtp_4
X_3736_ cordic_inst.deg_handler_inst.theta_norm\[22\] _1850_ VGND VGND VPWR VPWR _0022_
+ sky130_fd_sc_hd__xnor2_1
X_3667_ _1783_ _1808_ _1812_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__o21ai_1
X_3598_ cordic_inst.deg_handler_inst.theta_abs\[9\] _1765_ VGND VGND VPWR VPWR _1766_
+ sky130_fd_sc_hd__or2_1
X_2618_ cordic_inst.cordic_inst.y\[9\] _0951_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_81_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2549_ _0599_ _0882_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__nand2_1
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4219_ cordic_inst.cordic_inst.sin_out\[23\] net258 _2180_ _2182_ VGND VGND VPWR
+ VPWR _2183_ sky130_fd_sc_hd__a31o_1
XFILLER_75_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout280 cordic_inst.cordic_inst.i\[4\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_2
Xfanout291 net292 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4570_ net370 _0302_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_3521_ net176 _1619_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3452_ net182 _1680_ _1684_ _1685_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a31o_1
X_3383_ _1551_ _1620_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__nor2_1
XFILLER_69_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2403_ net247 _0659_ _0736_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__o22a_1
X_2334_ _0660_ _0668_ net235 VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux2_1
XFILLER_84_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2265_ cordic_inst.cordic_inst.x\[5\] VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__inv_2
XFILLER_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4004_ net146 _1943_ _2002_ _2007_ net350 VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o221a_1
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4906_ net391 _0036_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4837_ net403 _0064_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[1\] sky130_fd_sc_hd__dfxtp_1
X_4768_ net366 _0495_ _0190_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_3719_ net256 _1839_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__nand2_1
X_4699_ net367 _0426_ _0121_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2952_ net276 _1170_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__nand2_1
X_2883_ net238 _1162_ _1070_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__a21bo_1
X_4622_ net381 _0353_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[7\] sky130_fd_sc_hd__dfxtp_1
X_4553_ net356 _0285_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[19\] sky130_fd_sc_hd__dfxtp_1
X_3504_ _1514_ _1627_ _1533_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__a21o_1
X_4484_ net327 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__inv_2
X_3435_ cordic_inst.cordic_inst.angle\[30\] net174 _1670_ _1672_ net163 VGND VGND
+ VPWR VPWR _1673_ sky130_fd_sc_hd__a221o_1
X_3366_ _1591_ _1602_ _1604_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__o21ai_1
X_3297_ net302 net314 _0706_ net293 _0713_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__a221o_1
X_2317_ net278 _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__nor2_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput101 wdata[8] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3220_ cordic_inst.cordic_inst.y\[13\] cordic_inst.cordic_inst.sin_out\[13\] net210
+ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__mux2_1
X_3151_ net180 _1430_ _1438_ net160 cordic_inst.cordic_inst.x\[16\] VGND VGND VPWR
+ VPWR _0514_ sky130_fd_sc_hd__a32o_1
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3082_ cordic_inst.cordic_inst.x\[27\] _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__xor2_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3984_ _1993_ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__inv_2
X_2935_ cordic_inst.cordic_inst.x\[29\] _1233_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nand2_1
X_2866_ _1165_ _1166_ _1168_ net281 VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__a2bb2o_1
X_4605_ net374 _0337_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_1
X_2797_ cordic_inst.cordic_inst.y\[7\] cordic_inst.cordic_inst.y\[8\] cordic_inst.cordic_inst.y\[9\]
+ cordic_inst.cordic_inst.y\[10\] net310 net300 VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__mux4_1
X_4536_ net356 _0268_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_4467_ net334 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4398_ net347 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__inv_2
X_3418_ net249 cordic_inst.cordic_inst.z\[23\] _1491_ _1656_ VGND VGND VPWR VPWR _1657_
+ sky130_fd_sc_hd__a211oi_1
X_3349_ net274 _1587_ _1585_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__a21oi_1
XFILLER_85_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2720_ _0947_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__nor2_1
X_2651_ cordic_inst.cordic_inst.y\[26\] _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__xor2_1
X_2582_ _0672_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__xnor2_2
X_4321_ net126 net191 net156 axi_controller.result_out\[22\] VGND VGND VPWR VPWR _0572_
+ sky130_fd_sc_hd__a22o_1
X_4252_ cordic_inst.cordic_inst.cos_out\[27\] _2210_ net316 VGND VGND VPWR VPWR _2212_
+ sky130_fd_sc_hd__a21o_1
XFILLER_4_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3203_ cordic_inst.cordic_inst.y\[30\] cordic_inst.cordic_inst.sin_out\[30\] net207
+ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__mux2_1
X_4183_ cordic_inst.cordic_inst.sin_out\[18\] _2143_ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__or2_1
X_3134_ _1341_ _1421_ _1348_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3065_ _1349_ _1359_ _1362_ _1367_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__nor4_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3967_ axi_controller.write_addr_reg\[16\] net43 net188 VGND VGND VPWR VPWR _0315_
+ sky130_fd_sc_hd__mux2_1
X_2918_ net269 _1090_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__a21o_1
XFILLER_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3898_ net77 _1965_ _1973_ net353 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__o211a_1
X_2849_ _1117_ _1122_ net236 VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__mux2_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4519_ net374 _0006_ _0085_ VGND VGND VPWR VPWR cordic_inst.state\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_85_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4870_ net380 axi_controller.reg_input_data\[2\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3821_ _1878_ _1898_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__nor2_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3752_ cordic_inst.deg_handler_inst.theta_norm\[28\] _1860_ VGND VGND VPWR VPWR _0028_
+ sky130_fd_sc_hd__xnor2_1
X_3683_ cordic_inst.deg_handler_inst.theta_norm\[2\] _1817_ VGND VGND VPWR VPWR _0030_
+ sky130_fd_sc_hd__xnor2_1
X_2703_ cordic_inst.cordic_inst.y\[21\] net160 _1027_ net180 VGND VGND VPWR VPWR _0551_
+ sky130_fd_sc_hd__a22o_1
X_2634_ cordic_inst.cordic_inst.y\[16\] _0859_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__or2_1
X_2565_ cordic_inst.cordic_inst.y\[2\] _0891_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__xor2_1
X_4304_ net86 _2243_ _2251_ net351 VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o211a_1
XFILLER_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2496_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__inv_2
XFILLER_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4235_ cordic_inst.cordic_inst.cos_out\[25\] net223 _2196_ VGND VGND VPWR VPWR _2197_
+ sky130_fd_sc_hd__and3_1
XFILLER_59_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4166_ cordic_inst.cordic_inst.sin_out\[16\] _2128_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__or2_1
X_3117_ cordic_inst.cordic_inst.x\[27\] net162 _1415_ net174 VGND VGND VPWR VPWR _0525_
+ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_66_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4097_ net261 _2075_ cordic_inst.cordic_inst.sin_out\[8\] VGND VGND VPWR VPWR _2076_
+ sky130_fd_sc_hd__a21oi_1
X_3048_ _1195_ _1198_ _1202_ _1204_ net271 VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__o41a_1
XFILLER_51_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2350_ _0653_ _0674_ net236 VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux2_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2281_ cordic_inst.deg_handler_inst.theta_abs\[22\] VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__inv_2
X_4020_ net94 _2009_ _2016_ net352 VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o211a_1
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4922_ net373 _0022_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_4853_ net387 _0061_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[17\] sky130_fd_sc_hd__dfxtp_1
X_3804_ _1874_ _1902_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__or2_1
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4784_ net401 _0511_ _0206_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[13\] sky130_fd_sc_hd__dfrtp_4
X_3735_ net253 _1849_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__nand2_1
X_3666_ _0616_ _1808_ cordic_inst.deg_handler_inst.theta_abs\[21\] VGND VGND VPWR
+ VPWR _1812_ sky130_fd_sc_hd__o21bai_1
X_3597_ cordic_inst.deg_handler_inst.theta_abs\[8\] _1764_ VGND VGND VPWR VPWR _1765_
+ sky130_fd_sc_hd__or2_1
X_2617_ cordic_inst.cordic_inst.y\[9\] _0951_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__nand2_1
X_2548_ _0599_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and2_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4218_ net317 _2181_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__nand2_1
X_2479_ _0806_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_87_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4149_ net225 _2120_ cordic_inst.cordic_inst.cos_out\[15\] VGND VGND VPWR VPWR _2121_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__buf_2
Xfanout292 net295 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_4
Xfanout281 net282 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_2
XFILLER_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3520_ net185 _1734_ _1735_ _1736_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__a31o_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3451_ cordic_inst.cordic_inst.angle\[26\] net170 net163 cordic_inst.cordic_inst.z\[26\]
+ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__a22o_1
X_3382_ _1550_ _1616_ _1620_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__a21oi_1
X_2402_ net286 _0675_ net220 _0687_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__a22o_1
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2333_ cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.x\[16\] cordic_inst.cordic_inst.x\[17\]
+ cordic_inst.cordic_inst.x\[18\] net308 net298 VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__mux4_1
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2264_ net267 VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__inv_2
X_4003_ net68 _0622_ _0624_ _1923_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4905_ net390 _0035_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4836_ net387 _0053_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4767_ net366 _0494_ _0189_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_3718_ cordic_inst.deg_handler_inst.theta_norm\[15\] _1837_ VGND VGND VPWR VPWR _1839_
+ sky130_fd_sc_hd__or2_1
X_4698_ net368 _0425_ _0120_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3649_ cordic_inst.deg_handler_inst.theta_abs\[13\] _1769_ VGND VGND VPWR VPWR _1803_
+ sky130_fd_sc_hd__nand2_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2951_ _1253_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__inv_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4621_ net380 _0352_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2882_ _1182_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or2_1
X_4552_ net356 _0284_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[18\] sky130_fd_sc_hd__dfxtp_1
X_3503_ _1514_ _1533_ _1627_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__nand3_1
X_4483_ net327 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__inv_2
X_3434_ _1474_ _1669_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__or2_1
X_3365_ _1575_ _1603_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__and2_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3296_ _1514_ _1534_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__nand2_1
X_2316_ net239 _0650_ _0637_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_0_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4819_ net395 _0546_ _0241_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput102 wdata[9] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3150_ _1332_ _1361_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__or2_1
X_3081_ _1224_ _1383_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3983_ axi_controller.write_addr_reg\[3\] axi_controller.write_addr_reg\[4\] _1953_
+ axi_controller.write_addr_reg\[5\] VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__or4b_1
X_2934_ cordic_inst.cordic_inst.x\[29\] _1233_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__and2_1
X_2865_ net285 _1094_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4604_ net371 _0336_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4535_ net358 _0267_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_2796_ _1093_ _1096_ net235 VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux2_1
X_4466_ net334 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__inv_2
X_4397_ net346 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
X_3417_ _1495_ _1497_ _1654_ _1496_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_90_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3348_ _1564_ _1586_ _1577_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__a21o_1
XFILLER_58_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3279_ cordic_inst.cordic_inst.z\[14\] _1517_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__and2_1
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2650_ _0797_ _0803_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__xor2_2
X_2581_ _0770_ _0780_ net252 VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a21oi_1
X_4320_ net127 net192 net156 axi_controller.result_out\[23\] VGND VGND VPWR VPWR _0571_
+ sky130_fd_sc_hd__a22o_1
X_4251_ cordic_inst.cordic_inst.cos_out\[27\] _2210_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3202_ net264 cordic_inst.cordic_inst.sin_out\[31\] net208 VGND VGND VPWR VPWR _0497_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4182_ _2146_ _2150_ axi_controller.result_out\[18\] net201 VGND VGND VPWR VPWR _0372_
+ sky130_fd_sc_hd__o2bb2a_1
X_3133_ net178 _1423_ _1426_ net159 cordic_inst.cordic_inst.x\[22\] VGND VGND VPWR
+ VPWR _0520_ sky130_fd_sc_hd__a32o_1
X_3064_ _1365_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__or2_1
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3966_ axi_controller.write_addr_reg\[15\] net42 net189 VGND VGND VPWR VPWR _0314_
+ sky130_fd_sc_hd__mux2_1
X_2917_ net272 _1210_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_61_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3897_ axi_controller.reg_input_data\[15\] _1964_ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__or2_1
XFILLER_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2848_ _1149_ _1150_ net285 VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__mux2_1
X_2779_ net246 _1081_ net215 VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__a21o_1
X_4518_ net337 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__inv_2
X_4449_ net321 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__inv_2
XFILLER_85_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3820_ axi_controller.reg_input_data\[30\] _1913_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__xor2_1
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3751_ net253 _1859_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__nand2_1
X_2702_ _0843_ _1022_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__xnor2_1
X_3682_ cordic_inst.deg_handler_inst.theta_norm\[0\] cordic_inst.deg_handler_inst.theta_norm\[1\]
+ net255 VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_30_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2633_ _0961_ _0966_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__and3_2
X_2564_ _0896_ _0897_ _0895_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__o21ai_1
X_4303_ axi_controller.reg_input_data\[23\] _2242_ VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__or2_1
XFILLER_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2495_ cordic_inst.cordic_inst.y\[23\] _0827_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4234_ cordic_inst.cordic_inst.cos_out\[24\] _2188_ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__or2_1
X_4165_ axi_controller.result_out\[16\] _2135_ net201 VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
X_3116_ _1385_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_66_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4096_ cordic_inst.cordic_inst.sin_out\[7\] _2065_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__or2_1
X_3047_ net271 _1202_ _1217_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3949_ _0619_ _1991_ axi_controller.reg_done_flag VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__o21a_1
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2280_ cordic_inst.deg_handler_inst.theta_abs\[20\] VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__inv_2
XFILLER_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4921_ net379 _0021_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_4852_ net387 _0060_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[16\] sky130_fd_sc_hd__dfxtp_1
X_3803_ axi_controller.reg_input_data\[23\] _1890_ axi_controller.reg_input_data\[24\]
+ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__o21a_1
X_4783_ net401 _0510_ _0205_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[12\] sky130_fd_sc_hd__dfrtp_4
X_3734_ cordic_inst.deg_handler_inst.theta_norm\[21\] _1847_ VGND VGND VPWR VPWR _1849_
+ sky130_fd_sc_hd__or2_1
XFILLER_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3665_ cordic_inst.deg_handler_inst.theta_abs\[20\] net150 net148 _1811_ VGND VGND
+ VPWR VPWR _0065_ sky130_fd_sc_hd__a22o_1
X_2616_ _0762_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__xnor2_1
X_3596_ cordic_inst.deg_handler_inst.theta_abs\[7\] _1763_ VGND VGND VPWR VPWR _1764_
+ sky130_fd_sc_hd__or2_1
X_2547_ _0756_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__xnor2_1
X_2478_ net169 _0807_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__nor2_1
X_4217_ net258 _2180_ cordic_inst.cordic_inst.sin_out\[23\] VGND VGND VPWR VPWR _2181_
+ sky130_fd_sc_hd__a21o_1
XFILLER_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4148_ cordic_inst.cordic_inst.cos_out\[14\] cordic_inst.cordic_inst.cos_out\[13\]
+ _2111_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__or3_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4079_ cordic_inst.cordic_inst.sin_out\[5\] cordic_inst.cordic_inst.sin_out\[4\]
+ _2045_ net262 VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__o31a_1
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_2
Xfanout271 net272 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__buf_2
Xfanout282 cordic_inst.cordic_inst.i\[4\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_2
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout293 net294 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__buf_2
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3450_ _1661_ _1663_ _1679_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__or3_1
X_3381_ cordic_inst.cordic_inst.z\[9\] _1549_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__and2_1
X_2401_ _0703_ _0709_ _0710_ _0713_ net282 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__a221o_1
X_2332_ net244 _0659_ net169 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__a21o_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4002_ _1921_ _2006_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nor2_1
X_2263_ cordic_inst.cordic_inst.y\[0\] VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4904_ net390 _0034_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4835_ net384 _0008_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.isNegative
+ sky130_fd_sc_hd__dfxtp_4
X_4766_ net365 _0493_ _0188_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_3717_ cordic_inst.deg_handler_inst.theta_norm\[15\] _1838_ VGND VGND VPWR VPWR _0014_
+ sky130_fd_sc_hd__xnor2_1
X_4697_ net367 _0424_ _0119_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_3648_ _1769_ net147 _1802_ net151 cordic_inst.deg_handler_inst.theta_abs\[12\] VGND
+ VGND VPWR VPWR _0056_ sky130_fd_sc_hd__a32o_1
XFILLER_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3579_ cordic_inst.cordic_inst.x\[0\] cordic_inst.cordic_inst.cos_out\[0\] net212
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2950_ _0602_ _1251_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__nor2_1
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2881_ net263 _1134_ _1136_ _1141_ net245 net241 VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__mux4_2
X_4620_ net381 _0351_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[5\] sky130_fd_sc_hd__dfxtp_1
X_4551_ net357 _0283_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[17\] sky130_fd_sc_hd__dfxtp_1
X_3502_ cordic_inst.cordic_inst.angle\[14\] net173 net168 cordic_inst.cordic_inst.z\[14\]
+ _1723_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a221o_1
X_4482_ net327 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__inv_2
X_3433_ net273 net157 _1671_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o21a_1
X_3364_ cordic_inst.cordic_inst.z\[4\] _1574_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__or2_1
X_3295_ cordic_inst.cordic_inst.z\[12\] _1513_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__or2_1
X_2315_ _0646_ _0649_ net291 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_69_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4818_ net401 _0545_ _0240_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[15\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_78_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4749_ net400 _0476_ _0171_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput103 wstrb[0] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3080_ net215 _1214_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__or2_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3982_ axi_controller.write_addr_reg\[31\] net60 net188 VGND VGND VPWR VPWR _0330_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2933_ cordic_inst.cordic_inst.x\[28\] _1235_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__nand2_1
X_2864_ net235 _1087_ _1071_ net241 VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a211o_1
X_2795_ cordic_inst.cordic_inst.y\[31\] _1091_ _1094_ _1097_ net241 net245 VGND VGND
+ VPWR VPWR _1098_ sky130_fd_sc_hd__mux4_1
X_4603_ net371 _0335_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
X_4534_ net360 _0266_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4465_ net334 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__inv_2
X_4396_ net346 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_2
X_3416_ _1532_ _1628_ _1649_ _1496_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_90_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ net242 net313 net293 VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__o21a_1
XFILLER_58_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3278_ net273 _1481_ _1516_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__mux2_1
XFILLER_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2580_ _0873_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nor2_1
X_4250_ cordic_inst.deg_handler_inst.kuadran\[0\] _2204_ VGND VGND VPWR VPWR _2210_
+ sky130_fd_sc_hd__nor2_1
X_4181_ _2148_ _2149_ net201 VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__o21a_1
X_3201_ cordic_inst.cordic_inst.state\[1\] cordic_inst.cordic_inst.state\[0\] VGND
+ VGND VPWR VPWR _1472_ sky130_fd_sc_hd__nand2_1
X_3132_ _1339_ _1422_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__nand2_1
XFILLER_67_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3063_ cordic_inst.cordic_inst.x\[17\] _1364_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__and2_1
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3965_ axi_controller.write_addr_reg\[14\] net41 net189 VGND VGND VPWR VPWR _0313_
+ sky130_fd_sc_hd__mux2_1
X_3896_ net76 _1965_ _1972_ net352 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__o211a_1
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2916_ net271 _1209_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_61_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2847_ net264 _1085_ _1086_ _1083_ net232 net231 VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__mux4_2
X_2778_ net238 _1080_ _1070_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__a21bo_1
X_4517_ net326 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__inv_2
X_4448_ net321 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__inv_2
X_4379_ net329 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3750_ cordic_inst.deg_handler_inst.theta_norm\[27\] _1857_ VGND VGND VPWR VPWR _1859_
+ sky130_fd_sc_hd__or2_1
X_2701_ cordic_inst.cordic_inst.y\[22\] net158 _1026_ net178 VGND VGND VPWR VPWR _0552_
+ sky130_fd_sc_hd__a22o_1
X_3681_ cordic_inst.deg_handler_inst.theta_norm\[1\] _1816_ VGND VGND VPWR VPWR _0019_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_9_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2632_ _0926_ _0933_ _0965_ _0964_ _0936_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__o32a_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2563_ _0896_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__or2_1
X_4302_ net85 _2243_ _2250_ net351 VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o211a_1
X_2494_ cordic_inst.cordic_inst.y\[23\] _0827_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__nor2_1
X_4233_ net200 _2195_ _2187_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4164_ _2133_ _2134_ _2131_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__o21ai_1
X_3115_ _1387_ _1413_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__nand2_1
X_4095_ cordic_inst.cordic_inst.cos_out\[8\] _2072_ _2073_ VGND VGND VPWR VPWR _2074_
+ sky130_fd_sc_hd__a21o_1
X_3046_ _1335_ _1339_ _1343_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__or4_1
XFILLER_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3948_ net70 _1990_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__nand2_1
X_3879_ net107 axi_controller.state\[3\] _1961_ _1942_ axi_controller.state\[0\] VGND
+ VGND VPWR VPWR _1962_ sky130_fd_sc_hd__a32o_1
XFILLER_73_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4920_ net379 _0020_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4851_ net387 _0059_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[15\] sky130_fd_sc_hd__dfxtp_1
X_3802_ axi_controller.reg_input_data\[25\] _1899_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__xnor2_1
X_4782_ net399 _0509_ _0204_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_60_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3733_ cordic_inst.deg_handler_inst.theta_norm\[21\] _1848_ VGND VGND VPWR VPWR _0021_
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_41_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3664_ _0616_ _1808_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__xnor2_1
X_2615_ net276 _0760_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a21oi_1
X_3595_ cordic_inst.deg_handler_inst.theta_abs\[6\] _1762_ VGND VGND VPWR VPWR _1763_
+ sky130_fd_sc_hd__or2_1
X_2546_ _0743_ _0750_ net250 VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__a21o_1
X_2477_ _0810_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nand2_1
X_4216_ cordic_inst.cordic_inst.sin_out\[22\] _2176_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__or2_1
X_4147_ axi_controller.result_out\[14\] _2119_ net201 VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4078_ cordic_inst.cordic_inst.cos_out\[6\] _2058_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__xor2_1
X_3029_ _1328_ _1331_ _1325_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__nand3b_2
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout250 net251 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_77_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout272 cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_2
Xfanout283 net290 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_4
Xfanout261 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__buf_2
XFILLER_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout294 net295 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__buf_2
XFILLER_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2400_ net248 _0725_ _0734_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__o21a_1
X_3380_ _1611_ _1618_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__and2_1
X_2331_ net169 _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nor2_1
X_2262_ cordic_inst.cordic_inst.y\[5\] VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__inv_2
XFILLER_84_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4001_ net111 _0610_ axi_controller.state\[2\] VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__a21oi_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4903_ net390 _0033_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4834_ net369 _0561_ _0256_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[31\] sky130_fd_sc_hd__dfrtp_1
X_4765_ net365 _0492_ _0187_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_3716_ net256 _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__nand2_1
X_4696_ net393 _0423_ _0118_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3647_ cordic_inst.deg_handler_inst.theta_abs\[12\] _1768_ VGND VGND VPWR VPWR _1802_
+ sky130_fd_sc_hd__nand2_1
X_3578_ cordic_inst.cordic_inst.x\[1\] cordic_inst.cordic_inst.cos_out\[1\] net211
+ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux2_1
XFILLER_88_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2529_ _0850_ _0854_ _0862_ _0863_ _0848_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__o32a_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ net238 _1136_ _1070_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4550_ net356 _0282_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[16\] sky130_fd_sc_hd__dfxtp_1
X_3501_ _1520_ _1717_ _1722_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__a21boi_1
X_4481_ net326 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__inv_2
X_3432_ _0614_ cordic_inst.cordic_inst.angle\[31\] _1473_ _1670_ net163 VGND VGND
+ VPWR VPWR _1671_ sky130_fd_sc_hd__a221o_1
X_3363_ _1594_ _1601_ _1592_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__a21oi_1
XFILLER_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3294_ _1506_ _1530_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__or2_1
X_2314_ cordic_inst.cordic_inst.x\[27\] cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.x\[29\]
+ cordic_inst.cordic_inst.x\[30\] net307 net297 VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux4_1
XFILLER_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4817_ net401 _0544_ _0239_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[14\] sky130_fd_sc_hd__dfrtp_4
X_4748_ net409 _0475_ _0170_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4679_ net410 _0406_ _0101_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput104 wstrb[1] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3981_ axi_controller.write_addr_reg\[30\] net59 net188 VGND VGND VPWR VPWR _0329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2932_ _1082_ _1225_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__xnor2_1
X_2863_ net286 _1097_ _1100_ net219 VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a22o_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2794_ _1095_ _1096_ net292 VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__mux2_1
X_4602_ net372 _0334_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
X_4533_ net381 _0265_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[15\] sky130_fd_sc_hd__dfxtp_1
X_4464_ net334 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__inv_2
X_4395_ net346 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
XFILLER_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3415_ _1637_ _1653_ _1652_ _1642_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_90_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _1583_ _1584_ net251 VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3277_ net220 _0712_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_56_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4180_ cordic_inst.cordic_inst.cos_out\[18\] net224 _2147_ net319 VGND VGND VPWR
+ VPWR _2149_ sky130_fd_sc_hd__a31o_1
X_3200_ _0603_ _1471_ _1470_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
X_3131_ _1424_ _1425_ cordic_inst.cordic_inst.x\[23\] net158 VGND VGND VPWR VPWR _0521_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3062_ cordic_inst.cordic_inst.x\[17\] _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__nor2_1
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3964_ axi_controller.write_addr_reg\[13\] net40 net189 VGND VGND VPWR VPWR _0312_
+ sky130_fd_sc_hd__mux2_1
X_3895_ axi_controller.reg_input_data\[14\] _1964_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__or2_1
X_2915_ _1195_ _1198_ _1205_ net271 VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_61_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2846_ _1118_ _1125_ net291 VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__mux2_1
X_2777_ net234 _1079_ _1071_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__a21o_1
X_4516_ net322 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__inv_2
X_4447_ net323 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__inv_2
X_4378_ net330 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
X_3329_ cordic_inst.cordic_inst.z\[5\] _1567_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2700_ _0825_ _1023_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__xor2_1
X_3680_ cordic_inst.deg_handler_inst.theta_norm\[0\] net255 VGND VGND VPWR VPWR _1816_
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2631_ _0918_ _0924_ _0919_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a21o_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2562_ cordic_inst.cordic_inst.y\[1\] _0894_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__xnor2_1
X_4301_ axi_controller.reg_input_data\[22\] _2242_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__or2_1
X_2493_ cordic_inst.cordic_inst.y\[23\] _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__nand2_1
X_4232_ _2189_ _2190_ _2194_ net228 VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__o22a_1
X_4163_ cordic_inst.cordic_inst.cos_out\[16\] net224 _2132_ net318 VGND VGND VPWR
+ VPWR _2134_ sky130_fd_sc_hd__a31o_1
X_3114_ _1390_ _1412_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__or2_1
X_4094_ cordic_inst.cordic_inst.cos_out\[8\] _2072_ net229 VGND VGND VPWR VPWR _2073_
+ sky130_fd_sc_hd__o21ai_1
X_3045_ _1346_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__nand2b_1
XFILLER_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3947_ _1979_ _1989_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__nor2_2
X_3878_ _0623_ _1950_ _1954_ _1960_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__or4_1
X_2829_ cordic_inst.cordic_inst.y\[16\] cordic_inst.cordic_inst.y\[17\] cordic_inst.cordic_inst.y\[18\]
+ cordic_inst.cordic_inst.y\[19\] net308 net301 VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux4_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout410 net411 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ net387 _0058_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3801_ _1899_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4781_ net399 _0508_ _0203_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[10\] sky130_fd_sc_hd__dfrtp_4
X_3732_ net254 _1847_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__nand2_1
X_3663_ cordic_inst.deg_handler_inst.theta_abs\[19\] net149 net148 _1810_ VGND VGND
+ VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
X_2614_ net153 _0758_ net250 VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__a21oi_1
X_3594_ cordic_inst.deg_handler_inst.theta_abs\[5\] _1761_ VGND VGND VPWR VPWR _1762_
+ sky130_fd_sc_hd__or2_1
X_2545_ net250 _0743_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nor2_1
X_2476_ cordic_inst.cordic_inst.y\[30\] _0809_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__or2_1
X_4215_ axi_controller.result_out\[22\] _2179_ net200 VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_1
X_4146_ _2116_ _2118_ net228 VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__mux2_1
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ cordic_inst.cordic_inst.cos_out\[5\] cordic_inst.cordic_inst.cos_out\[4\]
+ _2048_ net226 VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__o31a_1
X_3028_ _1329_ _1330_ _1313_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__a21bo_1
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout240 net241 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout273 net277 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__buf_4
Xfanout251 net252 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_2
XFILLER_59_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout262 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout284 net290 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_2
Xfanout295 cordic_inst.cordic_inst.i\[2\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__buf_2
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2330_ net279 _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__nor2_1
X_2261_ cordic_inst.cordic_inst.y\[8\] VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__inv_2
XFILLER_84_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4000_ _0621_ _2005_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nor2_1
XFILLER_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4902_ net389 _0030_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4833_ net366 _0560_ _0255_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[30\] sky130_fd_sc_hd__dfrtp_2
X_4764_ net367 _0491_ _0186_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_3715_ cordic_inst.deg_handler_inst.theta_norm\[14\] cordic_inst.deg_handler_inst.theta_norm\[13\]
+ _1834_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__or3_1
X_4695_ net394 _0422_ _0117_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_3646_ _1768_ net147 _1801_ net151 cordic_inst.deg_handler_inst.theta_abs\[11\] VGND
+ VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a32o_1
X_3577_ cordic_inst.cordic_inst.x\[2\] cordic_inst.cordic_inst.cos_out\[2\] net211
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2528_ cordic_inst.cordic_inst.y\[19\] _0847_ _0851_ _0596_ VGND VGND VPWR VPWR _0863_
+ sky130_fd_sc_hd__o2bb2a_1
X_2459_ net243 _0692_ _0630_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4129_ net225 _2103_ cordic_inst.cordic_inst.cos_out\[12\] VGND VGND VPWR VPWR _2104_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3500_ net176 _1718_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__nor2_1
X_4480_ net326 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__inv_2
X_3431_ _1474_ _1669_ net174 VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__a21oi_1
X_3362_ _1596_ _1599_ _1600_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__o21ai_1
X_2313_ cordic_inst.cordic_inst.x\[29\] cordic_inst.cordic_inst.x\[30\] net307 VGND
+ VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux2_1
XFILLER_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3293_ _1515_ _1529_ _1530_ _1531_ _1526_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__o311a_1
XFILLER_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4816_ net400 _0543_ _0238_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_61_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4747_ net409 _0474_ _0169_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4678_ net407 _0405_ _0100_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3629_ cordic_inst.deg_handler_inst.theta_abs\[3\] _1759_ VGND VGND VPWR VPWR _1793_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput105 wstrb[2] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_1
XFILLER_29_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ axi_controller.write_addr_reg\[29\] net57 net188 VGND VGND VPWR VPWR _0328_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2931_ cordic_inst.cordic_inst.x\[29\] _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__nor2_1
XFILLER_43_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2862_ net216 _1120_ _1154_ _0713_ net281 VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a221o_1
X_4601_ net371 _0333_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_1
X_2793_ cordic_inst.cordic_inst.y\[15\] cordic_inst.cordic_inst.y\[16\] cordic_inst.cordic_inst.y\[17\]
+ cordic_inst.cordic_inst.y\[18\] net311 net301 VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux4_1
X_4532_ net376 _0264_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[14\] sky130_fd_sc_hd__dfxtp_1
X_4463_ net335 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__inv_2
X_3414_ cordic_inst.cordic_inst.z\[19\] _1636_ _1640_ cordic_inst.cordic_inst.z\[18\]
+ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__a22o_1
X_4394_ net341 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _1511_ _0707_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__nand2b_1
X_3276_ _1506_ _1514_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_56_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3130_ _1335_ _1337_ _1423_ net174 VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__a31o_1
XFILLER_79_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3061_ _1200_ _1363_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3963_ axi_controller.write_addr_reg\[12\] net39 net189 VGND VGND VPWR VPWR _0311_
+ sky130_fd_sc_hd__mux2_1
X_3894_ net75 _1965_ _1971_ net355 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__o211a_1
X_2914_ _1195_ _1198_ net271 VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__o21a_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2845_ _1138_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__and2_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4515_ net321 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__inv_2
X_2776_ cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.y\[29\] cordic_inst.cordic_inst.y\[30\]
+ net264 net305 net296 VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__mux4_2
X_4446_ net323 VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__inv_2
X_4377_ net330 VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
X_3328_ net274 _1481_ _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__mux2_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ net237 _0609_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__nor2_1
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2630_ cordic_inst.cordic_inst.y\[13\] _0932_ _0928_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2561_ cordic_inst.cordic_inst.y\[0\] _0718_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__nand2_1
X_2492_ _0800_ _0826_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__xnor2_1
X_4300_ net84 _2243_ _2249_ net351 VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o211a_1
X_4231_ _2192_ _2193_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__or2_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4162_ net224 _2132_ cordic_inst.cordic_inst.cos_out\[16\] VGND VGND VPWR VPWR _2133_
+ sky130_fd_sc_hd__a21oi_1
X_3113_ _1382_ _1397_ _1394_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__a21o_1
X_4093_ cordic_inst.cordic_inst.cos_out\[7\] _2068_ net226 VGND VGND VPWR VPWR _2072_
+ sky130_fd_sc_hd__o21a_1
X_3044_ cordic_inst.cordic_inst.x\[21\] _1345_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3946_ axi_controller.read_addr_reg\[17\] _1980_ _1988_ axi_controller.read_addr_reg\[2\]
+ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__or4b_1
X_3877_ axi_controller.write_addr_reg\[5\] _1959_ axi_controller.write_addr_reg\[3\]
+ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__or3b_1
X_2828_ net245 _1130_ _1124_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__o21ai_2
X_2759_ net184 _0901_ _1064_ net166 cordic_inst.cordic_inst.y\[2\] VGND VGND VPWR
+ VPWR _0532_ sky130_fd_sc_hd__a32o_1
XFILLER_78_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4429_ net344 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
Xfanout400 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_2
Xfanout411 net412 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3800_ _1880_ _1898_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__or2_1
X_4780_ net401 _0507_ _0202_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ cordic_inst.deg_handler_inst.theta_norm\[20\] cordic_inst.deg_handler_inst.theta_norm\[19\]
+ _1844_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__or3_1
XFILLER_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3662_ _1808_ _1809_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__nor2_1
X_3593_ cordic_inst.deg_handler_inst.theta_abs\[4\] _1760_ VGND VGND VPWR VPWR _1761_
+ sky130_fd_sc_hd__or2_1
X_2613_ _0940_ _0941_ _0947_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__or3_1
X_2544_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__inv_2
X_2475_ cordic_inst.cordic_inst.y\[30\] _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nand2_1
X_4214_ net317 _2177_ _2178_ _2174_ _2175_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__a32o_1
X_4145_ cordic_inst.cordic_inst.cos_out\[14\] _2117_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_87_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4076_ axi_controller.result_out\[5\] _2057_ net203 VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
X_3027_ _1287_ _1294_ _1318_ _1323_ _1293_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__a2111o_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3929_ axi_controller.read_addr_reg\[30\] net25 net195 VGND VGND VPWR VPWR _0296_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout230 _0612_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_2
Xfanout241 net242 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout263 net264 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_2
Xfanout252 _0604_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_2
Xfanout274 net276 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__buf_2
XFILLER_86_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout296 net297 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_2
Xfanout285 net290 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2260_ cordic_inst.cordic_inst.y\[10\] VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__inv_2
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4901_ net389 _0019_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4832_ net366 _0559_ _0254_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[29\] sky130_fd_sc_hd__dfrtp_4
X_4763_ net367 _0490_ _0185_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_3714_ cordic_inst.deg_handler_inst.theta_norm\[14\] _1836_ VGND VGND VPWR VPWR _0013_
+ sky130_fd_sc_hd__xnor2_1
X_4694_ net394 _0421_ _0116_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_3645_ cordic_inst.deg_handler_inst.theta_abs\[11\] _1767_ VGND VGND VPWR VPWR _1801_
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3576_ cordic_inst.cordic_inst.x\[3\] cordic_inst.cordic_inst.cos_out\[3\] net211
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_1
X_2527_ _0860_ _0861_ _0858_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__a21o_1
X_2458_ net278 _0749_ _0631_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2389_ net265 _0647_ _0648_ _0645_ net233 net231 VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__mux4_1
X_4128_ cordic_inst.cordic_inst.cos_out\[11\] cordic_inst.cordic_inst.cos_out\[10\]
+ _2089_ VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__or3_1
X_4059_ _2040_ _2042_ net229 VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__mux2_1
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap216 _0709_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
X_3430_ _1476_ _1477_ _1666_ _1668_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__o31ai_1
X_3361_ cordic_inst.cordic_inst.z\[2\] _1593_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_29_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2312_ cordic_inst.cordic_inst.x\[27\] cordic_inst.cordic_inst.x\[28\] net307 VGND
+ VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux2_1
X_3292_ _1518_ _1525_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__nand2_1
XFILLER_85_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4815_ net401 _0542_ _0237_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[12\] sky130_fd_sc_hd__dfrtp_2
X_4746_ net409 _0473_ _0168_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4677_ net407 _0404_ _0099_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3628_ _1759_ net147 _1792_ net152 cordic_inst.deg_handler_inst.theta_abs\[2\] VGND
+ VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a32o_1
X_3559_ cordic_inst.cordic_inst.x\[20\] cordic_inst.cordic_inst.cos_out\[20\] net209
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
Xinput106 wstrb[3] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2930_ _1226_ _1232_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4600_ net374 _0332_ VGND VGND VPWR VPWR axi_controller.mode sky130_fd_sc_hd__dfxtp_1
X_2861_ _1159_ _1160_ _1163_ net247 VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__o22a_1
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2792_ cordic_inst.cordic_inst.y\[11\] cordic_inst.cordic_inst.y\[12\] cordic_inst.cordic_inst.y\[13\]
+ cordic_inst.cordic_inst.y\[14\] net309 net299 VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux4_1
X_4531_ net380 _0263_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4462_ net342 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__inv_2
X_3413_ _1651_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__inv_2
X_4393_ net341 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ net294 _1509_ net206 net287 VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__a211o_1
XFILLER_85_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3275_ cordic_inst.cordic_inst.z\[12\] _1513_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__nand2_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4729_ net386 _0456_ _0151_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3060_ net252 _1201_ _1217_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__o21bai_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3962_ axi_controller.write_addr_reg\[11\] net38 net189 VGND VGND VPWR VPWR _0310_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3893_ axi_controller.reg_input_data\[13\] _1964_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__or2_1
X_2913_ net271 _1195_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2844_ net288 _1141_ _1145_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__a211o_1
X_4514_ net322 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__inv_2
X_2775_ cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.y\[29\] net305 VGND
+ VGND VPWR VPWR _1078_ sky130_fd_sc_hd__mux2_1
X_4445_ net324 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__inv_2
X_4376_ net332 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
X_3327_ _1564_ _1565_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _1485_ _1488_ _1484_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__o21ba_1
X_3189_ _1278_ _1464_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__and2_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2560_ cordic_inst.cordic_inst.y\[1\] _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__nand2_1
X_2491_ net169 _0652_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__nor2_1
X_4230_ cordic_inst.cordic_inst.sin_out\[24\] net257 _2191_ VGND VGND VPWR VPWR _2193_
+ sky130_fd_sc_hd__and3_1
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4161_ cordic_inst.cordic_inst.cos_out\[15\] cordic_inst.cordic_inst.cos_out\[14\]
+ cordic_inst.cordic_inst.cos_out\[13\] _2111_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__or4_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3112_ net179 _1401_ _1411_ net159 cordic_inst.cordic_inst.x\[28\] VGND VGND VPWR
+ VPWR _0526_ sky130_fd_sc_hd__a32o_1
X_4092_ net203 _2071_ _2064_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3043_ cordic_inst.cordic_inst.x\[21\] _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_66_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3945_ _0625_ _1982_ _1984_ _1985_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__or4_1
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3876_ _1955_ _1956_ _1957_ _1958_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__or4_1
X_2827_ net263 _1126_ _1128_ _1125_ net239 net232 VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux4_2
X_2758_ _0899_ _0900_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__or2_1
X_2689_ _0989_ _0990_ _1010_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a21o_1
X_4428_ net343 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__inv_2
Xfanout412 net413 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_2
Xfanout401 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__buf_2
XFILLER_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4359_ net347 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ cordic_inst.deg_handler_inst.theta_norm\[20\] _1846_ VGND VGND VPWR VPWR _0020_
+ sky130_fd_sc_hd__xnor2_1
X_3661_ cordic_inst.deg_handler_inst.theta_abs\[18\] cordic_inst.deg_handler_inst.theta_abs\[19\]
+ _1787_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__and3_1
XFILLER_9_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3592_ cordic_inst.deg_handler_inst.theta_abs\[3\] _1759_ VGND VGND VPWR VPWR _1760_
+ sky130_fd_sc_hd__or2_1
X_2612_ _0945_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__or2_1
X_2543_ cordic_inst.cordic_inst.y\[6\] _0875_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_10_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2474_ _0639_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__xnor2_1
X_4213_ cordic_inst.cordic_inst.sin_out\[22\] net258 _2176_ VGND VGND VPWR VPWR _2178_
+ sky130_fd_sc_hd__nand3_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4144_ cordic_inst.cordic_inst.cos_out\[13\] _2111_ net224 VGND VGND VPWR VPWR _2117_
+ sky130_fd_sc_hd__o21a_1
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4075_ net319 _2053_ _2055_ _2056_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__a22o_1
X_3026_ _1317_ _1321_ _1316_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__a21o_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3928_ axi_controller.read_addr_reg\[29\] net23 net195 VGND VGND VPWR VPWR _0295_
+ sky130_fd_sc_hd__mux2_1
X_3859_ _1932_ _1939_ _1941_ net107 net68 VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__o311a_1
XFILLER_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout220 _0680_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_2
Xfanout231 _0609_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_4
Xfanout242 _0607_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout264 cordic_inst.cordic_inst.y\[31\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_2
Xfanout253 cordic_inst.deg_handler_inst.theta_norm\[31\] VGND VGND VPWR VPWR net253
+ sky130_fd_sc_hd__buf_2
XFILLER_86_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout297 cordic_inst.cordic_inst.i\[1\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__buf_2
Xfanout286 net290 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
Xfanout275 net276 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_1
XFILLER_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4900_ net389 cordic_inst.deg_handler_inst.theta_norm\[0\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4831_ net366 _0558_ _0253_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4762_ net393 _0489_ _0184_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3713_ cordic_inst.deg_handler_inst.theta_norm\[13\] _1834_ net255 VGND VGND VPWR
+ VPWR _1836_ sky130_fd_sc_hd__o21ai_1
X_4693_ net396 _0420_ _0115_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_3644_ _1767_ net147 _1800_ net151 cordic_inst.deg_handler_inst.theta_abs\[10\] VGND
+ VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a32o_1
X_3575_ cordic_inst.cordic_inst.x\[4\] cordic_inst.cordic_inst.cos_out\[4\] net211
+ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux2_1
X_2526_ cordic_inst.cordic_inst.y\[17\] _0857_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nand2_1
X_2457_ _0631_ _0790_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__nand2_1
XFILLER_68_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2388_ net231 _0648_ _0633_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a21o_1
XFILLER_68_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4127_ net230 _2100_ _2101_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__or3_1
X_4058_ cordic_inst.cordic_inst.cos_out\[3\] _2041_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__xor2_1
XFILLER_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3009_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap206 _1502_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_1
Xmax_cap217 net218 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_1
X_3360_ _1597_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__nor2_1
X_2311_ cordic_inst.cordic_inst.x\[23\] cordic_inst.cordic_inst.x\[24\] cordic_inst.cordic_inst.x\[25\]
+ cordic_inst.cordic_inst.x\[26\] net306 net296 VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux4_1
X_3291_ cordic_inst.cordic_inst.z\[13\] _1505_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__nor2_1
XFILLER_38_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4814_ net400 _0541_ _0236_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[11\] sky130_fd_sc_hd__dfrtp_2
X_4745_ net408 _0472_ _0167_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4676_ net412 _0403_ _0098_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3627_ cordic_inst.deg_handler_inst.theta_abs\[2\] _1758_ VGND VGND VPWR VPWR _1792_
+ sky130_fd_sc_hd__nand2_1
X_3558_ cordic_inst.cordic_inst.x\[21\] cordic_inst.cordic_inst.cos_out\[21\] net209
+ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
X_2509_ _0832_ _0837_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__or3_1
XFILLER_88_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput107 wvalid VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
X_3489_ cordic_inst.cordic_inst.angle\[17\] net170 net163 cordic_inst.cordic_inst.z\[17\]
+ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__a22o_1
XFILLER_84_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2860_ _1161_ _1162_ net285 VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__mux2_1
X_2791_ _1084_ _1093_ net235 VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__mux2_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4530_ net381 _0262_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4461_ net342 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__inv_2
X_3412_ _1632_ _1647_ _1645_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__o21a_1
X_4392_ net348 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ net289 _1577_ _1580_ _1511_ _1522_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__o32a_1
X_3274_ net277 _1507_ _1512_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__mux2_1
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2989_ _1182_ _1291_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__xnor2_1
X_4728_ net385 _0455_ _0150_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[21\] sky130_fd_sc_hd__dfrtp_1
X_4659_ net406 _0389_ _0091_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_49_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3961_ axi_controller.write_addr_reg\[10\] net37 net189 VGND VGND VPWR VPWR _0309_
+ sky130_fd_sc_hd__mux2_1
X_2912_ net272 _1189_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__nand2_1
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3892_ net74 _1965_ _1970_ net352 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o211a_1
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2843_ cordic_inst.cordic_inst.y\[0\] net222 _0711_ _1143_ net220 VGND VGND VPWR
+ VPWR _1146_ sky130_fd_sc_hd__a32o_1
X_2774_ net246 _1076_ net215 VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__a21o_1
X_4513_ net323 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__inv_2
X_4444_ net324 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__inv_2
X_4375_ net331 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_84_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3326_ _1498_ _1558_ _0706_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__o21ai_1
XFILLER_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3257_ _1486_ _1490_ _1495_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__or3_1
X_3188_ _1260_ _1263_ _1277_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__nand3_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2490_ _0823_ _0824_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__and2_1
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4160_ cordic_inst.cordic_inst.sin_out\[16\] net259 _2128_ _2130_ VGND VGND VPWR
+ VPWR _2131_ sky130_fd_sc_hd__a31o_1
X_3111_ _1240_ _1396_ _1398_ _1400_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__or4_1
XFILLER_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4091_ net230 _2066_ _2067_ _2069_ _2070_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__o32a_1
X_3042_ _1207_ _1344_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3944_ axi_controller.read_addr_reg\[25\] _1981_ _1983_ _1986_ VGND VGND VPWR VPWR
+ _1987_ sky130_fd_sc_hd__nor4_1
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3875_ axi_controller.write_addr_reg\[17\] axi_controller.write_addr_reg\[16\] axi_controller.write_addr_reg\[19\]
+ axi_controller.write_addr_reg\[18\] VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__or4_1
X_2826_ net232 _1128_ _1071_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__a21o_1
X_2757_ net185 _0905_ _1063_ net166 cordic_inst.cordic_inst.y\[3\] VGND VGND VPWR
+ VPWR _0533_ sky130_fd_sc_hd__a32o_1
X_2688_ _0989_ _0990_ _1010_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__nand3_1
X_4427_ net343 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__inv_2
Xfanout413 net414 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_2
Xfanout402 net414 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_2
XFILLER_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4358_ net346 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
X_4289_ axi_controller.reg_input_data\[16\] _2242_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__or2_1
X_3309_ net293 _0706_ _0712_ net221 _0705_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__a311o_1
XFILLER_58_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ cordic_inst.deg_handler_inst.theta_abs\[18\] _1787_ cordic_inst.deg_handler_inst.theta_abs\[19\]
+ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__a21oi_2
X_3591_ cordic_inst.deg_handler_inst.theta_abs\[0\] cordic_inst.deg_handler_inst.theta_abs\[1\]
+ cordic_inst.deg_handler_inst.theta_abs\[2\] VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__or3_1
X_2611_ _0597_ _0944_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__and2_1
X_2542_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__inv_2
X_4212_ net258 _2176_ cordic_inst.cordic_inst.sin_out\[22\] VGND VGND VPWR VPWR _2177_
+ sky130_fd_sc_hd__a21o_1
X_2473_ net268 _0807_ _0806_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_79_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4143_ cordic_inst.cordic_inst.sin_out\[14\] _2115_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__xor2_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4074_ cordic_inst.cordic_inst.cos_out\[5\] _2054_ net319 VGND VGND VPWR VPWR _2056_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_87_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3025_ _1304_ _1307_ _1326_ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_34_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3927_ axi_controller.read_addr_reg\[28\] net22 net197 VGND VGND VPWR VPWR _0294_
+ sky130_fd_sc_hd__mux2_1
X_3858_ net47 net36 _1933_ _1940_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__or4_1
X_3789_ axi_controller.reg_input_data\[20\] axi_controller.reg_input_data\[19\] axi_controller.reg_input_data\[22\]
+ axi_controller.reg_input_data\[21\] VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__o211a_1
X_2809_ cordic_inst.cordic_inst.y\[26\] cordic_inst.cordic_inst.y\[27\] net305 VGND
+ VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux2_1
Xfanout221 _0678_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_2
Xfanout232 net234 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_4
Xfanout210 net214 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_4
Xfanout254 cordic_inst.deg_handler_inst.theta_norm\[31\] VGND VGND VPWR VPWR net254
+ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_6_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout243 net246 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_4
Xfanout265 net266 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_2
Xfanout287 net288 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_2
Xfanout298 net301 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_2
Xfanout276 net277 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_2
XFILLER_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ net367 _0557_ _0252_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4761_ net393 _0488_ _0183_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_3712_ cordic_inst.deg_handler_inst.theta_norm\[13\] _1835_ VGND VGND VPWR VPWR _0012_
+ sky130_fd_sc_hd__xnor2_1
X_4692_ net397 _0419_ _0114_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_3643_ cordic_inst.deg_handler_inst.theta_abs\[10\] _1766_ VGND VGND VPWR VPWR _1800_
+ sky130_fd_sc_hd__nand2_1
X_3574_ cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.cos_out\[5\] net211
+ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux2_1
X_2525_ cordic_inst.cordic_inst.y\[16\] _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__nand2_1
X_2456_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4126_ net261 _2099_ cordic_inst.cordic_inst.sin_out\[12\] VGND VGND VPWR VPWR _2101_
+ sky130_fd_sc_hd__a21oi_1
X_2387_ _0645_ _0647_ net297 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux2_1
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4057_ cordic_inst.cordic_inst.cos_out\[2\] cordic_inst.cordic_inst.cos_out\[1\]
+ cordic_inst.cordic_inst.cos_out\[0\] net227 VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__o31a_1
X_3008_ cordic_inst.cordic_inst.x\[12\] _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_82_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4959_ net411 _0588_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_1
XFILLER_10_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap218 _0708_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_1
X_3290_ _1528_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__inv_2
X_2310_ cordic_inst.cordic_inst.x\[25\] cordic_inst.cordic_inst.x\[26\] net307 VGND
+ VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4813_ net400 _0540_ _0235_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_61_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4744_ net407 _0471_ _0166_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4675_ net405 _0402_ _0097_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3626_ _1758_ _1790_ _1791_ net151 cordic_inst.deg_handler_inst.theta_abs\[1\] VGND
+ VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a32o_1
X_3557_ cordic_inst.cordic_inst.x\[22\] cordic_inst.cordic_inst.cos_out\[22\] net207
+ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
XFILLER_88_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2508_ _0841_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nand2_1
X_3488_ _1632_ _1648_ _1705_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__or3_1
X_2439_ net284 _0754_ _0637_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__o21a_1
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4109_ cordic_inst.cordic_inst.sin_out\[9\] cordic_inst.cordic_inst.sin_out\[8\]
+ cordic_inst.cordic_inst.sin_out\[7\] _2065_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__or4_1
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ cordic_inst.cordic_inst.y\[19\] cordic_inst.cordic_inst.y\[20\] cordic_inst.cordic_inst.y\[21\]
+ cordic_inst.cordic_inst.y\[22\] net308 net298 VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__mux4_1
X_4460_ net342 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__inv_2
X_4391_ net347 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
X_3411_ _1532_ _1628_ _1649_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__a21o_1
X_3342_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _1510_ _1511_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__nand2b_1
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2988_ _1180_ _1184_ net271 VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__o21ai_1
X_4727_ net385 _0454_ _0149_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[20\] sky130_fd_sc_hd__dfrtp_1
X_4658_ net406 _0388_ _0090_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[2\] sky130_fd_sc_hd__dfrtp_1
Xinput90 wdata[27] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
X_3609_ cordic_inst.deg_handler_inst.theta_abs\[28\] cordic_inst.deg_handler_inst.theta_abs\[29\]
+ cordic_inst.deg_handler_inst.theta_abs\[30\] cordic_inst.deg_handler_inst.theta_abs\[31\]
+ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__or4_1
XFILLER_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4589_ net360 _0321_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3960_ axi_controller.write_addr_reg\[9\] net67 net190 VGND VGND VPWR VPWR _0308_
+ sky130_fd_sc_hd__mux2_1
X_2911_ _1070_ _1092_ net280 VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__a21oi_1
X_3891_ axi_controller.reg_input_data\[12\] _1964_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_61_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2842_ cordic_inst.cordic_inst.y\[1\] net217 net216 _1144_ net281 VGND VGND VPWR
+ VPWR _1145_ sky130_fd_sc_hd__a221o_1
X_2773_ net238 _1075_ _1070_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__a21bo_1
X_4512_ net323 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__inv_2
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4443_ net329 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__inv_2
X_4374_ net331 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
X_3325_ net287 _0707_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__or2_1
X_3256_ _1491_ _1492_ _1494_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_69_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ cordic_inst.cordic_inst.x\[5\] net157 _1462_ _1463_ VGND VGND VPWR VPWR _0503_
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3110_ net179 _1409_ _1410_ net162 cordic_inst.cordic_inst.x\[29\] VGND VGND VPWR
+ VPWR _0527_ sky130_fd_sc_hd__a32o_1
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4090_ cordic_inst.cordic_inst.cos_out\[7\] net226 _2068_ net319 VGND VGND VPWR VPWR
+ _2070_ sky130_fd_sc_hd__a31o_1
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3041_ net252 _1208_ _1218_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_66_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3943_ axi_controller.read_addr_reg\[20\] axi_controller.read_addr_reg\[23\] axi_controller.read_addr_reg\[22\]
+ _1984_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__or4_1
X_3874_ axi_controller.write_addr_reg\[25\] axi_controller.write_addr_reg\[24\] axi_controller.write_addr_reg\[27\]
+ axi_controller.write_addr_reg\[26\] VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__or4_1
X_2825_ net231 _1086_ _1072_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__a21o_1
X_2756_ _0902_ _0904_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__or2_1
X_2687_ cordic_inst.cordic_inst.y\[26\] net158 _1015_ _1016_ VGND VGND VPWR VPWR _0556_
+ sky130_fd_sc_hd__a22o_1
X_4426_ net343 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__inv_2
Xfanout414 net1 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_4
Xfanout403 net404 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4357_ net339 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
XFILLER_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3308_ _1540_ _1546_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__nor2_1
X_4288_ net105 _1963_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__nand2_2
XFILLER_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3239_ net251 cordic_inst.cordic_inst.z\[24\] VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__nand2_1
XFILLER_27_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3590_ cordic_inst.deg_handler_inst.theta_abs\[0\] cordic_inst.deg_handler_inst.theta_abs\[1\]
+ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__or2_1
X_2610_ _0597_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__nor2_1
X_2541_ cordic_inst.cordic_inst.y\[6\] _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nor2_1
X_2472_ net278 _0774_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__nor2_1
X_4211_ cordic_inst.cordic_inst.sin_out\[21\] _2169_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__or2_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4142_ cordic_inst.cordic_inst.sin_out\[13\] _2107_ net260 VGND VGND VPWR VPWR _2115_
+ sky130_fd_sc_hd__o21a_1
X_4073_ cordic_inst.cordic_inst.cos_out\[5\] _2054_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__or2_1
X_3024_ _1298_ _1302_ _1297_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3926_ axi_controller.read_addr_reg\[27\] net21 net197 VGND VGND VPWR VPWR _0293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3857_ net39 net42 net41 _1934_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__or4_1
XFILLER_50_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2808_ cordic_inst.cordic_inst.y\[22\] cordic_inst.cordic_inst.y\[23\] cordic_inst.cordic_inst.y\[24\]
+ cordic_inst.cordic_inst.y\[25\] net306 net296 VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__mux4_1
X_3788_ axi_controller.reg_input_data\[22\] _1889_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__xnor2_1
X_2739_ net174 _1039_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nor2_1
XFILLER_59_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout200 net205 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout211 net212 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_4
Xfanout222 _0678_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_2
X_4409_ net340 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
Xfanout255 net256 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout244 net246 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_2
Xfanout233 net234 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_4
Xfanout266 net267 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__buf_1
Xfanout299 net300 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_2
Xfanout277 cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_2
Xfanout288 net289 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_2
XFILLER_27_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4760_ net393 _0487_ _0182_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3711_ net255 _1834_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__nand2_1
X_4691_ net396 _0418_ _0113_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3642_ _1766_ net147 _1799_ net151 cordic_inst.deg_handler_inst.theta_abs\[9\] VGND
+ VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3573_ cordic_inst.cordic_inst.x\[6\] cordic_inst.cordic_inst.cos_out\[6\] net211
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
X_2524_ _0785_ _0855_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__xor2_1
X_2455_ net247 _0755_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__nand2_1
X_2386_ _0719_ _0720_ net292 VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux2_1
X_4125_ cordic_inst.cordic_inst.sin_out\[12\] net261 _2099_ VGND VGND VPWR VPWR _2100_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4056_ cordic_inst.cordic_inst.sin_out\[3\] _2039_ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3007_ _1190_ _1215_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__xor2_1
XFILLER_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4958_ net410 _0587_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_1
X_4889_ net378 _0042_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_3909_ axi_controller.read_addr_reg\[10\] net3 net195 VGND VGND VPWR VPWR _0276_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4812_ net407 _0539_ _0234_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[9\] sky130_fd_sc_hd__dfrtp_2
X_4743_ net410 _0470_ _0165_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4674_ net385 _0401_ _0096_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.done sky130_fd_sc_hd__dfrtp_1
X_3625_ cordic_inst.deg_handler_inst.theta_abs\[0\] cordic_inst.deg_handler_inst.theta_abs\[1\]
+ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__nand2_1
X_3556_ cordic_inst.cordic_inst.x\[23\] cordic_inst.cordic_inst.cos_out\[23\] net207
+ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
X_2507_ cordic_inst.cordic_inst.y\[21\] _0840_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__or2_1
XFILLER_88_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3487_ _1632_ _1705_ _1648_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__o21ai_1
X_2438_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__inv_2
X_2369_ cordic_inst.cordic_inst.x\[4\] cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.x\[6\]
+ cordic_inst.cordic_inst.x\[7\] net312 net302 VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__mux4_1
X_4108_ axi_controller.result_out\[10\] net203 VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__nor2_1
X_4039_ axi_controller.reg_input_data\[7\] _2018_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__or2_1
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4390_ net348 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
X_3410_ _1647_ _1642_ _1634_ _1645_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__or4bb_1
X_3341_ net294 net304 net315 VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__and3_1
X_3272_ net294 net304 net289 VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2987_ _1244_ _1247_ _1282_ _1289_ _1243_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a311o_1
X_4726_ net385 _0453_ _0148_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[19\] sky130_fd_sc_hd__dfrtp_1
X_4657_ net405 _0387_ _0089_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[1\] sky130_fd_sc_hd__dfrtp_2
Xinput91 wdata[28] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
Xinput80 wdata[18] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
X_3608_ cordic_inst.deg_handler_inst.theta_abs\[19\] cordic_inst.deg_handler_inst.theta_abs\[20\]
+ _1775_ cordic_inst.deg_handler_inst.theta_abs\[21\] VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__a31o_1
XFILLER_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4588_ net360 _0320_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[21\] sky130_fd_sc_hd__dfxtp_1
X_3539_ _1596_ _1599_ _1600_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__or3_1
XFILLER_72_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2910_ net246 _1186_ net215 VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__a21o_1
X_3890_ net73 _1965_ _1969_ net355 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__o211a_1
XFILLER_31_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2841_ cordic_inst.cordic_inst.y\[2\] cordic_inst.cordic_inst.y\[3\] net314 VGND
+ VGND VPWR VPWR _1144_ sky130_fd_sc_hd__mux2_1
X_2772_ net232 _1074_ _1071_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__a21o_1
X_4511_ net323 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__inv_2
X_4442_ net329 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__inv_2
X_4373_ net331 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
X_3324_ _1561_ _1562_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__or2_1
X_3255_ net273 cordic_inst.cordic_inst.z\[23\] VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3186_ _1279_ _1280_ net177 VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__a21o_1
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4709_ net403 _0436_ _0131_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3040_ _1341_ _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3942_ axi_controller.read_addr_reg\[20\] axi_controller.read_addr_reg\[23\] axi_controller.read_addr_reg\[22\]
+ axi_controller.read_addr_reg\[25\] VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__or4_1
X_3873_ axi_controller.write_addr_reg\[28\] axi_controller.write_addr_reg\[29\] axi_controller.write_addr_reg\[30\]
+ axi_controller.write_addr_reg\[31\] VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__nand4_1
X_2824_ _1125_ _1126_ net291 VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__mux2_1
X_2755_ net185 _0909_ _1062_ net166 cordic_inst.cordic_inst.y\[4\] VGND VGND VPWR
+ VPWR _0534_ sky130_fd_sc_hd__a32o_1
X_2686_ net174 _1012_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__nor2_1
X_4425_ net346 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
Xfanout404 net405 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlymetal6s2s_1
X_4356_ net337 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3307_ _1544_ _1545_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__nand2b_1
XFILLER_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4287_ net105 _1963_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__and2_1
XFILLER_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3238_ net273 cordic_inst.cordic_inst.z\[28\] VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__xor2_1
XFILLER_27_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3169_ _1321_ _1441_ _1318_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__a21boi_1
XFILLER_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2540_ _0693_ _0870_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__xnor2_1
X_2471_ _0644_ _0805_ net268 VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__o21a_1
X_4210_ cordic_inst.cordic_inst.cos_out\[22\] _0613_ _2173_ net317 VGND VGND VPWR
+ VPWR _2175_ sky130_fd_sc_hd__a31oi_1
XFILLER_79_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4141_ axi_controller.result_out\[13\] _2114_ net202 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux2_1
XFILLER_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4072_ cordic_inst.cordic_inst.cos_out\[4\] _2048_ net226 VGND VGND VPWR VPWR _2054_
+ sky130_fd_sc_hd__o21a_1
XFILLER_83_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3023_ cordic_inst.cordic_inst.x\[13\] _1306_ _1310_ cordic_inst.cordic_inst.x\[12\]
+ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3925_ axi_controller.read_addr_reg\[26\] net20 net197 VGND VGND VPWR VPWR _0292_
+ sky130_fd_sc_hd__mux2_1
X_3856_ _1935_ _1936_ _1937_ _1938_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__or4b_1
X_3787_ axi_controller.reg_input_data\[21\] _1880_ _1883_ _1887_ VGND VGND VPWR VPWR
+ _1889_ sky130_fd_sc_hd__o31a_1
X_2807_ net285 _1106_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a21o_1
X_2738_ _0947_ _1038_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__nand2_1
X_4408_ net341 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
X_2669_ _0810_ _1000_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__a21oi_1
Xfanout223 _0613_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_2
Xfanout201 net202 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_2
Xfanout212 net213 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
Xfanout256 cordic_inst.deg_handler_inst.theta_norm\[31\] VGND VGND VPWR VPWR net256
+ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout245 net246 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_2
Xfanout234 net236 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4339_ net138 net193 net154 axi_controller.result_out\[4\] VGND VGND VPWR VPWR _0590_
+ sky130_fd_sc_hd__a22o_1
Xfanout278 net280 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_4
Xfanout267 cordic_inst.cordic_inst.x\[31\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__buf_2
Xfanout289 net290 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_2
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3710_ cordic_inst.deg_handler_inst.theta_norm\[12\] _1832_ VGND VGND VPWR VPWR _1834_
+ sky130_fd_sc_hd__or2_1
X_4690_ net396 _0417_ _0112_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3641_ cordic_inst.deg_handler_inst.theta_abs\[9\] _1765_ VGND VGND VPWR VPWR _1799_
+ sky130_fd_sc_hd__nand2_1
X_3572_ cordic_inst.cordic_inst.x\[7\] cordic_inst.cordic_inst.cos_out\[7\] net213
+ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux2_1
X_2523_ cordic_inst.cordic_inst.y\[17\] _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__nor2_1
X_2454_ _0771_ _0781_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__or3_1
X_2385_ cordic_inst.cordic_inst.x\[21\] cordic_inst.cordic_inst.x\[22\] cordic_inst.cordic_inst.x\[23\]
+ cordic_inst.cordic_inst.x\[24\] net306 net297 VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux4_1
X_4124_ cordic_inst.cordic_inst.sin_out\[11\] cordic_inst.cordic_inst.sin_out\[10\]
+ _2086_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__or3_1
Xinput1 aclk VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4055_ cordic_inst.cordic_inst.sin_out\[2\] cordic_inst.cordic_inst.sin_out\[1\]
+ cordic_inst.cordic_inst.sin_out\[0\] net262 VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__o31a_1
X_3006_ _1307_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4957_ net410 _0586_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_1
X_4888_ net378 _0041_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_3908_ axi_controller.read_addr_reg\[9\] net33 net196 VGND VGND VPWR VPWR _0275_
+ sky130_fd_sc_hd__mux2_1
X_3839_ _1924_ _1925_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__or2_1
XFILLER_10_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4811_ net407 _0538_ _0233_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[8\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_16_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4742_ net412 _0469_ _0164_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4673_ net374 _0400_ _0095_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.start sky130_fd_sc_hd__dfrtp_1
X_3624_ net148 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
X_3555_ cordic_inst.cordic_inst.x\[24\] cordic_inst.cordic_inst.cos_out\[24\] net207
+ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
X_2506_ cordic_inst.cordic_inst.y\[21\] _0840_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nand2_1
X_3486_ cordic_inst.cordic_inst.angle\[18\] net170 net164 cordic_inst.cordic_inst.z\[18\]
+ _1711_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__a221o_1
X_2437_ net265 _0642_ _0747_ _0744_ net240 net246 VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__mux4_2
XFILLER_69_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2368_ cordic_inst.cordic_inst.x\[4\] cordic_inst.cordic_inst.x\[5\] net312 VGND
+ VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux2_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2299_ net231 _0632_ _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__a21o_1
X_4107_ axi_controller.result_out\[9\] _2084_ net203 VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__mux2_1
X_4038_ net99 _2019_ _2026_ net354 VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__o211a_1
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3340_ net287 _1521_ _1578_ net220 _1500_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_90_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ net222 _0707_ _1509_ net220 VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__a22o_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2986_ _1287_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__nand2_1
X_4725_ net391 _0452_ _0147_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[18\] sky130_fd_sc_hd__dfrtp_1
X_4656_ net385 _0386_ _0088_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[0\] sky130_fd_sc_hd__dfrtp_1
Xinput70 rready VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
Xinput81 wdata[19] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
X_4587_ net360 _0319_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[20\] sky130_fd_sc_hd__dfxtp_1
X_3607_ _0615_ _1774_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__nand2_1
Xinput92 wdata[29] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
X_3538_ net176 _1602_ _1747_ _1748_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__o31ai_1
XFILLER_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3469_ cordic_inst.cordic_inst.angle\[22\] net171 net163 cordic_inst.cordic_inst.z\[22\]
+ _1698_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a221o_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2840_ cordic_inst.cordic_inst.y\[4\] cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.y\[6\]
+ cordic_inst.cordic_inst.y\[7\] net312 net302 VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__mux4_1
X_2771_ net231 _1073_ _1072_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__a21o_1
X_4510_ net325 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__inv_2
X_4441_ net329 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_44_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4372_ net331 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
X_3323_ cordic_inst.cordic_inst.z\[6\] _1560_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__nor2_1
XFILLER_39_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3254_ _1491_ _1492_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__or2_1
X_3185_ _1279_ _1280_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__nor2_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2969_ _1270_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__nand2b_1
X_4708_ net403 _0435_ _0130_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_62_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4639_ net398 _0370_ net331 VGND VGND VPWR VPWR axi_controller.result_out\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_80_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3941_ axi_controller.read_addr_reg\[24\] axi_controller.read_addr_reg\[27\] axi_controller.read_addr_reg\[26\]
+ axi_controller.read_addr_reg\[28\] VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__or4b_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3872_ axi_controller.write_addr_reg\[21\] axi_controller.write_addr_reg\[20\] axi_controller.write_addr_reg\[23\]
+ axi_controller.write_addr_reg\[22\] VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__or4_1
X_2823_ _1083_ _1085_ net296 VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__mux2_1
X_2754_ _0906_ _0907_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__or2_1
X_2685_ _0986_ _1011_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__or2_1
X_4424_ net347 VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__inv_2
Xfanout405 net413 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__buf_2
X_4355_ net339 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
X_3306_ cordic_inst.cordic_inst.z\[10\] _1543_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__or2_1
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4286_ _2240_ _2241_ axi_controller.result_out\[31\] net199 VGND VGND VPWR VPWR _0385_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3237_ _1475_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__inv_2
X_3168_ cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.next_state\[1\] _1451_
+ net175 VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__o22a_1
XFILLER_54_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3099_ _1236_ _1238_ _1401_ _1234_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__a31o_1
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ net268 _0798_ _0804_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a21o_1
XFILLER_55_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4140_ _2112_ _2113_ _2110_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4071_ cordic_inst.cordic_inst.sin_out\[5\] _2052_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3022_ _1290_ _1295_ _1313_ _1324_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__or4bb_1
XFILLER_63_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3924_ axi_controller.read_addr_reg\[25\] net19 net196 VGND VGND VPWR VPWR _0291_
+ sky130_fd_sc_hd__mux2_1
X_3855_ net56 net57 net59 net60 VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__and4_1
X_3786_ _1887_ _1888_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and2_1
X_2806_ net219 _1107_ _1108_ net221 net279 VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a221o_1
X_2737_ net181 _1050_ _1051_ net162 cordic_inst.cordic_inst.y\[11\] VGND VGND VPWR
+ VPWR _0541_ sky130_fd_sc_hd__a32o_1
X_2668_ _1001_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__xor2_1
XFILLER_59_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4407_ net339 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__inv_2
Xfanout213 net214 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
Xfanout202 net205 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__buf_2
X_2599_ cordic_inst.cordic_inst.y\[13\] _0932_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout224 net225 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_2
Xfanout246 net248 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
Xfanout235 net236 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4338_ net139 net193 net154 axi_controller.result_out\[5\] VGND VGND VPWR VPWR _0589_
+ sky130_fd_sc_hd__a22o_1
Xfanout257 net258 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_2
X_4269_ cordic_inst.cordic_inst.cos_out\[28\] net223 _2218_ cordic_inst.cordic_inst.cos_out\[29\]
+ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__a211o_1
Xfanout268 net270 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__buf_2
Xfanout279 net280 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_2
XFILLER_86_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _1765_ net147 _1798_ net151 cordic_inst.deg_handler_inst.theta_abs\[8\] VGND
+ VGND VPWR VPWR _0083_ sky130_fd_sc_hd__a32o_1
X_3571_ cordic_inst.cordic_inst.x\[8\] cordic_inst.cordic_inst.cos_out\[8\] net213
+ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
X_2522_ _0784_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2453_ _0665_ _0667_ _0786_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__or3b_1
X_2384_ cordic_inst.cordic_inst.x\[17\] cordic_inst.cordic_inst.x\[18\] cordic_inst.cordic_inst.x\[19\]
+ cordic_inst.cordic_inst.x\[20\] net308 net298 VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__mux4_1
X_4123_ axi_controller.result_out\[11\] _2098_ net203 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 araddr[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4054_ axi_controller.result_out\[2\] _2038_ net204 VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
X_3005_ cordic_inst.cordic_inst.x\[13\] _1306_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__nand2_1
X_4956_ net409 _0585_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_1
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4887_ net378 _0040_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_3907_ axi_controller.read_addr_reg\[8\] net32 net196 VGND VGND VPWR VPWR _0274_
+ sky130_fd_sc_hd__mux2_1
X_3838_ net145 axi_controller.state\[1\] net70 _1921_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__a31o_1
X_3769_ axi_controller.reg_input_data\[24\] _1873_ axi_controller.reg_input_data\[31\]
+ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__o21bai_2
XFILLER_3_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4810_ net406 _0537_ _0232_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[7\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_16_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ net412 _0468_ _0163_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4672_ net385 net157 _0094_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3623_ _1785_ _1789_ _1780_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__a21oi_2
X_3554_ cordic_inst.cordic_inst.x\[25\] cordic_inst.cordic_inst.cos_out\[25\] net207
+ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
X_2505_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__inv_2
X_3485_ _1706_ _1710_ net182 VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__and3b_1
XFILLER_88_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2436_ net153 _0758_ _0765_ _0769_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__nand4_2
XFILLER_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2367_ _0700_ _0701_ net292 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__mux2_1
X_2298_ net265 net297 VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__and2_1
X_4106_ _2083_ _2082_ _2080_ net229 VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__a2bb2o_1
X_4037_ axi_controller.reg_input_data\[6\] _2018_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__or2_1
XFILLER_37_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4939_ net365 _0568_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_1
XFILLER_20_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3270_ net303 net314 VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_90_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2985_ cordic_inst.cordic_inst.x\[8\] _1286_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__or2_1
X_4724_ net385 _0451_ _0146_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[17\] sky130_fd_sc_hd__dfrtp_1
X_4655_ net374 net205 net337 VGND VGND VPWR VPWR axi_controller.done sky130_fd_sc_hd__dfrtp_1
Xinput60 awaddr[31] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
Xinput71 wdata[0] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
Xinput82 wdata[1] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
X_3606_ cordic_inst.deg_handler_inst.theta_abs\[17\] _1773_ VGND VGND VPWR VPWR _1774_
+ sky130_fd_sc_hd__nand2_1
X_4586_ net361 _0318_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[19\] sky130_fd_sc_hd__dfxtp_1
Xinput93 wdata[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
X_3537_ cordic_inst.cordic_inst.angle\[3\] net172 net165 cordic_inst.cordic_inst.z\[3\]
+ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__a22oi_1
X_3468_ _1693_ _1697_ net182 VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__and3b_1
XFILLER_88_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2419_ net233 _0723_ _0635_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a21oi_1
X_3399_ cordic_inst.cordic_inst.z\[19\] _1636_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__nand2_1
XFILLER_17_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2770_ cordic_inst.cordic_inst.y\[30\] net264 net305 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__mux2_1
X_4440_ net330 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__inv_2
X_4371_ net334 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
X_3322_ cordic_inst.cordic_inst.z\[6\] _1560_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__and2_1
XFILLER_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3253_ net249 cordic_inst.cordic_inst.z\[22\] VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__nor2_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3184_ net184 _1461_ net157 cordic_inst.cordic_inst.x\[6\] VGND VGND VPWR VPWR _0504_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2968_ cordic_inst.cordic_inst.x\[1\] _1268_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__xor2_1
X_4707_ net404 _0434_ _0129_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[0\] sky130_fd_sc_hd__dfrtp_1
X_4638_ net398 _0369_ net332 VGND VGND VPWR VPWR axi_controller.result_out\[15\] sky130_fd_sc_hd__dfrtp_1
X_2899_ _1199_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nand2_1
X_4569_ net370 _0301_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3940_ _0625_ _1982_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__or2_1
XFILLER_51_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3871_ axi_controller.write_addr_reg\[12\] axi_controller.write_addr_reg\[15\] axi_controller.write_addr_reg\[14\]
+ _1951_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__or4_1
X_2822_ cordic_inst.cordic_inst.y\[21\] cordic_inst.cordic_inst.y\[22\] cordic_inst.cordic_inst.y\[23\]
+ cordic_inst.cordic_inst.y\[24\] net306 net296 VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__mux4_1
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2753_ cordic_inst.cordic_inst.y\[5\] net166 _1061_ net184 VGND VGND VPWR VPWR _0535_
+ sky130_fd_sc_hd__a22o_1
X_2684_ cordic_inst.cordic_inst.y\[27\] net158 _1014_ net178 VGND VGND VPWR VPWR _0557_
+ sky130_fd_sc_hd__a22o_1
X_4423_ net347 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__inv_2
X_4354_ net339 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
X_3305_ cordic_inst.cordic_inst.z\[10\] _1543_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__and2_1
Xfanout406 net413 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_2
X_4285_ net316 _2236_ _2237_ net199 VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__o31a_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3236_ net270 cordic_inst.cordic_inst.z\[29\] VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__xnor2_1
X_3167_ _1312_ _1442_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__xnor2_1
X_3098_ _1396_ _1398_ _1400_ _1240_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__o31ai_4
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4070_ cordic_inst.cordic_inst.sin_out\[4\] _2045_ net262 VGND VGND VPWR VPWR _2052_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_83_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3021_ _1318_ _1323_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__nor2_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3923_ axi_controller.read_addr_reg\[24\] net18 net197 VGND VGND VPWR VPWR _0290_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3854_ net53 net52 net55 net54 VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__or4_1
X_2805_ cordic_inst.cordic_inst.y\[6\] cordic_inst.cordic_inst.y\[7\] cordic_inst.cordic_inst.y\[8\]
+ cordic_inst.cordic_inst.y\[9\] net309 net300 VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__mux4_1
X_3785_ _1884_ _1885_ _1886_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__or3_1
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2736_ _0942_ _0945_ _1039_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__or3_1
X_2667_ net264 net267 VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__xnor2_2
X_4406_ net348 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
Xfanout214 _1472_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_4
X_2598_ cordic_inst.cordic_inst.y\[13\] _0932_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nor2_1
Xfanout203 net205 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_4
Xfanout225 net227 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
Xfanout247 net248 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_4
X_4337_ net140 net193 net154 axi_controller.result_out\[6\] VGND VGND VPWR VPWR _0588_
+ sky130_fd_sc_hd__a22o_1
X_4268_ cordic_inst.cordic_inst.cos_out\[28\] cordic_inst.cordic_inst.cos_out\[27\]
+ _2210_ net223 cordic_inst.cordic_inst.cos_out\[29\] VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__o311a_1
Xfanout258 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__buf_2
Xfanout269 net270 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3219_ cordic_inst.cordic_inst.y\[14\] cordic_inst.cordic_inst.sin_out\[14\] net214
+ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
XFILLER_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4199_ _2162_ _2165_ axi_controller.result_out\[20\] net202 VGND VGND VPWR VPWR _0374_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3570_ cordic_inst.cordic_inst.x\[9\] cordic_inst.cordic_inst.cos_out\[9\] net213
+ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
X_2521_ _0782_ _0785_ net252 VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a21o_1
X_2452_ _0782_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ net248 _0699_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__o21a_1
X_4122_ _2094_ _2095_ _2097_ net320 VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__o22ai_1
X_4053_ _2035_ _2037_ net229 VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__mux2_1
XFILLER_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput3 araddr[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_3004_ cordic_inst.cordic_inst.x\[13\] _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__or2_1
XFILLER_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4955_ net401 _0584_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_1
X_3906_ axi_controller.read_addr_reg\[7\] net31 net198 VGND VGND VPWR VPWR _0273_
+ sky130_fd_sc_hd__mux2_1
X_4886_ net378 axi_controller.reg_input_data\[18\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_3837_ net35 _1922_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__nor2_1
X_3768_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1871_
+ _1872_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__or4_1
X_2719_ _0955_ _1037_ _0962_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o21a_1
X_3699_ cordic_inst.deg_handler_inst.theta_norm\[8\] cordic_inst.deg_handler_inst.theta_norm\[7\]
+ _1824_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__or3_1
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4740_ net412 _0467_ _0162_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4671_ net385 cordic_inst.cordic_inst.next_state\[0\] _0093_ VGND VGND VPWR VPWR
+ cordic_inst.cordic_inst.state\[0\] sky130_fd_sc_hd__dfrtp_1
X_3622_ _1779_ _1783_ _1787_ _1788_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3553_ cordic_inst.cordic_inst.x\[26\] cordic_inst.cordic_inst.cos_out\[26\] net208
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux2_1
X_2504_ _0792_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__xnor2_1
X_3484_ _1648_ _1705_ _1651_ _1641_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__a211o_1
X_2435_ net153 _0758_ _0765_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__and4_1
XFILLER_84_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2366_ cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.x\[13\] cordic_inst.cordic_inst.x\[14\]
+ cordic_inst.cordic_inst.x\[15\] net309 net299 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux4_1
X_4105_ cordic_inst.cordic_inst.sin_out\[9\] net261 _2081_ net229 VGND VGND VPWR VPWR
+ _2083_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2297_ cordic_inst.cordic_inst.x\[30\] net265 net307 VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux2_1
X_4036_ net98 _2019_ _2025_ net354 VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o211a_1
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4938_ net366 _0567_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_1
X_4869_ net380 axi_controller.reg_input_data\[1\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2984_ cordic_inst.cordic_inst.x\[8\] _1286_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__nand2_1
X_4723_ net391 _0450_ _0145_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[16\] sky130_fd_sc_hd__dfrtp_1
X_4654_ net363 _0385_ net326 VGND VGND VPWR VPWR axi_controller.result_out\[31\] sky130_fd_sc_hd__dfrtp_1
Xinput72 wdata[10] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
Xinput50 awaddr[22] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
X_3605_ cordic_inst.deg_handler_inst.theta_abs\[16\] _1772_ VGND VGND VPWR VPWR _1773_
+ sky130_fd_sc_hd__or2_1
X_4585_ net361 _0317_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[18\] sky130_fd_sc_hd__dfxtp_1
Xinput61 awaddr[3] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
Xinput94 wdata[30] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
X_3536_ _1592_ _1594_ _1601_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__and3_1
Xinput83 wdata[20] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
X_3467_ _1493_ _1692_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__nand2_1
X_2418_ net285 _0751_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a21o_1
X_3398_ cordic_inst.cordic_inst.z\[19\] _1636_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__or2_1
XFILLER_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2349_ net280 _0651_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a21o_1
X_4019_ axi_controller.reg_input_data\[30\] _2008_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__or2_1
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4370_ net334 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
X_3321_ net274 _1504_ _1559_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__mux2_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3252_ net249 cordic_inst.cordic_inst.z\[22\] VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__and2_1
XFILLER_39_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3183_ _1249_ _1281_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2967_ _0603_ _1138_ _1147_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__and3_1
X_4706_ net363 _0433_ _0128_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_2898_ net244 _1137_ _1068_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__a21oi_2
X_4637_ net398 _0368_ net332 VGND VGND VPWR VPWR axi_controller.result_out\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4568_ net370 _0300_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_3519_ cordic_inst.cordic_inst.angle\[9\] net173 net167 cordic_inst.cordic_inst.z\[9\]
+ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__a22o_1
X_4499_ net335 VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__inv_2
XFILLER_57_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3870_ _1948_ _1950_ _1951_ _1952_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__or4_1
X_2821_ net285 _1119_ _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a21o_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2752_ _0910_ _0912_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__xor2_1
X_4422_ net346 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__inv_2
X_2683_ _0984_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__xnor2_1
X_4353_ net340 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
X_3304_ _1481_ net274 _1542_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__mux2_1
X_4284_ cordic_inst.cordic_inst.sin_out\[31\] _2238_ _2239_ VGND VGND VPWR VPWR _2240_
+ sky130_fd_sc_hd__o21ai_1
Xfanout407 net411 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_2
X_3235_ net273 cordic_inst.cordic_inst.z\[30\] VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__xnor2_1
X_3166_ cordic_inst.cordic_inst.x\[13\] net160 _1450_ net180 VGND VGND VPWR VPWR _0511_
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3097_ cordic_inst.cordic_inst.x\[27\] _1384_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__a21o_1
X_3999_ net108 _0610_ _1924_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3020_ _1321_ _1322_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nand2_1
XFILLER_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3922_ axi_controller.read_addr_reg\[23\] net17 net197 VGND VGND VPWR VPWR _0289_
+ sky130_fd_sc_hd__mux2_1
X_3853_ net44 net43 net46 net45 VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__or4_1
X_2804_ cordic_inst.cordic_inst.y\[10\] cordic_inst.cordic_inst.y\[11\] cordic_inst.cordic_inst.y\[12\]
+ cordic_inst.cordic_inst.y\[13\] net309 net299 VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__mux4_1
X_3784_ axi_controller.reg_input_data\[21\] _1886_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__nand2_1
X_2735_ _0945_ _1039_ _0942_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__o21ai_1
X_2666_ _0639_ _0806_ _0807_ net268 VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__o31a_1
X_4405_ net341 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__inv_2
X_2597_ _0778_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__xnor2_1
X_4336_ net141 net194 _2256_ axi_controller.result_out\[7\] VGND VGND VPWR VPWR _0587_
+ sky130_fd_sc_hd__a22o_1
Xfanout204 net205 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
Xfanout237 _0608_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
Xfanout215 _1068_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_2
Xfanout226 net227 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_2
X_4267_ cordic_inst.cordic_inst.sin_out\[29\] net258 _2221_ VGND VGND VPWR VPWR _2225_
+ sky130_fd_sc_hd__nand3_1
Xfanout259 net260 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__buf_2
Xfanout248 _0606_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_2
X_4198_ net318 _2164_ net202 VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__o21a_1
X_3218_ cordic_inst.cordic_inst.y\[15\] cordic_inst.cordic_inst.sin_out\[15\] net210
+ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_1
X_3149_ cordic_inst.cordic_inst.x\[17\] net161 _1437_ net180 VGND VGND VPWR VPWR _0515_
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2520_ net252 _0782_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__or2_1
XFILLER_60_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2451_ _0783_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2382_ net288 _0702_ _0715_ _0716_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__a211o_1
X_4121_ cordic_inst.cordic_inst.cos_out\[11\] _2096_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__xnor2_1
X_4052_ cordic_inst.cordic_inst.cos_out\[2\] _2036_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__xor2_1
Xinput4 araddr[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_3003_ _1192_ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4954_ net400 _0583_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_1
X_3905_ axi_controller.read_addr_reg\[6\] net30 net198 VGND VGND VPWR VPWR _0272_
+ sky130_fd_sc_hd__mux2_1
X_4885_ net378 axi_controller.reg_input_data\[17\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3836_ net68 net35 VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__nor2_1
X_3767_ axi_controller.reg_input_data\[30\] axi_controller.reg_input_data\[29\] axi_controller.reg_input_data\[28\]
+ axi_controller.reg_input_data\[27\] VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__or4_1
X_2718_ _0915_ _0959_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__or2_1
X_3698_ cordic_inst.deg_handler_inst.theta_norm\[8\] _1826_ VGND VGND VPWR VPWR _0038_
+ sky130_fd_sc_hd__xnor2_1
X_2649_ _0982_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__and2b_1
X_4319_ net128 net191 net156 axi_controller.result_out\[24\] VGND VGND VPWR VPWR _0570_
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4670_ net371 _0399_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
X_3621_ _0615_ cordic_inst.deg_handler_inst.theta_abs\[19\] cordic_inst.deg_handler_inst.theta_abs\[22\]
+ cordic_inst.deg_handler_inst.theta_abs\[23\] VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__or4b_1
X_3552_ cordic_inst.cordic_inst.x\[27\] cordic_inst.cordic_inst.cos_out\[27\] net208
+ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
X_2503_ _0789_ _0793_ net269 VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__o21a_1
X_3483_ cordic_inst.cordic_inst.angle\[19\] net170 net164 cordic_inst.cordic_inst.z\[19\]
+ _1709_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a221o_1
X_2434_ net278 _0766_ _0767_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a22o_1
X_2365_ cordic_inst.cordic_inst.x\[8\] cordic_inst.cordic_inst.x\[9\] cordic_inst.cordic_inst.x\[10\]
+ cordic_inst.cordic_inst.x\[11\] net309 net299 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__mux4_1
X_4104_ net261 _2081_ cordic_inst.cordic_inst.sin_out\[9\] VGND VGND VPWR VPWR _2082_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2296_ net267 net278 VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nand2_2
X_4035_ axi_controller.reg_input_data\[5\] _2018_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__or2_1
XFILLER_52_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4937_ net365 _0566_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_1
XFILLER_52_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4868_ net380 axi_controller.reg_input_data\[0\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3819_ _1912_ _1910_ axi_controller.reg_input_data\[29\] VGND VGND VPWR VPWR _1913_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4799_ net369 _0526_ _0221_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2983_ _1184_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__xor2_1
X_4722_ net391 _0449_ _0144_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4653_ net359 _0384_ net321 VGND VGND VPWR VPWR axi_controller.result_out\[30\] sky130_fd_sc_hd__dfrtp_1
Xinput40 awaddr[13] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput73 wdata[11] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
X_3604_ cordic_inst.deg_handler_inst.theta_abs\[15\] _1771_ VGND VGND VPWR VPWR _1772_
+ sky130_fd_sc_hd__or2_1
Xinput51 awaddr[23] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
X_4584_ net361 _0316_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[17\] sky130_fd_sc_hd__dfxtp_1
Xinput62 awaddr[4] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
Xinput95 wdata[31] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
X_3535_ net185 _1605_ _1745_ _1746_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a31o_1
Xinput84 wdata[21] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
X_3466_ net182 _1694_ _1695_ _1696_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a31o_1
XFILLER_88_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2417_ net219 _0726_ _0730_ net221 net281 VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a221o_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3397_ net277 _1635_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__xnor2_1
X_2348_ net283 _0669_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2279_ cordic_inst.deg_handler_inst.theta_abs\[18\] VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__inv_2
XFILLER_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4018_ net92 _2009_ _2015_ net352 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o211a_1
XFILLER_25_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3320_ net220 _1557_ _1558_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_13_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3251_ _1488_ _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__nand2_1
XFILLER_78_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3182_ _1459_ _1460_ cordic_inst.cordic_inst.x\[7\] net166 VGND VGND VPWR VPWR _0505_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2966_ cordic_inst.cordic_inst.x\[1\] _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__nand2_1
X_2897_ _1069_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4705_ net364 _0432_ _0127_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_4636_ net399 _0367_ net334 VGND VGND VPWR VPWR axi_controller.result_out\[13\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_31_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4567_ net370 _0299_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3518_ _1616_ _1619_ _1622_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__o21ai_1
X_4498_ net335 VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__inv_2
X_3449_ net182 _1682_ _1683_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2820_ net221 _1121_ _1122_ net219 net281 VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__a221o_1
X_2751_ net184 _1057_ _1060_ net166 cordic_inst.cordic_inst.y\[6\] VGND VGND VPWR
+ VPWR _0536_ sky130_fd_sc_hd__a32o_1
X_2682_ cordic_inst.cordic_inst.y\[26\] _0985_ _1012_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a21oi_1
X_4421_ net339 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__inv_2
X_4352_ net340 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
X_3303_ net221 _0706_ _0712_ _1541_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__and4b_1
X_4283_ cordic_inst.cordic_inst.sin_out\[31\] _2238_ net228 VGND VGND VPWR VPWR _2239_
+ sky130_fd_sc_hd__a21oi_1
Xfanout408 net411 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_1
X_3234_ net249 cordic_inst.cordic_inst.z\[30\] VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__nand2_1
X_3165_ _1309_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3096_ cordic_inst.cordic_inst.x\[27\] _1384_ _1387_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_37_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3998_ _0611_ _2002_ _2004_ _0621_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a211oi_1
XFILLER_10_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2949_ _0602_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__and2_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4619_ net381 _0350_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3921_ axi_controller.read_addr_reg\[22\] net16 net197 VGND VGND VPWR VPWR _0288_
+ sky130_fd_sc_hd__mux2_1
X_3852_ net49 net48 net51 net50 VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__or4_1
X_2803_ _1104_ _1105_ net292 VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux2_1
X_3783_ axi_controller.reg_input_data\[20\] axi_controller.reg_input_data\[19\] _1874_
+ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_42_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2734_ net181 _1041_ _1049_ net162 cordic_inst.cordic_inst.y\[12\] VGND VGND VPWR
+ VPWR _0542_ sky130_fd_sc_hd__a32o_1
X_2665_ _0819_ _0997_ _0812_ _0815_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__a211o_1
X_4404_ net341 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__inv_2
X_2596_ _0770_ _0773_ net252 VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a21o_1
Xfanout205 cordic_inst.sign_handler_inst.done_pulse VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_4
X_4335_ net142 net193 net154 axi_controller.result_out\[8\] VGND VGND VPWR VPWR _0586_
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout238 net239 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_2
Xfanout227 _0613_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4266_ net257 _2221_ cordic_inst.cordic_inst.sin_out\[29\] VGND VGND VPWR VPWR _2224_
+ sky130_fd_sc_hd__a21o_1
Xfanout249 net251 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_2
X_3217_ cordic_inst.cordic_inst.y\[16\] cordic_inst.cordic_inst.sin_out\[16\] net210
+ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
X_4197_ cordic_inst.cordic_inst.cos_out\[20\] _2163_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__xnor2_1
X_3148_ _1367_ _1436_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ _1377_ _1381_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__nand2_1
XFILLER_42_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2450_ net244 _0699_ _0630_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a21oi_1
X_2381_ cordic_inst.cordic_inst.x\[0\] net222 _0711_ _0704_ _0680_ VGND VGND VPWR
+ VPWR _0716_ sky130_fd_sc_hd__a32o_1
XFILLER_68_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4120_ cordic_inst.cordic_inst.cos_out\[10\] _2089_ net224 VGND VGND VPWR VPWR _2096_
+ sky130_fd_sc_hd__o21a_1
X_4051_ cordic_inst.cordic_inst.cos_out\[1\] cordic_inst.cordic_inst.cos_out\[0\]
+ net227 VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__o21a_1
Xinput5 araddr[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_3002_ _1189_ _1190_ net272 VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__o21a_1
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4953_ net401 _0582_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3904_ axi_controller.read_addr_reg\[5\] net29 net196 VGND VGND VPWR VPWR _0271_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4884_ net378 axi_controller.reg_input_data\[16\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3835_ _0610_ net68 VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__or2_1
X_3766_ axi_controller.reg_input_data\[22\] _1870_ axi_controller.reg_input_data\[23\]
+ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__o21a_1
X_2717_ net180 _0972_ _1036_ net160 cordic_inst.cordic_inst.y\[16\] VGND VGND VPWR
+ VPWR _0546_ sky130_fd_sc_hd__a32o_1
X_3697_ cordic_inst.deg_handler_inst.theta_norm\[7\] _1824_ net255 VGND VGND VPWR
+ VPWR _1826_ sky130_fd_sc_hd__o21ai_1
X_2648_ cordic_inst.cordic_inst.y\[27\] _0981_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__nand2_1
X_2579_ cordic_inst.cordic_inst.y\[7\] _0872_ _0879_ _0913_ _0877_ VGND VGND VPWR
+ VPWR _0914_ sky130_fd_sc_hd__o221a_1
X_4318_ net129 net191 net156 axi_controller.result_out\[25\] VGND VGND VPWR VPWR _0569_
+ sky130_fd_sc_hd__a22o_1
X_4249_ axi_controller.result_out\[26\] _2209_ net199 VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux2_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3620_ cordic_inst.deg_handler_inst.theta_abs\[17\] _1773_ VGND VGND VPWR VPWR _1787_
+ sky130_fd_sc_hd__or2_2
X_3551_ cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.cos_out\[28\] net208
+ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
X_2502_ _0835_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nand2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3482_ _1639_ _1707_ _1708_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__o21a_1
X_2433_ net242 _0739_ net279 VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__a21oi_1
X_2364_ _0696_ _0698_ net284 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__mux2_2
X_4103_ cordic_inst.cordic_inst.sin_out\[8\] _2075_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_87_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2295_ _0601_ net243 VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__nor2_1
X_4034_ net97 _2019_ _2024_ net354 VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o211a_1
XFILLER_52_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4936_ net365 _0565_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_1
X_4867_ net383 _0077_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[31\] sky130_fd_sc_hd__dfxtp_1
X_3818_ _1911_ _1912_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_50_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4798_ net363 _0525_ _0220_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[27\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3749_ cordic_inst.deg_handler_inst.theta_norm\[27\] _1858_ VGND VGND VPWR VPWR _0027_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_79_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2982_ net272 _1180_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__nand2_1
X_4721_ net391 _0448_ _0143_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_61_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4652_ net359 _0383_ net321 VGND VGND VPWR VPWR axi_controller.result_out\[29\] sky130_fd_sc_hd__dfrtp_1
X_3603_ cordic_inst.deg_handler_inst.theta_abs\[14\] _1770_ VGND VGND VPWR VPWR _1771_
+ sky130_fd_sc_hd__or2_1
Xinput30 araddr[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput52 awaddr[24] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
X_4583_ net361 _0315_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[16\] sky130_fd_sc_hd__dfxtp_1
Xinput41 awaddr[14] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput63 awaddr[5] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
Xinput96 wdata[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput74 wdata[12] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
X_3534_ cordic_inst.cordic_inst.angle\[4\] net172 net165 cordic_inst.cordic_inst.z\[4\]
+ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__a22o_1
Xinput85 wdata[22] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
X_3465_ cordic_inst.cordic_inst.angle\[23\] net171 net163 cordic_inst.cordic_inst.z\[23\]
+ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__a22o_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2416_ _0719_ _0727_ net235 VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__mux2_1
X_3396_ net289 _1576_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__nor2_1
XFILLER_29_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2347_ net221 _0679_ net219 _0681_ net279 VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a221o_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2278_ cordic_inst.cordic_inst.state\[1\] VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__inv_2
X_4017_ axi_controller.reg_input_data\[29\] _2008_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__or2_1
XFILLER_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4919_ net379 _0018_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3250_ cordic_inst.cordic_inst.z\[20\] _1487_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__or2_1
X_3181_ _1247_ _1282_ _1283_ net177 VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__a31o_1
XFILLER_78_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4704_ net363 _0431_ _0126_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2965_ _1157_ _1267_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__xnor2_1
X_2896_ net244 _1151_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4635_ net399 _0366_ net334 VGND VGND VPWR VPWR axi_controller.result_out\[12\] sky130_fd_sc_hd__dfrtp_1
X_4566_ net374 _0298_ VGND VGND VPWR VPWR axi_controller.reg_done_flag sky130_fd_sc_hd__dfxtp_1
X_3517_ _1616_ _1619_ _1622_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__or3_1
X_4497_ net335 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_2
X_3448_ cordic_inst.cordic_inst.angle\[27\] net170 net163 cordic_inst.cordic_inst.z\[27\]
+ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__a22o_1
X_3379_ _1616_ _1617_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2750_ _0877_ _0878_ _0913_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__a21o_1
X_2681_ _0986_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__and2_1
XFILLER_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4420_ net337 VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__inv_2
X_4351_ net339 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
X_3302_ net287 net293 VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__nand2_1
X_4282_ cordic_inst.cordic_inst.sin_out\[30\] _2224_ net258 VGND VGND VPWR VPWR _2238_
+ sky130_fd_sc_hd__o21a_1
Xfanout409 net410 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_2
X_3233_ cordic_inst.cordic_inst.y\[0\] cordic_inst.cordic_inst.sin_out\[0\] net212
+ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
X_3164_ cordic_inst.cordic_inst.x\[12\] _1310_ _1443_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__a21oi_1
X_3095_ _1394_ _1397_ _1385_ _1389_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_65_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3997_ _1961_ _1995_ _2003_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__a21oi_1
X_2948_ _1131_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__xor2_1
X_4618_ net380 _0349_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[3\] sky130_fd_sc_hd__dfxtp_1
X_2879_ net263 _1149_ _1150_ _1152_ net245 net241 VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__mux4_1
X_4549_ net358 _0281_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3920_ axi_controller.read_addr_reg\[21\] net15 net195 VGND VGND VPWR VPWR _0287_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3851_ net66 net38 net37 net40 VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__or4_1
X_3782_ _1880_ _1883_ axi_controller.reg_input_data\[21\] VGND VGND VPWR VPWR _1885_
+ sky130_fd_sc_hd__o21a_1
X_2802_ cordic_inst.cordic_inst.y\[18\] cordic_inst.cordic_inst.y\[19\] cordic_inst.cordic_inst.y\[20\]
+ cordic_inst.cordic_inst.y\[21\] net308 net298 VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_42_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2733_ _0930_ _1040_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__or2_1
X_2664_ _0819_ _0997_ _0815_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a21o_1
X_4403_ net341 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__inv_2
X_2595_ _0928_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nor2_1
X_4334_ net143 net193 net154 axi_controller.result_out\[9\] VGND VGND VPWR VPWR _0585_
+ sky130_fd_sc_hd__a22o_1
Xfanout228 net230 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4265_ axi_controller.result_out\[28\] _2223_ net199 VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
Xfanout239 net240 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_2
X_3216_ cordic_inst.cordic_inst.y\[17\] cordic_inst.cordic_inst.sin_out\[17\] net209
+ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
X_4196_ cordic_inst.cordic_inst.cos_out\[19\] _2155_ net225 VGND VGND VPWR VPWR _2163_
+ sky130_fd_sc_hd__o21a_1
X_3147_ cordic_inst.cordic_inst.x\[16\] _1360_ _1361_ _1332_ VGND VGND VPWR VPWR _1436_
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3078_ _1379_ _1380_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__nor2_1
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2380_ cordic_inst.cordic_inst.x\[1\] net218 _0709_ _0710_ net281 VGND VGND VPWR
+ VPWR _0715_ sky130_fd_sc_hd__a221o_1
X_4050_ cordic_inst.cordic_inst.sin_out\[2\] _2034_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 araddr[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_3001_ _1299_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__and2_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4952_ net399 _0581_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_64_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4883_ net379 axi_controller.reg_input_data\[15\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3903_ axi_controller.read_addr_reg\[4\] net28 net198 VGND VGND VPWR VPWR _0270_
+ sky130_fd_sc_hd__mux2_1
X_3834_ net111 axi_controller.state\[2\] net69 _0621_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__a31o_1
X_3765_ axi_controller.reg_input_data\[19\] _1869_ axi_controller.reg_input_data\[21\]
+ axi_controller.reg_input_data\[20\] VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__o211a_1
X_3696_ cordic_inst.deg_handler_inst.theta_norm\[7\] _1825_ VGND VGND VPWR VPWR _0037_
+ sky130_fd_sc_hd__xnor2_1
X_2716_ _0968_ _0970_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__nand2_1
X_2647_ cordic_inst.cordic_inst.y\[27\] _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nor2_1
X_2578_ _0906_ _0907_ _0912_ _0911_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__a31o_1
X_4317_ net130 net191 net156 axi_controller.result_out\[26\] VGND VGND VPWR VPWR _0568_
+ sky130_fd_sc_hd__a22o_1
X_4248_ net316 _2208_ _2206_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__a21o_1
XFILLER_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4179_ net224 _2147_ cordic_inst.cordic_inst.cos_out\[18\] VGND VGND VPWR VPWR _2148_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3550_ cordic_inst.cordic_inst.x\[29\] cordic_inst.cordic_inst.cos_out\[29\] net214
+ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
X_2501_ cordic_inst.cordic_inst.y\[20\] _0834_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__or2_1
X_3481_ _1639_ _1707_ net176 VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__a21oi_1
X_2432_ net283 _0661_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2363_ _0641_ _0697_ net233 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__mux2_1
X_4102_ cordic_inst.cordic_inst.cos_out\[9\] _2079_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__xor2_1
X_4033_ axi_controller.reg_input_data\[4\] _2018_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__or2_1
X_2294_ net164 VGND VGND VPWR VPWR cordic_inst.cordic_inst.next_state\[1\] sky130_fd_sc_hd__inv_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4935_ net365 _0564_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_1
X_4866_ net383 _0076_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[30\] sky130_fd_sc_hd__dfxtp_1
X_3817_ axi_controller.reg_input_data\[28\] axi_controller.reg_input_data\[27\] _1908_
+ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__nor3_1
X_4797_ net363 _0524_ _0219_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[26\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_50_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3748_ net253 _1857_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__nand2_1
X_3679_ cordic_inst.deg_handler_inst.theta_abs\[30\] net149 VGND VGND VPWR VPWR _0076_
+ sky130_fd_sc_hd__and2_1
Xoutput140 net140 VGND VGND VPWR VPWR rdata[6] sky130_fd_sc_hd__buf_2
XFILLER_75_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2981_ _1244_ _1247_ _1282_ _1243_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__a31o_1
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4720_ net391 _0447_ _0142_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[13\] sky130_fd_sc_hd__dfrtp_1
X_4651_ net359 _0382_ net321 VGND VGND VPWR VPWR axi_controller.result_out\[28\] sky130_fd_sc_hd__dfrtp_1
X_3602_ cordic_inst.deg_handler_inst.theta_abs\[13\] _1769_ VGND VGND VPWR VPWR _1770_
+ sky130_fd_sc_hd__or2_1
Xinput20 araddr[26] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 araddr[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput53 awaddr[25] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput42 awaddr[15] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
X_4582_ net361 _0314_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[15\] sky130_fd_sc_hd__dfxtp_1
Xinput64 awaddr[6] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xinput75 wdata[13] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
Xinput97 wdata[4] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
X_3533_ _1591_ _1602_ _1604_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__or3_1
Xinput86 wdata[23] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
X_3464_ _1491_ _1494_ _1693_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__or3_1
X_2415_ _0746_ _0749_ net281 VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__mux2_2
X_3395_ _1632_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__nor2_1
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2346_ cordic_inst.cordic_inst.x\[11\] cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.x\[13\]
+ cordic_inst.cordic_inst.x\[14\] net309 net299 VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux4_1
XFILLER_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2277_ cordic_inst.deg_handler_inst.kuadran\[0\] VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__inv_2
X_4016_ net91 _2009_ _2014_ net352 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o211a_1
XFILLER_84_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4918_ net387 _0017_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_40_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4849_ net391 _0057_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3180_ _1247_ _1282_ _1283_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2964_ net275 _1138_ _1147_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__and3_1
X_4703_ net363 _0430_ _0125_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2895_ net244 _1196_ _1197_ net215 VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_32_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4634_ net400 _0365_ net335 VGND VGND VPWR VPWR axi_controller.result_out\[11\] sky130_fd_sc_hd__dfrtp_1
X_4565_ net357 _0297_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3516_ cordic_inst.cordic_inst.angle\[10\] net172 net167 cordic_inst.cordic_inst.z\[10\]
+ _1733_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4496_ net335 VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__inv_2
XFILLER_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3447_ _1660_ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__xnor2_1
X_3378_ cordic_inst.cordic_inst.z\[8\] _1615_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__nor2_1
X_2329_ net283 _0661_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_68_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2680_ _0979_ _0993_ _0989_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__o21a_1
XFILLER_12_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4350_ net346 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
X_3301_ _1538_ _1539_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__nand2_1
X_4281_ cordic_inst.cordic_inst.cos_out\[30\] _2227_ net223 cordic_inst.cordic_inst.cos_out\[31\]
+ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__o211a_1
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3232_ cordic_inst.cordic_inst.y\[1\] cordic_inst.cordic_inst.sin_out\[1\] net211
+ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
X_3163_ net181 _1445_ _1448_ net161 cordic_inst.cordic_inst.x\[14\] VGND VGND VPWR
+ VPWR _0512_ sky130_fd_sc_hd__a32o_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3094_ _1379_ _1393_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3996_ _0624_ _1942_ _1998_ _2002_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__a31o_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947_ net250 _1178_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__or2_1
X_4617_ net380 _0348_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_2878_ net238 _1150_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__nand2_1
XFILLER_89_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4548_ net358 _0280_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[14\] sky130_fd_sc_hd__dfxtp_1
X_4479_ net326 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__inv_2
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3850_ net58 net65 net64 net67 VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__or4_1
X_3781_ axi_controller.reg_input_data\[21\] _1880_ _1883_ VGND VGND VPWR VPWR _1884_
+ sky130_fd_sc_hd__nor3_1
X_2801_ cordic_inst.cordic_inst.y\[14\] cordic_inst.cordic_inst.y\[15\] cordic_inst.cordic_inst.y\[16\]
+ cordic_inst.cordic_inst.y\[17\] net311 net301 VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__mux4_1
X_2732_ cordic_inst.cordic_inst.y\[13\] net161 _1048_ net181 VGND VGND VPWR VPWR _0543_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2663_ _0815_ _0818_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__and2b_1
X_4402_ net341 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__inv_2
X_2594_ cordic_inst.cordic_inst.y\[12\] _0927_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__and2b_1
X_4333_ net113 net193 net154 axi_controller.result_out\[10\] VGND VGND VPWR VPWR _0584_
+ sky130_fd_sc_hd__a22o_1
X_4264_ net316 _2219_ _2222_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__o21ai_1
Xfanout207 net208 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_4
Xfanout229 net230 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_2
XFILLER_59_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3215_ cordic_inst.cordic_inst.y\[18\] cordic_inst.cordic_inst.sin_out\[18\] net209
+ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
X_4195_ cordic_inst.cordic_inst.sin_out\[20\] net259 _2159_ _2161_ VGND VGND VPWR
+ VPWR _2162_ sky130_fd_sc_hd__a31o_1
X_3146_ net180 _1432_ _1435_ net161 cordic_inst.cordic_inst.x\[18\] VGND VGND VPWR
+ VPWR _0516_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_19_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3077_ cordic_inst.cordic_inst.x\[24\] _1378_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__nor2_1
XFILLER_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3979_ axi_controller.write_addr_reg\[28\] net56 net187 VGND VGND VPWR VPWR _0327_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 araddr[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_3000_ cordic_inst.cordic_inst.x\[14\] _1301_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__xor2_1
XFILLER_76_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4951_ net402 _0580_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_1
X_4882_ net379 axi_controller.reg_input_data\[14\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3902_ axi_controller.read_addr_reg\[3\] net27 net196 VGND VGND VPWR VPWR _0269_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3833_ net111 net69 VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__nand2_1
X_3764_ axi_controller.reg_input_data\[17\] axi_controller.reg_input_data\[16\] _1868_
+ axi_controller.reg_input_data\[18\] VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__o31a_1
X_3695_ net256 _1824_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__nand2_1
X_2715_ cordic_inst.cordic_inst.y\[17\] net160 _1035_ net180 VGND VGND VPWR VPWR _0547_
+ sky130_fd_sc_hd__a22o_1
X_2646_ _0804_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2577_ _0883_ _0885_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__nor2_1
X_4316_ net131 net191 net156 axi_controller.result_out\[27\] VGND VGND VPWR VPWR _0567_
+ sky130_fd_sc_hd__a22o_1
X_4247_ cordic_inst.cordic_inst.sin_out\[26\] _2207_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__xnor2_1
X_4178_ cordic_inst.cordic_inst.cos_out\[17\] cordic_inst.cordic_inst.cos_out\[16\]
+ _2132_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_2_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3129_ _1337_ _1423_ _1335_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2500_ cordic_inst.cordic_inst.y\[20\] _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__nand2_1
X_3480_ cordic_inst.cordic_inst.z\[18\] _1640_ _1706_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__a21o_1
X_2431_ net283 _0662_ _0637_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__o21a_1
X_2362_ cordic_inst.cordic_inst.x\[24\] cordic_inst.cordic_inst.x\[25\] cordic_inst.cordic_inst.x\[26\]
+ cordic_inst.cordic_inst.x\[27\] net305 net296 VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux4_1
X_4101_ cordic_inst.cordic_inst.cos_out\[8\] cordic_inst.cordic_inst.cos_out\[7\]
+ _2068_ net226 VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__o31a_1
X_2293_ net182 net170 VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__nor2_1
X_4032_ net96 _2019_ _2023_ net354 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__o211a_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4934_ net363 _0563_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4865_ net383 _0074_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[29\] sky130_fd_sc_hd__dfxtp_1
X_3816_ axi_controller.reg_input_data\[29\] _1910_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__xnor2_1
X_4796_ net369 _0523_ _0218_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[25\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3747_ cordic_inst.deg_handler_inst.theta_norm\[26\] cordic_inst.deg_handler_inst.theta_norm\[25\]
+ _1854_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__or3_1
X_3678_ cordic_inst.deg_handler_inst.theta_abs\[29\] net149 VGND VGND VPWR VPWR _0074_
+ sky130_fd_sc_hd__and2_1
Xoutput130 net130 VGND VGND VPWR VPWR rdata[26] sky130_fd_sc_hd__buf_2
X_2629_ _0939_ _0963_ _0962_ _0948_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__o2bb2a_1
Xoutput141 net141 VGND VGND VPWR VPWR rdata[7] sky130_fd_sc_hd__buf_2
XFILLER_75_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout390 net391 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2980_ _1243_ _1244_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__nand2b_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4650_ net365 _0381_ net321 VGND VGND VPWR VPWR axi_controller.result_out\[27\] sky130_fd_sc_hd__dfrtp_1
X_3601_ cordic_inst.deg_handler_inst.theta_abs\[12\] _1768_ VGND VGND VPWR VPWR _1769_
+ sky130_fd_sc_hd__or2_1
Xinput10 araddr[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 araddr[27] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput54 awaddr[26] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
Xinput32 araddr[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 awaddr[16] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
X_4581_ net361 _0313_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[14\] sky130_fd_sc_hd__dfxtp_1
Xinput98 wdata[5] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
Xinput76 wdata[14] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xinput87 wdata[24] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
X_3532_ cordic_inst.cordic_inst.angle\[5\] net172 net167 cordic_inst.cordic_inst.z\[5\]
+ _1744_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__a221o_1
Xinput65 awaddr[7] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
X_3463_ _1491_ _1693_ _1494_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__o21ai_1
XFILLER_88_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2414_ net283 _0747_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__o21ai_2
X_3394_ cordic_inst.cordic_inst.z\[16\] _1631_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__and2b_1
XFILLER_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2345_ net288 net293 VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__and2b_1
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2276_ net337 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
X_4015_ axi_controller.reg_input_data\[28\] _2008_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4917_ net387 _0016_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4848_ net390 _0056_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4779_ net407 _0506_ _0201_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2963_ cordic_inst.cordic_inst.x\[2\] _1265_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__nand2_1
X_4702_ net363 _0429_ _0124_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2894_ net241 _1088_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__or2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ net400 _0364_ net335 VGND VGND VPWR VPWR axi_controller.result_out\[10\] sky130_fd_sc_hd__dfrtp_1
X_4564_ net356 _0296_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[30\] sky130_fd_sc_hd__dfxtp_1
X_3515_ net177 _1732_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__nor2_1
XFILLER_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4495_ net345 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__inv_2
X_3446_ net249 cordic_inst.cordic_inst.z\[26\] _1680_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__a21boi_1
X_3377_ cordic_inst.cordic_inst.z\[8\] _1615_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__and2_1
X_2328_ net234 _0649_ _0635_ net238 VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_68_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2259_ cordic_inst.cordic_inst.y\[18\] VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__inv_2
XFILLER_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3300_ cordic_inst.cordic_inst.z\[11\] _1537_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__nand2_1
X_4280_ cordic_inst.deg_handler_inst.kuadran\[0\] _2232_ cordic_inst.cordic_inst.cos_out\[31\]
+ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__o21ba_1
XFILLER_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3231_ cordic_inst.cordic_inst.y\[2\] cordic_inst.cordic_inst.sin_out\[2\] net212
+ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
X_3162_ _1303_ _1444_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__or2_1
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3093_ _1382_ _1385_ _1389_ _1395_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__and4b_1
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3995_ net107 _0624_ _1943_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__o21ai_1
X_2946_ _1247_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__nand2_1
X_2877_ _1170_ _1179_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__or2_1
X_4616_ net381 _0347_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[1\] sky130_fd_sc_hd__dfxtp_1
X_4547_ net358 _0279_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4478_ net326 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__inv_2
X_3429_ cordic_inst.cordic_inst.z\[29\] cordic_inst.cordic_inst.z\[28\] net249 VGND
+ VGND VPWR VPWR _1668_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3780_ axi_controller.reg_input_data\[20\] axi_controller.reg_input_data\[19\] VGND
+ VGND VPWR VPWR _1883_ sky130_fd_sc_hd__and2_1
X_2800_ net279 _1089_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a21o_1
X_2731_ _0935_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_42_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4401_ net346 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__inv_2
X_2662_ _0983_ _0992_ _0994_ _0995_ _0821_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a41o_1
X_2593_ _0927_ cordic_inst.cordic_inst.y\[12\] VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__and2b_1
X_4332_ net114 net193 net154 axi_controller.result_out\[11\] VGND VGND VPWR VPWR _0583_
+ sky130_fd_sc_hd__a22o_1
X_4263_ net228 _2220_ _2221_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__or3b_1
Xfanout208 net214 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_4
Xfanout219 net220 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_2
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3214_ cordic_inst.cordic_inst.y\[19\] cordic_inst.cordic_inst.sin_out\[19\] net209
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
X_4194_ net318 _2160_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__nand2_1
XFILLER_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3145_ _1358_ _1431_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__nand2_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3076_ cordic_inst.cordic_inst.x\[24\] _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__and2_1
XFILLER_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3978_ axi_controller.write_addr_reg\[27\] net55 net187 VGND VGND VPWR VPWR _0326_
+ sky130_fd_sc_hd__mux2_1
X_2929_ net215 _1227_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__or2_1
XFILLER_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput8 araddr[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4950_ net398 _0579_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_1
X_4881_ net380 axi_controller.reg_input_data\[13\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3901_ axi_controller.read_addr_reg\[2\] net24 net196 VGND VGND VPWR VPWR _0268_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3832_ _0620_ _1919_ _1918_ cordic_inst.state\[0\] VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3763_ _1864_ _1865_ _1866_ _1867_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__or4_1
X_3694_ cordic_inst.deg_handler_inst.theta_norm\[6\] _1822_ VGND VGND VPWR VPWR _1824_
+ sky130_fd_sc_hd__or2_1
X_2714_ _0868_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__xor2_1
X_2645_ net169 _0798_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__nor2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4315_ net132 net191 net156 axi_controller.result_out\[28\] VGND VGND VPWR VPWR _0566_
+ sky130_fd_sc_hd__a22o_1
X_2576_ cordic_inst.cordic_inst.y\[4\] _0884_ _0886_ _0885_ VGND VGND VPWR VPWR _0911_
+ sky130_fd_sc_hd__a31o_1
X_4246_ cordic_inst.cordic_inst.sin_out\[25\] _2199_ net257 VGND VGND VPWR VPWR _2207_
+ sky130_fd_sc_hd__o21ai_1
X_4177_ cordic_inst.cordic_inst.sin_out\[18\] net259 _2143_ _2145_ VGND VGND VPWR
+ VPWR _2146_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_2_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3128_ _1339_ _1422_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__or2_1
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3059_ cordic_inst.cordic_inst.x\[16\] _1360_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2430_ _0677_ _0763_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nor2_1
X_2361_ _0694_ _0695_ net292 VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux2_1
X_2292_ _0614_ cordic_inst.cordic_inst.state\[0\] VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__and2_1
X_4100_ axi_controller.result_out\[8\] net203 _2078_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__o21ba_1
X_4031_ axi_controller.reg_input_data\[3\] _2018_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__or2_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4933_ net374 axi_controller.done _0257_ VGND VGND VPWR VPWR cordic_inst.done_d sky130_fd_sc_hd__dfrtp_1
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4864_ net383 _0073_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[28\] sky130_fd_sc_hd__dfxtp_1
X_3815_ _1877_ _1900_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__and2_1
X_4795_ net369 _0522_ _0217_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[24\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3746_ cordic_inst.deg_handler_inst.theta_norm\[26\] _1856_ VGND VGND VPWR VPWR _0026_
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_65_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3677_ cordic_inst.deg_handler_inst.theta_abs\[28\] net149 VGND VGND VPWR VPWR _0073_
+ sky130_fd_sc_hd__and2_1
Xoutput120 net120 VGND VGND VPWR VPWR rdata[17] sky130_fd_sc_hd__buf_2
Xoutput131 net131 VGND VGND VPWR VPWR rdata[27] sky130_fd_sc_hd__buf_2
X_2628_ _0941_ _0945_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__or2_1
Xoutput142 net142 VGND VGND VPWR VPWR rdata[8] sky130_fd_sc_hd__buf_2
X_2559_ _0735_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__xor2_1
XFILLER_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4229_ net257 _2191_ cordic_inst.cordic_inst.sin_out\[24\] VGND VGND VPWR VPWR _2192_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_75_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_83_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout380 net381 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_2
Xfanout391 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_2
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3600_ cordic_inst.deg_handler_inst.theta_abs\[11\] _1767_ VGND VGND VPWR VPWR _1768_
+ sky130_fd_sc_hd__or2_1
Xinput22 araddr[28] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 araddr[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_4580_ net370 _0312_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[13\] sky130_fd_sc_hd__dfxtp_1
X_3531_ net176 _1606_ _1743_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__nor3_1
Xinput33 araddr[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput55 awaddr[27] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xinput44 awaddr[17] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput77 wdata[15] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
Xinput88 wdata[25] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
Xinput66 awaddr[8] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput99 wdata[6] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3462_ _1493_ _1692_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__nor2_1
X_3393_ _1631_ cordic_inst.cordic_inst.z\[16\] VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__and2b_1
X_2413_ net234 _0641_ _0635_ net240 VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a211o_1
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2344_ cordic_inst.cordic_inst.x\[7\] cordic_inst.cordic_inst.x\[8\] cordic_inst.cordic_inst.x\[9\]
+ cordic_inst.cordic_inst.x\[10\] net309 net299 VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux4_1
X_2275_ net319 VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__inv_2
X_4014_ net90 _2009_ _2013_ net352 VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o211a_1
XFILLER_25_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4916_ net387 _0015_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4847_ net404 _0055_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[11\] sky130_fd_sc_hd__dfxtp_1
X_4778_ net407 _0505_ _0200_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[7\] sky130_fd_sc_hd__dfrtp_2
X_3729_ cordic_inst.deg_handler_inst.theta_norm\[19\] _1844_ net254 VGND VGND VPWR
+ VPWR _1846_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2962_ _1164_ _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__xnor2_1
X_4701_ net363 _0428_ _0123_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2893_ net285 _1099_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__or2_1
XFILLER_30_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4632_ net409 _0363_ net342 VGND VGND VPWR VPWR axi_controller.result_out\[9\] sky130_fd_sc_hd__dfrtp_1
X_4563_ net357 _0295_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[29\] sky130_fd_sc_hd__dfxtp_1
X_3514_ _1546_ _1623_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__xor2_1
X_4494_ net345 VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__inv_2
XFILLER_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3445_ _1663_ _1679_ _1661_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__o21ai_1
X_3376_ net275 _1614_ _1613_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__mux2_1
XFILLER_69_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2327_ net232 _0649_ _0635_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2258_ cordic_inst.cordic_inst.y\[28\] VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3230_ cordic_inst.cordic_inst.y\[3\] cordic_inst.cordic_inst.sin_out\[3\] net212
+ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
XFILLER_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3161_ cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.next_state\[1\] _1446_
+ _1447_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o22a_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3092_ _1393_ _1394_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3994_ _0610_ net145 _0619_ net350 _1928_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a41o_1
X_2945_ cordic_inst.cordic_inst.x\[6\] _1246_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__nand2b_1
X_2876_ _1103_ _1116_ _1131_ _1177_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__nand4_1
X_4615_ net381 _0346_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[0\] sky130_fd_sc_hd__dfxtp_1
X_4546_ net356 _0278_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[12\] sky130_fd_sc_hd__dfxtp_1
X_4477_ net325 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__inv_2
X_3428_ _1477_ _1666_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__nor2_1
X_3359_ cordic_inst.cordic_inst.z\[1\] _1595_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2730_ _0928_ _1041_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_42_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2661_ _0983_ _0992_ _0994_ _0995_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__and4_1
X_4400_ net346 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2592_ _0772_ _0921_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4331_ net115 net192 net155 axi_controller.result_out\[12\] VGND VGND VPWR VPWR _0582_
+ sky130_fd_sc_hd__a22o_1
X_4262_ net257 _2214_ cordic_inst.cordic_inst.sin_out\[28\] VGND VGND VPWR VPWR _2221_
+ sky130_fd_sc_hd__a21o_1
Xfanout209 net210 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_4
X_3213_ cordic_inst.cordic_inst.y\[20\] cordic_inst.cordic_inst.sin_out\[20\] net209
+ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_4193_ net259 _2159_ cordic_inst.cordic_inst.sin_out\[20\] VGND VGND VPWR VPWR _2160_
+ sky130_fd_sc_hd__a21o_1
XFILLER_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3144_ _1433_ _1434_ cordic_inst.cordic_inst.x\[19\] net161 VGND VGND VPWR VPWR _0517_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3075_ _1211_ _1221_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3977_ axi_controller.write_addr_reg\[26\] net54 net187 VGND VGND VPWR VPWR _0325_
+ sky130_fd_sc_hd__mux2_1
X_2928_ cordic_inst.cordic_inst.x\[30\] _1229_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__xor2_1
X_2859_ net264 _1073_ _1078_ _1112_ net231 net232 VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__mux4_2
XFILLER_40_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4529_ net388 _0261_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 araddr[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ net380 axi_controller.reg_input_data\[12\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3900_ axi_controller.read_addr_reg\[1\] net13 net198 VGND VGND VPWR VPWR _0267_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3831_ cordic_inst.state\[1\] _1919_ cordic_inst.state\[2\] VGND VGND VPWR VPWR _0007_
+ sky130_fd_sc_hd__a21o_1
X_3762_ axi_controller.reg_input_data\[7\] axi_controller.reg_input_data\[6\] axi_controller.reg_input_data\[5\]
+ axi_controller.reg_input_data\[4\] VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__or4_1
XFILLER_20_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3693_ cordic_inst.deg_handler_inst.theta_norm\[6\] _1823_ VGND VGND VPWR VPWR _0036_
+ sky130_fd_sc_hd__xnor2_1
X_2713_ _0860_ _0972_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__nand2_1
X_2644_ _0974_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2575_ cordic_inst.cordic_inst.y\[4\] _0886_ _0908_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a21o_1
X_4314_ net133 net191 net156 axi_controller.result_out\[29\] VGND VGND VPWR VPWR _0565_
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4245_ _0605_ cordic_inst.deg_handler_inst.kuadran\[0\] _2203_ _2205_ VGND VGND VPWR
+ VPWR _2206_ sky130_fd_sc_hd__o31a_1
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4176_ net319 _2144_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3127_ _1369_ _1421_ _1346_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__a21o_1
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3058_ cordic_inst.cordic_inst.x\[16\] _1360_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__xor2_1
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2360_ cordic_inst.cordic_inst.x\[20\] cordic_inst.cordic_inst.x\[21\] cordic_inst.cordic_inst.x\[22\]
+ cordic_inst.cordic_inst.x\[23\] net306 net297 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux4_1
X_2291_ _0614_ cordic_inst.cordic_inst.state\[0\] VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or2_2
X_4030_ net93 _2019_ _2022_ net354 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4932_ net375 _0562_ VGND VGND VPWR VPWR axi_controller.start_pulse_reg sky130_fd_sc_hd__dfxtp_1
X_4863_ net383 _0072_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[27\] sky130_fd_sc_hd__dfxtp_1
X_3814_ axi_controller.reg_input_data\[28\] _1909_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__xnor2_1
X_4794_ net402 _0521_ _0216_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[23\] sky130_fd_sc_hd__dfrtp_4
X_3745_ cordic_inst.deg_handler_inst.theta_norm\[25\] _1854_ net253 VGND VGND VPWR
+ VPWR _1856_ sky130_fd_sc_hd__o21ai_1
Xoutput110 net110 VGND VGND VPWR VPWR bresp[1] sky130_fd_sc_hd__buf_2
X_3676_ cordic_inst.deg_handler_inst.theta_abs\[27\] net149 VGND VGND VPWR VPWR _0072_
+ sky130_fd_sc_hd__and2_1
Xoutput132 net132 VGND VGND VPWR VPWR rdata[28] sky130_fd_sc_hd__buf_2
Xoutput121 net121 VGND VGND VPWR VPWR rdata[18] sky130_fd_sc_hd__buf_2
X_2627_ _0953_ _0957_ _0952_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__o21a_1
Xoutput143 net143 VGND VGND VPWR VPWR rdata[9] sky130_fd_sc_hd__buf_2
X_2558_ net248 _0699_ _0717_ net276 VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__o211a_1
X_2489_ cordic_inst.cordic_inst.y\[22\] _0822_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__or2_1
X_4228_ cordic_inst.cordic_inst.sin_out\[23\] cordic_inst.cordic_inst.sin_out\[22\]
+ _2176_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__or3_1
XFILLER_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4159_ net318 _2129_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__nand2_1
XFILLER_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout392 net414 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_2
Xfanout381 net382 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_2
Xfanout370 net372 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 araddr[19] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput34 aresetn VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_1
X_3530_ _1570_ _1575_ _1605_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__and3b_1
Xinput23 araddr[29] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput45 awaddr[18] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput89 wdata[26] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
Xinput56 awaddr[28] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 wdata[16] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
Xinput67 awaddr[9] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3461_ _1486_ _1691_ _1497_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__o21a_1
X_3392_ _1507_ net274 _1630_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__mux2_1
X_2412_ _0695_ _0697_ net291 VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__mux2_1
X_2343_ net288 net294 VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__nor2_1
X_4013_ axi_controller.reg_input_data\[27\] _2008_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__or2_1
X_2274_ net110 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__inv_2
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4915_ net387 _0014_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4846_ net404 _0054_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4777_ net407 _0504_ _0199_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[6\] sky130_fd_sc_hd__dfrtp_2
X_3728_ cordic_inst.deg_handler_inst.theta_norm\[19\] _1845_ VGND VGND VPWR VPWR _0018_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3659_ cordic_inst.deg_handler_inst.theta_abs\[18\] net150 net148 _1807_ VGND VGND
+ VPWR VPWR _0062_ sky130_fd_sc_hd__a22o_1
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2961_ _1148_ _1157_ net276 VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__o21a_1
X_4700_ net365 _0427_ _0122_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2892_ _1170_ _1179_ _1188_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__or4_2
X_4631_ net409 _0362_ net342 VGND VGND VPWR VPWR axi_controller.result_out\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4562_ net359 _0294_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[28\] sky130_fd_sc_hd__dfxtp_1
X_3513_ cordic_inst.cordic_inst.angle\[11\] net172 net167 cordic_inst.cordic_inst.z\[11\]
+ _1731_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a221o_1
X_4493_ net345 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__inv_2
X_3444_ _1658_ _1659_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__nor2_1
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3375_ net275 _0712_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__nand2_1
X_2326_ _0646_ _0660_ net232 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4829_ net367 _0556_ _0251_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[26\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_31_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3160_ _1299_ _1302_ _1445_ net175 VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__a31o_1
X_3091_ cordic_inst.cordic_inst.x\[25\] _1392_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3993_ net351 _2001_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and2_1
XFILLER_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2944_ _1246_ cordic_inst.cordic_inst.x\[6\] VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__nand2b_1
X_2875_ _1170_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__and2b_1
X_4614_ net369 _0005_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.kuadran\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_4545_ net356 _0277_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[11\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap153 _0743_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
X_4476_ net325 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3427_ _1658_ _1659_ _1662_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__o31a_1
X_3358_ _1583_ _1584_ cordic_inst.cordic_inst.z\[0\] VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__a21oi_1
X_2309_ net243 _0643_ net169 VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__a21o_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3289_ _1520_ _1527_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__nor2_1
XFILLER_57_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2660_ _0982_ _0985_ cordic_inst.cordic_inst.y\[26\] VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__nand3b_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2591_ _0920_ _0925_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__or2_1
XFILLER_5_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4330_ net116 net192 net155 axi_controller.result_out\[13\] VGND VGND VPWR VPWR _0581_
+ sky130_fd_sc_hd__a22o_1
X_4261_ cordic_inst.cordic_inst.sin_out\[28\] net257 _2214_ VGND VGND VPWR VPWR _2220_
+ sky130_fd_sc_hd__and3_1
X_3212_ cordic_inst.cordic_inst.y\[21\] cordic_inst.cordic_inst.sin_out\[21\] net209
+ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux2_1
X_4192_ cordic_inst.cordic_inst.sin_out\[19\] _2151_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__or2_1
XFILLER_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3143_ _1355_ _1357_ _1432_ net175 VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__a31o_1
XFILLER_27_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3074_ _1332_ _1368_ _1376_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__a21bo_1
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3976_ axi_controller.write_addr_reg\[25\] net53 net187 VGND VGND VPWR VPWR _0324_
+ sky130_fd_sc_hd__mux2_1
X_2927_ _1229_ cordic_inst.cordic_inst.x\[30\] VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and2b_1
X_2858_ _1105_ _1111_ net291 VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__mux2_1
X_2789_ net238 _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__nand2_1
X_4528_ net388 _0260_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4459_ net342 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__inv_2
XFILLER_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3830_ cordic_inst.done_d axi_controller.done VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__nand2b_1
X_3761_ axi_controller.reg_input_data\[3\] axi_controller.reg_input_data\[2\] axi_controller.reg_input_data\[1\]
+ axi_controller.reg_input_data\[0\] VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__or4_1
XFILLER_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2712_ net180 _1030_ _1033_ net160 cordic_inst.cordic_inst.y\[18\] VGND VGND VPWR
+ VPWR _0548_ sky130_fd_sc_hd__a32o_1
X_3692_ net256 _1822_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__nand2_1
X_2643_ _0976_ _0977_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_10_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2574_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__inv_2
X_4313_ net135 net191 net156 axi_controller.result_out\[30\] VGND VGND VPWR VPWR _0564_
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4244_ net316 _2204_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__nor2_1
X_4175_ net260 _2143_ cordic_inst.cordic_inst.sin_out\[18\] VGND VGND VPWR VPWR _2144_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3126_ _1375_ _1420_ _1343_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__a21o_1
X_3057_ _1201_ _1217_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__xor2_2
XFILLER_23_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3959_ axi_controller.write_addr_reg\[8\] net66 net189 VGND VGND VPWR VPWR _0307_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2290_ _0614_ cordic_inst.cordic_inst.state\[0\] VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__nor2_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4931_ net374 _0032_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4862_ net384 _0071_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[26\] sky130_fd_sc_hd__dfxtp_1
X_3813_ _1908_ _1906_ axi_controller.reg_input_data\[27\] VGND VGND VPWR VPWR _1909_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4793_ net368 _0520_ _0215_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[22\] sky130_fd_sc_hd__dfrtp_4
XFILLER_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3744_ cordic_inst.deg_handler_inst.theta_norm\[25\] _1855_ VGND VGND VPWR VPWR _0025_
+ sky130_fd_sc_hd__xnor2_1
X_3675_ cordic_inst.deg_handler_inst.theta_abs\[26\] net149 VGND VGND VPWR VPWR _0071_
+ sky130_fd_sc_hd__and2_1
X_2626_ _0915_ _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__or2_1
Xoutput111 net111 VGND VGND VPWR VPWR bvalid sky130_fd_sc_hd__buf_2
Xoutput133 net133 VGND VGND VPWR VPWR rdata[29] sky130_fd_sc_hd__buf_2
Xoutput122 net122 VGND VGND VPWR VPWR rdata[19] sky130_fd_sc_hd__buf_2
Xoutput144 net144 VGND VGND VPWR VPWR rresp[1] sky130_fd_sc_hd__buf_2
X_2557_ cordic_inst.cordic_inst.y\[2\] _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__and2_1
X_2488_ cordic_inst.cordic_inst.y\[22\] _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__nand2_1
X_4227_ cordic_inst.cordic_inst.cos_out\[24\] net223 _2188_ net317 VGND VGND VPWR
+ VPWR _2190_ sky130_fd_sc_hd__a31o_1
XFILLER_28_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ net260 _2128_ cordic_inst.cordic_inst.sin_out\[16\] VGND VGND VPWR VPWR _2129_
+ sky130_fd_sc_hd__a21o_1
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3109_ _1236_ _1401_ _1237_ _1234_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__a211o_1
XFILLER_43_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4089_ net226 _2068_ cordic_inst.cordic_inst.cos_out\[7\] VGND VGND VPWR VPWR _2069_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout382 net392 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_2
Xfanout393 net402 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_2
Xfanout360 net362 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_2
Xfanout371 net372 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput13 araddr[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xinput35 arvalid VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
Xinput24 araddr[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput46 awaddr[19] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput79 wdata[17] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
Xinput68 awvalid VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xinput57 awaddr[29] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
X_3460_ _1650_ _1654_ _1490_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__a21o_1
X_3391_ net242 _1578_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__nand2_1
X_2411_ net286 _0744_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2342_ net266 _0655_ _0658_ _0675_ net247 net240 VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux4_1
XFILLER_69_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4012_ net89 _2009_ _2012_ net352 VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o211a_1
X_2273_ axi_controller.state\[0\] VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__inv_2
XFILLER_80_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4914_ net387 _0013_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4845_ net404 _0084_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4776_ net407 _0503_ _0198_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[5\] sky130_fd_sc_hd__dfrtp_4
X_3727_ net254 _1844_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__nand2_1
X_3658_ cordic_inst.deg_handler_inst.theta_abs\[18\] _1787_ VGND VGND VPWR VPWR _1807_
+ sky130_fd_sc_hd__xnor2_1
X_2609_ _0677_ _0943_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__xor2_1
X_3589_ net183 net164 net315 VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux2_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout190 _1929_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_2
XFILLER_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2960_ cordic_inst.cordic_inst.x\[3\] _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__nand2_1
X_2891_ _1190_ _1192_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__or3_1
XFILLER_30_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4630_ net409 _0361_ net342 VGND VGND VPWR VPWR axi_controller.result_out\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4561_ net359 _0293_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[27\] sky130_fd_sc_hd__dfxtp_1
X_3512_ _1540_ _1729_ _1730_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__o21ba_1
X_4492_ net345 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__inv_2
X_3443_ cordic_inst.cordic_inst.angle\[28\] net170 net159 cordic_inst.cordic_inst.z\[28\]
+ _1678_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a221o_1
X_3374_ _1498_ _1510_ _1577_ _1612_ _0609_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__o32a_1
XFILLER_69_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2325_ cordic_inst.cordic_inst.x\[19\] cordic_inst.cordic_inst.x\[20\] cordic_inst.cordic_inst.x\[21\]
+ cordic_inst.cordic_inst.x\[22\] net306 net298 VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux4_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4828_ net367 _0555_ _0250_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[25\] sky130_fd_sc_hd__dfrtp_2
X_4759_ net394 _0486_ _0181_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_89_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3090_ cordic_inst.cordic_inst.x\[25\] _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__and2_1
XFILLER_66_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3992_ net93 net320 _1999_ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2943_ _1116_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__xor2_1
X_2874_ _1173_ _1176_ net279 VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux2_1
X_4613_ net377 _0345_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[31\] sky130_fd_sc_hd__dfxtp_1
X_4544_ net357 _0276_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[10\] sky130_fd_sc_hd__dfxtp_1
X_4475_ net333 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__inv_2
X_3426_ _1663_ _1664_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__nor2_1
X_3357_ cordic_inst.cordic_inst.z\[1\] _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__and2_1
X_2308_ net238 _0642_ _0637_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a21bo_1
X_3288_ _1525_ _1526_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__nand2_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ cordic_inst.cordic_inst.y\[14\] _0923_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__xnor2_1
X_4260_ cordic_inst.cordic_inst.cos_out\[28\] _2218_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3211_ cordic_inst.cordic_inst.y\[22\] cordic_inst.cordic_inst.sin_out\[22\] net208
+ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux2_1
X_4191_ _2154_ _2158_ axi_controller.result_out\[19\] net202 VGND VGND VPWR VPWR _0373_
+ sky130_fd_sc_hd__o2bb2a_1
X_3142_ _1357_ _1432_ _1355_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_78_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3073_ _1349_ _1375_ _1372_ _1370_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__o211a_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3975_ axi_controller.write_addr_reg\[24\] net52 net187 VGND VGND VPWR VPWR _0323_
+ sky130_fd_sc_hd__mux2_1
X_2926_ _1077_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__xnor2_1
X_2857_ net219 _1108_ _1158_ net286 VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__a22o_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2788_ net232 _1087_ _1071_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a21o_1
X_4527_ net388 _0259_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[9\] sky130_fd_sc_hd__dfxtp_1
X_4458_ net343 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__inv_2
X_3409_ _1646_ _1647_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ net326 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
XFILLER_85_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3760_ axi_controller.reg_input_data\[15\] axi_controller.reg_input_data\[14\] axi_controller.reg_input_data\[13\]
+ axi_controller.reg_input_data\[12\] VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__or4_1
X_2711_ _0858_ _1029_ _0854_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3691_ cordic_inst.deg_handler_inst.theta_norm\[5\] cordic_inst.deg_handler_inst.theta_norm\[4\]
+ _1819_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__or3_1
X_2642_ cordic_inst.cordic_inst.y\[24\] _0975_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__nor2_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2573_ _0906_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and2_1
X_4312_ net136 net191 net156 axi_controller.result_out\[31\] VGND VGND VPWR VPWR _0563_
+ sky130_fd_sc_hd__a22o_1
X_4243_ cordic_inst.deg_handler_inst.kuadran\[0\] _2203_ _0605_ VGND VGND VPWR VPWR
+ _2204_ sky130_fd_sc_hd__o21a_1
XFILLER_87_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4174_ cordic_inst.cordic_inst.sin_out\[17\] cordic_inst.cordic_inst.sin_out\[16\]
+ _2128_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__or3_1
XFILLER_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3125_ _1359_ _1362_ _1367_ _1332_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__or4b_1
X_3056_ _1355_ _1358_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__or2_1
XFILLER_82_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3958_ axi_controller.write_addr_reg\[7\] net65 net190 VGND VGND VPWR VPWR _0306_
+ sky130_fd_sc_hd__mux2_1
X_3889_ axi_controller.reg_input_data\[11\] _1964_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__or2_1
X_2909_ _1070_ _1181_ net278 VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ net373 _0031_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_4861_ net384 _0070_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[25\] sky130_fd_sc_hd__dfxtp_1
X_3812_ _1907_ _1908_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_15_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4792_ net395 _0519_ _0214_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[21\] sky130_fd_sc_hd__dfrtp_4
X_3743_ net253 _1854_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__nand2_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3674_ cordic_inst.deg_handler_inst.theta_abs\[25\] net149 VGND VGND VPWR VPWR _0070_
+ sky130_fd_sc_hd__and2_1
X_2625_ _0936_ _0948_ _0955_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__or4_1
Xoutput112 net112 VGND VGND VPWR VPWR rdata[0] sky130_fd_sc_hd__buf_2
Xoutput123 net123 VGND VGND VPWR VPWR rdata[1] sky130_fd_sc_hd__buf_2
Xoutput134 net134 VGND VGND VPWR VPWR rdata[2] sky130_fd_sc_hd__buf_2
Xoutput145 net145 VGND VGND VPWR VPWR rvalid sky130_fd_sc_hd__buf_2
X_2556_ _0738_ _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__xnor2_1
X_2487_ _0794_ _0799_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_34_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4226_ net223 _2188_ cordic_inst.cordic_inst.cos_out\[24\] VGND VGND VPWR VPWR _2189_
+ sky130_fd_sc_hd__a21oi_1
X_4157_ cordic_inst.cordic_inst.sin_out\[15\] _2123_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__or2_1
X_3108_ _1234_ _1237_ _1401_ _1236_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__o211ai_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4088_ cordic_inst.cordic_inst.cos_out\[6\] cordic_inst.cordic_inst.cos_out\[5\]
+ cordic_inst.cordic_inst.cos_out\[4\] _2048_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__or4_2
X_3039_ cordic_inst.cordic_inst.x\[20\] _1340_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__or2_1
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout350 net351 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_2
Xfanout361 net362 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_2
Xfanout383 net386 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_2
Xfanout372 net375 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_2
Xfanout394 net395 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_61_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput25 araddr[30] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 araddr[20] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput36 awaddr[0] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput69 bready VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_70_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput58 awaddr[2] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput47 awaddr[1] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
X_2410_ net220 _0700_ _0704_ net221 VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a22o_1
X_3390_ _1532_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__nand2_1
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2341_ net240 _0658_ _0637_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a21bo_1
XFILLER_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2272_ net302 VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__inv_2
X_4011_ axi_controller.reg_input_data\[26\] _2008_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__or2_1
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4913_ net389 _0012_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4844_ net413 _0083_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4775_ net408 _0502_ _0197_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[4\] sky130_fd_sc_hd__dfrtp_2
X_3726_ cordic_inst.deg_handler_inst.theta_norm\[18\] _1842_ VGND VGND VPWR VPWR _1844_
+ sky130_fd_sc_hd__or2_1
X_3657_ _1774_ _1787_ net148 net150 cordic_inst.deg_handler_inst.theta_abs\[17\] VGND
+ VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a32o_1
X_3588_ net302 net167 _1509_ net185 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a22o_1
X_2608_ net153 _0758_ _0764_ net250 VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__a31o_1
XFILLER_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2539_ cordic_inst.cordic_inst.y\[7\] _0872_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__nor2_1
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4209_ _0613_ _2173_ cordic_inst.cordic_inst.cos_out\[22\] VGND VGND VPWR VPWR _2174_
+ sky130_fd_sc_hd__a21o_1
XFILLER_73_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcordic_system_415 VGND VGND VPWR VPWR cordic_system_415/HI bresp[0] sky130_fd_sc_hd__conb_1
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout180 net181 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_2
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout191 net194 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2890_ net263 _1075_ _1114_ _1106_ net239 net243 VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__mux4_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ net359 _0292_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[26\] sky130_fd_sc_hd__dfxtp_1
X_3511_ _1540_ _1729_ net177 VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__a21o_1
X_4491_ net345 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__inv_2
X_3442_ _1477_ _1666_ _1677_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__a21oi_1
X_3373_ net287 net313 VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__or2_1
X_2324_ _0655_ _0658_ net283 VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux2_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4827_ net368 _0554_ _0249_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[24\] sky130_fd_sc_hd__dfrtp_2
X_4758_ net394 _0485_ _0180_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3709_ cordic_inst.deg_handler_inst.theta_norm\[12\] _1833_ VGND VGND VPWR VPWR _0011_
+ sky130_fd_sc_hd__xnor2_1
X_4689_ net396 _0416_ _0111_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3991_ net351 _2000_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2942_ _1131_ _1178_ net250 VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a21o_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2873_ net285 _1174_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__o21ai_1
X_4612_ net377 _0344_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[30\] sky130_fd_sc_hd__dfxtp_1
X_4543_ net356 _0275_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4474_ net333 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__inv_2
X_3425_ cordic_inst.cordic_inst.z\[27\] cordic_inst.cordic_inst.z\[26\] net249 VGND
+ VGND VPWR VPWR _1664_ sky130_fd_sc_hd__o21a_1
X_3356_ _1585_ _1587_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__xnor2_1
X_3287_ cordic_inst.cordic_inst.z\[15\] _1524_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__nand2_1
X_2307_ net233 _0641_ _0635_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__a21o_1
XFILLER_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4190_ _2156_ _2157_ net202 VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__o21a_1
X_3210_ cordic_inst.cordic_inst.y\[23\] cordic_inst.cordic_inst.sin_out\[23\] net208
+ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux2_1
XFILLER_79_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3141_ _1358_ _1431_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3072_ _1359_ _1365_ _1373_ _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__o31a_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3974_ axi_controller.write_addr_reg\[23\] net51 net187 VGND VGND VPWR VPWR _0322_
+ sky130_fd_sc_hd__mux2_1
X_2925_ net270 _1227_ _1226_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__a21oi_1
X_2856_ net216 _1142_ _1144_ _0713_ net282 VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a221o_1
X_2787_ net278 _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__nor2_1
X_4526_ net388 _0258_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[8\] sky130_fd_sc_hd__dfxtp_1
X_4457_ net343 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__inv_2
X_3408_ cordic_inst.cordic_inst.z\[17\] _1644_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__and2_1
X_4388_ net327 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
X_3339_ _1498_ _1577_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2710_ _1031_ _1032_ cordic_inst.cordic_inst.y\[19\] net160 VGND VGND VPWR VPWR _0549_
+ sky130_fd_sc_hd__a2bb2o_1
X_3690_ cordic_inst.deg_handler_inst.theta_norm\[5\] _1821_ VGND VGND VPWR VPWR _0035_
+ sky130_fd_sc_hd__xnor2_1
X_2641_ cordic_inst.cordic_inst.y\[24\] _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2572_ cordic_inst.cordic_inst.y\[4\] _0886_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__xor2_1
X_4311_ net191 _1976_ _1987_ _2252_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__and4b_4
X_4242_ cordic_inst.cordic_inst.cos_out\[25\] _2196_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__nor2_1
X_4173_ _2139_ _2142_ axi_controller.result_out\[17\] net201 VGND VGND VPWR VPWR _0371_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_2_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3124_ net178 _1382_ _1419_ net158 cordic_inst.cordic_inst.x\[24\] VGND VGND VPWR
+ VPWR _0522_ sky130_fd_sc_hd__a32o_1
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3055_ cordic_inst.cordic_inst.x\[18\] _1356_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_18_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3957_ axi_controller.write_addr_reg\[6\] net64 net190 VGND VGND VPWR VPWR _0305_
+ sky130_fd_sc_hd__mux2_1
X_2908_ net243 _1183_ net215 VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__a21o_1
X_3888_ net72 _1965_ _1968_ net354 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__o211a_1
X_2839_ cordic_inst.cordic_inst.y\[4\] cordic_inst.cordic_inst.y\[5\] net314 VGND
+ VGND VPWR VPWR _1142_ sky130_fd_sc_hd__mux2_1
X_4509_ net324 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__inv_2
XFILLER_86_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4860_ net384 _0069_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3811_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1903_
+ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_15_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4791_ net395 _0518_ _0213_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[20\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3742_ cordic_inst.deg_handler_inst.theta_norm\[24\] _1852_ VGND VGND VPWR VPWR _1854_
+ sky130_fd_sc_hd__or2_1
X_3673_ cordic_inst.deg_handler_inst.theta_abs\[24\] net149 VGND VGND VPWR VPWR _0069_
+ sky130_fd_sc_hd__and2_1
X_2624_ _0957_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nand2_1
Xoutput124 net124 VGND VGND VPWR VPWR rdata[20] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR rdata[10] sky130_fd_sc_hd__buf_2
Xoutput135 net135 VGND VGND VPWR VPWR rdata[30] sky130_fd_sc_hd__buf_2
Xoutput146 net146 VGND VGND VPWR VPWR wready sky130_fd_sc_hd__buf_2
X_2555_ _0718_ _0735_ net276 VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__o21ai_1
X_2486_ _0817_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__or2_1
XFILLER_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4225_ cordic_inst.cordic_inst.cos_out\[23\] cordic_inst.cordic_inst.cos_out\[22\]
+ _2173_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__or3_1
X_4156_ axi_controller.result_out\[15\] net201 _2127_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__o21ba_1
X_3107_ cordic_inst.cordic_inst.x\[30\] net159 _1408_ net179 VGND VGND VPWR VPWR _0528_
+ sky130_fd_sc_hd__a22o_1
X_4087_ net262 _2065_ cordic_inst.cordic_inst.sin_out\[7\] VGND VGND VPWR VPWR _2067_
+ sky130_fd_sc_hd__a21oi_1
X_3038_ cordic_inst.cordic_inst.x\[20\] _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__nand2_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout340 net341 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__buf_2
Xfanout351 net34 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_2
Xfanout362 net364 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout384 net386 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_2
Xfanout373 net375 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout395 net402 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput26 araddr[31] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 araddr[21] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput37 awaddr[10] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 awaddr[20] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput59 awaddr[30] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2340_ _0673_ _0674_ net292 VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__mux2_1
X_2271_ net294 VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__inv_2
XFILLER_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4010_ net88 _2009_ _2011_ net352 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__o211a_1
XFILLER_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4912_ net389 _0011_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4843_ net403 _0082_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[7\] sky130_fd_sc_hd__dfxtp_1
X_4774_ net408 _0501_ _0196_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[3\] sky130_fd_sc_hd__dfrtp_2
X_3725_ cordic_inst.deg_handler_inst.theta_norm\[18\] _1843_ VGND VGND VPWR VPWR _0017_
+ sky130_fd_sc_hd__xnor2_1
X_3656_ _1773_ net148 _1806_ net150 cordic_inst.deg_handler_inst.theta_abs\[16\] VGND
+ VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a32o_1
X_2607_ _0940_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__nor2_1
X_3587_ net182 _1576_ _1581_ net163 net294 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a32o_1
XFILLER_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2538_ cordic_inst.cordic_inst.y\[7\] _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__and2_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4208_ cordic_inst.cordic_inst.cos_out\[21\] _2166_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__or2_1
X_2469_ net268 _0797_ _0803_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a21o_1
XFILLER_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4139_ cordic_inst.cordic_inst.cos_out\[13\] net224 _2111_ net318 VGND VGND VPWR
+ VPWR _2113_ sky130_fd_sc_hd__a31o_1
XFILLER_71_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcordic_system_416 VGND VGND VPWR VPWR cordic_system_416/HI rresp[0] sky130_fd_sc_hd__conb_1
Xfanout192 net194 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_4
Xfanout181 net186 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xfanout170 net171 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3510_ _1545_ _1623_ _1544_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__a21oi_1
X_4490_ net345 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
X_3441_ net174 _1667_ VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__or2_1
X_3372_ _1554_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__or2_1
X_2323_ net265 _0632_ _0640_ _0656_ net231 net233 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_68_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4826_ net368 _0553_ _0248_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[23\] sky130_fd_sc_hd__dfrtp_4
X_4757_ net396 _0484_ _0179_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3708_ net255 _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__nand2_1
X_4688_ net399 _0415_ _0110_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_3639_ cordic_inst.deg_handler_inst.theta_abs\[8\] _1764_ VGND VGND VPWR VPWR _1798_
+ sky130_fd_sc_hd__nand2_1
XFILLER_88_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3990_ net71 net338 _1999_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2941_ cordic_inst.cordic_inst.x\[7\] _1242_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__nand2_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4611_ net377 _0343_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[29\] sky130_fd_sc_hd__dfxtp_1
X_2872_ net235 _1079_ _1071_ net241 VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__a211o_1
X_4542_ net356 _0274_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[8\] sky130_fd_sc_hd__dfxtp_1
X_4473_ net330 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__inv_2
X_3424_ cordic_inst.cordic_inst.z\[25\] cordic_inst.cordic_inst.z\[24\] net249 VGND
+ VGND VPWR VPWR _1663_ sky130_fd_sc_hd__o21a_1
X_3355_ cordic_inst.cordic_inst.z\[2\] _1593_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__nand2_1
X_3286_ cordic_inst.cordic_inst.z\[15\] _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__or2_1
X_2306_ cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.x\[29\] cordic_inst.cordic_inst.x\[30\]
+ net265 net307 net297 VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux4_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4809_ net406 _0536_ _0231_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ _1373_ _1430_ _1365_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__a21o_1
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3071_ _1354_ _1357_ _1353_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__a21o_1
XFILLER_54_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3973_ axi_controller.write_addr_reg\[22\] net50 net187 VGND VGND VPWR VPWR _0321_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2924_ net280 _1191_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__nor2_1
X_2855_ _1104_ _1107_ net235 VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__mux2_1
X_2786_ net239 _1088_ _1070_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__a21boi_1
X_4525_ net371 _0004_ VGND VGND VPWR VPWR axi_controller.state\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4456_ net343 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4387_ net327 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
X_3407_ _1645_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__inv_2
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3338_ _0711_ _1576_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3269_ net222 _0707_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__nand2_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2640_ _0795_ _0801_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2571_ _0902_ _0904_ _0889_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__a21o_1
X_4310_ net82 net103 _1930_ _1994_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__and4_1
X_4241_ axi_controller.result_out\[25\] _2202_ net199 VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux2_1
X_4172_ net319 _2141_ net201 VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3123_ _1377_ _1381_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__or2_1
X_3054_ cordic_inst.cordic_inst.x\[18\] _1356_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__nand2_1
XFILLER_82_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3956_ axi_controller.write_addr_reg\[5\] net63 net189 VGND VGND VPWR VPWR _0304_
+ sky130_fd_sc_hd__mux2_1
X_2907_ net243 _1115_ net215 VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a21o_1
XFILLER_31_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3887_ axi_controller.reg_input_data\[10\] _1964_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__or2_1
X_2838_ _1139_ _1140_ net292 VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__mux2_1
X_2769_ net264 net296 VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__and2_1
X_4508_ net324 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__inv_2
X_4439_ net332 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__inv_2
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3810_ axi_controller.reg_input_data\[27\] _1905_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_15_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4790_ net394 _0517_ _0212_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3741_ cordic_inst.deg_handler_inst.theta_norm\[24\] _1853_ VGND VGND VPWR VPWR _0024_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3672_ cordic_inst.deg_handler_inst.theta_abs\[23\] cordic_inst.deg_handler_inst.theta_abs\[31\]
+ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__and2_1
X_2623_ _0598_ _0956_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__nand2_1
Xoutput125 net125 VGND VGND VPWR VPWR rdata[21] sky130_fd_sc_hd__buf_2
Xoutput114 net114 VGND VGND VPWR VPWR rdata[11] sky130_fd_sc_hd__buf_2
X_2554_ cordic_inst.cordic_inst.y\[3\] _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__and2_1
Xoutput136 net136 VGND VGND VPWR VPWR rdata[31] sky130_fd_sc_hd__buf_2
X_2485_ _0595_ _0816_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__and2_1
X_4224_ axi_controller.result_out\[24\] net200 VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__nor2_1
X_4155_ _2121_ _2122_ _2126_ net201 VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__o211a_1
X_3106_ _1231_ _1402_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__xor2_1
XFILLER_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4086_ cordic_inst.cordic_inst.sin_out\[7\] net262 _2065_ VGND VGND VPWR VPWR _2066_
+ sky130_fd_sc_hd__and3_1
XFILLER_70_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3037_ _1208_ _1218_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__xor2_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3939_ axi_controller.read_addr_reg\[29\] axi_controller.read_addr_reg\[30\] VGND
+ VGND VPWR VPWR _1982_ sky130_fd_sc_hd__nand2_1
XFILLER_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout330 net333 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__buf_2
Xfanout341 net348 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__buf_4
Xfanout352 net353 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_2
Xfanout363 net364 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
Xfanout374 net375 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout396 net398 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_2
Xfanout385 net386 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_2
XFILLER_46_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 araddr[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 araddr[22] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput49 awaddr[21] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 awaddr[11] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2270_ net289 VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__inv_2
XFILLER_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4911_ net390 _0010_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4842_ net403 _0081_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[6\] sky130_fd_sc_hd__dfxtp_1
X_4773_ net408 _0500_ _0195_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[2\] sky130_fd_sc_hd__dfrtp_2
X_3724_ net254 _1842_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__nand2_1
X_3655_ cordic_inst.deg_handler_inst.theta_abs\[16\] _1772_ VGND VGND VPWR VPWR _1806_
+ sky130_fd_sc_hd__nand2_1
X_2606_ _0938_ cordic_inst.cordic_inst.y\[11\] VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__and2b_1
X_3586_ _1756_ _1757_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and2_1
X_2537_ _0684_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__xor2_1
X_2468_ net269 _0796_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21o_1
X_4207_ axi_controller.result_out\[21\] _2172_ net202 VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
X_2399_ net288 _0728_ _0732_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__a211o_1
X_4138_ net224 _2111_ cordic_inst.cordic_inst.cos_out\[13\] VGND VGND VPWR VPWR _2112_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_54_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4069_ net204 _2051_ _2044_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_26_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout160 net161 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
XFILLER_19_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout171 _0628_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xfanout182 net183 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_2
XFILLER_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout193 net194 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
XFILLER_74_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3440_ net179 _1675_ _1676_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a21o_1
X_3371_ _1561_ _1608_ _1556_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__o21ba_1
X_2322_ _0640_ _0656_ net231 VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__mux2_1
XFILLER_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4825_ net393 _0552_ _0247_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[22\] sky130_fd_sc_hd__dfrtp_2
X_4756_ net396 _0483_ _0178_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3707_ cordic_inst.deg_handler_inst.theta_norm\[11\] cordic_inst.deg_handler_inst.theta_norm\[10\]
+ _1829_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__or3_1
X_4687_ net399 _0414_ _0109_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3638_ _1764_ net147 _1797_ net151 cordic_inst.deg_handler_inst.theta_abs\[7\] VGND
+ VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a32o_1
X_3569_ cordic_inst.cordic_inst.x\[10\] cordic_inst.cordic_inst.cos_out\[10\] net210
+ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_68_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2940_ cordic_inst.cordic_inst.x\[7\] _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__nor2_1
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2871_ _1133_ _1135_ net291 VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__mux2_1
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4610_ net377 _0342_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4541_ net360 _0273_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_4472_ net331 VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__inv_2
X_3423_ _1660_ _1661_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__nand2_1
X_3354_ _1582_ _1588_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__xor2_1
X_3285_ net277 _1481_ _1523_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__mux2_1
X_2305_ cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.x\[29\] net307 VGND
+ VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux2_1
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4808_ net407 _0535_ _0230_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[5\] sky130_fd_sc_hd__dfrtp_2
X_4739_ net405 _0466_ _0161_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3070_ cordic_inst.cordic_inst.x\[16\] _1360_ _1364_ cordic_inst.cordic_inst.x\[17\]
+ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__a22oi_1
XFILLER_47_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3972_ axi_controller.write_addr_reg\[21\] net49 net187 VGND VGND VPWR VPWR _0320_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2923_ _1082_ _1225_ net270 VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__o21a_1
X_2854_ _1153_ _1155_ _1156_ _1151_ net247 VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__o32a_1
X_2785_ _1084_ _1087_ net292 VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4524_ net371 _0003_ VGND VGND VPWR VPWR axi_controller.state\[2\] sky130_fd_sc_hd__dfxtp_1
X_4455_ net345 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__inv_2
X_4386_ net327 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
X_3406_ cordic_inst.cordic_inst.z\[17\] _1644_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__or2_1
X_3337_ net304 net313 net294 VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_5_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3268_ net251 _0705_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__or2_1
XFILLER_73_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3199_ _0603_ net171 VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__nor2_1
XFILLER_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2570_ _0902_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4240_ net316 _2197_ _2198_ _2200_ _2201_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__o32ai_1
X_4171_ cordic_inst.cordic_inst.cos_out\[17\] _2140_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__xnor2_1
X_3122_ cordic_inst.cordic_inst.x\[25\] net158 _1418_ net178 VGND VGND VPWR VPWR _0523_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3053_ _1204_ _1350_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__xor2_1
XFILLER_67_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3955_ axi_controller.write_addr_reg\[4\] net62 net189 VGND VGND VPWR VPWR _0303_
+ sky130_fd_sc_hd__mux2_1
X_2906_ _1206_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__nand2_1
X_3886_ net102 _1965_ _1967_ net354 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o211a_1
X_2837_ cordic_inst.cordic_inst.y\[12\] cordic_inst.cordic_inst.y\[13\] cordic_inst.cordic_inst.y\[14\]
+ cordic_inst.cordic_inst.y\[15\] net309 net299 VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__mux4_1
X_2768_ net263 net291 VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and2_1
X_4507_ net329 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__inv_2
X_2699_ cordic_inst.cordic_inst.y\[23\] net159 _1025_ net178 VGND VGND VPWR VPWR _0553_
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4438_ net332 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
X_4369_ net334 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
XFILLER_73_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3740_ net253 _1852_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__nand2_1
X_3671_ net148 _1814_ _1815_ net149 cordic_inst.deg_handler_inst.theta_abs\[22\] VGND
+ VGND VPWR VPWR _0067_ sky130_fd_sc_hd__a32o_1
X_2622_ _0598_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__or2_1
Xoutput115 net115 VGND VGND VPWR VPWR rdata[12] sky130_fd_sc_hd__buf_2
X_2553_ _0742_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__xnor2_1
Xoutput137 net137 VGND VGND VPWR VPWR rdata[3] sky130_fd_sc_hd__buf_2
Xoutput126 net126 VGND VGND VPWR VPWR rdata[22] sky130_fd_sc_hd__buf_2
X_2484_ cordic_inst.cordic_inst.y\[29\] _0814_ _0817_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4223_ _2183_ _2186_ axi_controller.result_out\[23\] net200 VGND VGND VPWR VPWR _0377_
+ sky130_fd_sc_hd__o2bb2a_1
X_4154_ _2124_ _2125_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__or2_1
X_3105_ net179 _1406_ _1407_ net159 net266 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a32o_1
X_4085_ cordic_inst.cordic_inst.sin_out\[6\] cordic_inst.cordic_inst.sin_out\[5\]
+ cordic_inst.cordic_inst.sin_out\[4\] _2045_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__or4_1
X_3036_ _1337_ _1338_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__nand2_1
XFILLER_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3938_ axi_controller.read_addr_reg\[17\] _1980_ axi_controller.read_addr_reg\[2\]
+ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__or3b_1
X_3869_ axi_controller.write_addr_reg\[12\] axi_controller.write_addr_reg\[15\] axi_controller.write_addr_reg\[14\]
+ axi_controller.write_addr_reg\[17\] VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__or4_1
XFILLER_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout331 net332 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__buf_4
Xfanout320 axi_controller.mode VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_4
Xfanout353 net355 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout364 net414 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_2
Xfanout342 net344 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_4
Xfanout375 net392 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout397 net398 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__buf_1
Xfanout386 net392 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 araddr[23] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 araddr[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 awaddr[12] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_20_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4910_ net390 _0009_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4841_ net403 _0080_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4772_ net408 _0499_ _0194_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[1\] sky130_fd_sc_hd__dfrtp_2
X_3723_ cordic_inst.deg_handler_inst.theta_norm\[17\] cordic_inst.deg_handler_inst.theta_norm\[16\]
+ _1839_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__or3_1
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3654_ _1772_ net148 _1805_ net152 cordic_inst.deg_handler_inst.theta_abs\[15\] VGND
+ VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a32o_1
X_2605_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__inv_2
X_3585_ net157 _1580_ net289 VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__a21o_1
X_2536_ _0693_ net153 _0757_ net250 VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__a31o_1
X_2467_ net269 _0795_ _0801_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__a21bo_1
X_4206_ net318 _2170_ _2171_ _2167_ _2168_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__a32o_1
XFILLER_68_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2398_ cordic_inst.cordic_inst.x\[1\] net222 _0711_ _0730_ net220 VGND VGND VPWR
+ VPWR _0733_ sky130_fd_sc_hd__a32o_1
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4137_ cordic_inst.cordic_inst.cos_out\[12\] cordic_inst.cordic_inst.cos_out\[11\]
+ cordic_inst.cordic_inst.cos_out\[10\] _2089_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__or4_2
XFILLER_56_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4068_ net230 _2046_ _2047_ _2049_ _2050_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__o32a_1
X_3019_ cordic_inst.cordic_inst.x\[10\] _1320_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_2
Xfanout161 net162 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net186 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_2
Xfanout150 _1781_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout194 _1927_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_8
XFILLER_74_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3370_ _1561_ _1608_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__nor2_1
XFILLER_69_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2321_ cordic_inst.cordic_inst.x\[26\] cordic_inst.cordic_inst.x\[27\] net307 VGND
+ VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4824_ net393 _0551_ _0246_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[21\] sky130_fd_sc_hd__dfrtp_2
X_4755_ net396 _0482_ _0177_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3706_ cordic_inst.deg_handler_inst.theta_norm\[11\] _1831_ VGND VGND VPWR VPWR _0010_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4686_ net399 _0413_ _0108_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3637_ cordic_inst.deg_handler_inst.theta_abs\[7\] _1763_ VGND VGND VPWR VPWR _1797_
+ sky130_fd_sc_hd__nand2_1
X_3568_ cordic_inst.cordic_inst.x\[11\] cordic_inst.cordic_inst.cos_out\[11\] net210
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
X_2519_ _0852_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__nand2_1
XFILLER_88_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3499_ cordic_inst.cordic_inst.angle\[15\] net173 net168 cordic_inst.cordic_inst.z\[15\]
+ _1721_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__a221o_1
XFILLER_75_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2870_ net285 _1171_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4540_ net360 _0272_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4471_ net331 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__inv_2
X_3422_ net273 cordic_inst.cordic_inst.z\[26\] VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__xnor2_1
X_3353_ cordic_inst.cordic_inst.z\[3\] _1590_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3284_ _0707_ _1521_ net289 VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__a21o_1
X_2304_ net243 _0638_ net169 VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a21o_1
XFILLER_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4807_ net406 _0534_ _0229_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2999_ cordic_inst.cordic_inst.x\[14\] _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__nand2_1
X_4738_ net385 _0465_ _0160_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[31\] sky130_fd_sc_hd__dfrtp_2
X_4669_ net376 _0398_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[23\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_8_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3971_ axi_controller.write_addr_reg\[20\] net48 net187 VGND VGND VPWR VPWR _0319_
+ sky130_fd_sc_hd__mux2_1
X_2922_ net268 _1214_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2853_ cordic_inst.cordic_inst.y\[1\] net222 _0711_ _1121_ net220 VGND VGND VPWR
+ VPWR _1156_ sky130_fd_sc_hd__a32o_1
X_2784_ cordic_inst.cordic_inst.y\[27\] cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.y\[29\]
+ cordic_inst.cordic_inst.y\[30\] net305 net296 VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_41_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4523_ net371 _0002_ VGND VGND VPWR VPWR axi_controller.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_4454_ net345 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__inv_2
X_4385_ net326 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
X_3405_ net251 _1643_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__xnor2_1
X_3336_ cordic_inst.cordic_inst.z\[4\] _1574_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__nand2_1
XFILLER_58_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3267_ cordic_inst.cordic_inst.z\[13\] _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__and2_1
X_3198_ net184 _1148_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__nand2_1
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4170_ cordic_inst.cordic_inst.cos_out\[16\] _2132_ net224 VGND VGND VPWR VPWR _2140_
+ sky130_fd_sc_hd__o21a_1
X_3121_ _1395_ _1417_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__xnor2_1
X_3052_ _1353_ _1354_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__nand2b_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3954_ axi_controller.write_addr_reg\[3\] net61 net189 VGND VGND VPWR VPWR _0302_
+ sky130_fd_sc_hd__mux2_1
X_3885_ axi_controller.reg_input_data\[9\] _1964_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__or2_1
X_2905_ net279 _1176_ _1069_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__o21a_1
XFILLER_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2836_ cordic_inst.cordic_inst.y\[8\] cordic_inst.cordic_inst.y\[9\] cordic_inst.cordic_inst.y\[10\]
+ cordic_inst.cordic_inst.y\[11\] net310 net299 VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__mux4_1
X_2767_ net263 net283 VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__nand2_2
X_2698_ _0830_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__xnor2_1
X_4506_ net324 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__inv_2
X_4437_ net332 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__inv_2
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4368_ net335 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
X_3319_ net237 net314 VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__and2_1
X_4299_ axi_controller.reg_input_data\[21\] _2242_ VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__or2_1
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3670_ _1783_ _1808_ _0617_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__o21ai_1
X_2621_ _0760_ _0949_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__xnor2_1
Xoutput116 net116 VGND VGND VPWR VPWR rdata[13] sky130_fd_sc_hd__buf_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2552_ _0718_ _0735_ _0738_ net276 VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__o31a_1
Xoutput127 net127 VGND VGND VPWR VPWR rdata[23] sky130_fd_sc_hd__buf_2
Xoutput138 net138 VGND VGND VPWR VPWR rdata[4] sky130_fd_sc_hd__buf_2
X_4222_ net317 _2185_ net200 VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__o21a_1
X_2483_ cordic_inst.cordic_inst.y\[29\] _0814_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_91_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4153_ cordic_inst.cordic_inst.sin_out\[15\] net260 _2123_ net228 VGND VGND VPWR
+ VPWR _2125_ sky130_fd_sc_hd__a31o_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3104_ _1230_ _1403_ _1405_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__or3_1
X_4084_ axi_controller.result_out\[7\] net203 VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__nor2_1
X_3035_ cordic_inst.cordic_inst.x\[22\] _1336_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__or2_1
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3937_ axi_controller.read_addr_reg\[16\] axi_controller.read_addr_reg\[19\] axi_controller.read_addr_reg\[18\]
+ axi_controller.read_addr_reg\[21\] VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__or4_1
X_3868_ axi_controller.write_addr_reg\[8\] axi_controller.write_addr_reg\[11\] axi_controller.write_addr_reg\[10\]
+ axi_controller.write_addr_reg\[13\] VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__or4_1
X_3799_ axi_controller.reg_input_data\[23\] _1892_ axi_controller.reg_input_data\[24\]
+ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__a21oi_1
X_2819_ cordic_inst.cordic_inst.y\[9\] cordic_inst.cordic_inst.y\[10\] cordic_inst.cordic_inst.y\[11\]
+ cordic_inst.cordic_inst.y\[12\] net310 net300 VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux4_1
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout321 net328 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_4
Xfanout332 net333 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_4
Xfanout310 net311 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_2
Xfanout354 net355 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_2
Xfanout365 net366 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_2
Xfanout343 net344 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__buf_4
Xfanout376 net382 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout387 net389 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout398 net402 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__buf_2
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 araddr[24] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 araddr[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4840_ net403 _0079_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4771_ net406 _0498_ _0193_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[0\] sky130_fd_sc_hd__dfrtp_1
X_3722_ cordic_inst.deg_handler_inst.theta_norm\[17\] _1841_ VGND VGND VPWR VPWR _0016_
+ sky130_fd_sc_hd__xnor2_1
X_3653_ cordic_inst.deg_handler_inst.theta_abs\[15\] _1771_ VGND VGND VPWR VPWR _1805_
+ sky130_fd_sc_hd__nand2_1
X_2604_ cordic_inst.cordic_inst.y\[11\] _0938_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nand2b_1
X_3584_ _1755_ _1756_ net282 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
X_2535_ _0743_ _0757_ net250 VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21oi_1
X_2466_ net269 _0652_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a21oi_1
X_4205_ cordic_inst.cordic_inst.sin_out\[21\] net259 _2169_ VGND VGND VPWR VPWR _2171_
+ sky130_fd_sc_hd__nand3_1
X_4136_ _2108_ _2109_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__or2_1
XFILLER_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2397_ cordic_inst.cordic_inst.x\[2\] net217 _0709_ _0731_ net281 VGND VGND VPWR
+ VPWR _0732_ sky130_fd_sc_hd__a221o_1
XFILLER_68_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4067_ cordic_inst.cordic_inst.cos_out\[4\] net226 _2048_ net320 VGND VGND VPWR VPWR
+ _2050_ sky130_fd_sc_hd__a31o_1
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3018_ cordic_inst.cordic_inst.x\[10\] _1320_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_54_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
Xfanout173 _0628_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_2
Xfanout162 _0629_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout195 net196 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2320_ _0653_ _0654_ net295 VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_38_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4823_ net393 _0550_ _0245_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4754_ net398 _0481_ _0176_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3705_ cordic_inst.deg_handler_inst.theta_norm\[10\] _1829_ net255 VGND VGND VPWR
+ VPWR _1831_ sky130_fd_sc_hd__o21ai_1
X_4685_ net400 _0412_ _0107_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3636_ _1763_ net147 _1796_ net151 cordic_inst.deg_handler_inst.theta_abs\[6\] VGND
+ VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a32o_1
X_3567_ cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.cos_out\[12\] net210
+ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_2518_ _0596_ _0851_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__nand2_1
X_3498_ _1527_ _1719_ _1720_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2449_ _0631_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nand2_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4119_ cordic_inst.cordic_inst.sin_out\[11\] net261 _2093_ net229 VGND VGND VPWR
+ VPWR _2095_ sky130_fd_sc_hd__a31o_1
XFILLER_83_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4470_ net331 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__inv_2
X_3421_ net273 cordic_inst.cordic_inst.z\[27\] VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__xnor2_1
X_3352_ cordic_inst.cordic_inst.z\[3\] _1590_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__and2_1
X_2303_ net283 _0636_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__o21ai_1
XFILLER_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3283_ _1521_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4806_ net405 _0533_ _0228_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2998_ _1193_ _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4737_ net383 _0464_ _0159_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[30\] sky130_fd_sc_hd__dfrtp_1
X_4668_ net376 _0397_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[22\] sky130_fd_sc_hd__dfxtp_1
X_3619_ net152 _1786_ cordic_inst.deg_handler_inst.theta_abs\[0\] VGND VGND VPWR VPWR
+ _0053_ sky130_fd_sc_hd__o21a_1
X_4599_ net375 _0331_ VGND VGND VPWR VPWR axi_controller.rst sky130_fd_sc_hd__dfxtp_1
XFILLER_76_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3970_ axi_controller.write_addr_reg\[19\] net46 net187 VGND VGND VPWR VPWR _0318_
+ sky130_fd_sc_hd__mux2_1
X_2921_ net268 _1213_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2852_ cordic_inst.cordic_inst.y\[2\] net217 net216 _1154_ net282 VGND VGND VPWR
+ VPWR _1155_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2783_ cordic_inst.cordic_inst.y\[29\] cordic_inst.cordic_inst.y\[30\] net305 VGND
+ VGND VPWR VPWR _1086_ sky130_fd_sc_hd__mux2_1
X_4522_ net371 _0001_ VGND VGND VPWR VPWR axi_controller.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_4453_ net326 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__inv_2
X_3404_ net293 net313 _1498_ _1502_ net287 VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__a2111o_1
X_4384_ net326 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
X_3335_ _1481_ net274 _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__mux2_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3266_ net274 _1503_ _1504_ _1501_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3197_ net184 _1272_ _1469_ net166 cordic_inst.cordic_inst.x\[1\] VGND VGND VPWR
+ VPWR _0499_ sky130_fd_sc_hd__a32o_1
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3120_ _1377_ _1381_ _1379_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__a21oi_1
X_3051_ cordic_inst.cordic_inst.x\[19\] _1352_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__nand2_1
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3953_ axi_controller.write_addr_reg\[2\] net58 net190 VGND VGND VPWR VPWR _0301_
+ sky130_fd_sc_hd__mux2_1
X_3884_ net101 _1965_ _1966_ net354 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__o211a_1
X_2904_ _1069_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__nand2_1
X_2835_ net248 _1137_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__or2_1
X_2766_ net263 net279 VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nand2_1
X_2697_ _0825_ _1023_ _0823_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__a21bo_1
X_4505_ net329 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__inv_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4436_ net336 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__inv_2
X_4367_ net342 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
XFILLER_86_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3318_ net288 net237 _0712_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4298_ net83 _2243_ _2248_ net351 VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o211a_1
XFILLER_58_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3249_ cordic_inst.cordic_inst.z\[20\] _1487_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__nand2_1
XFILLER_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2620_ _0952_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nand2_1
X_2551_ _0750_ _0880_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__xnor2_2
Xoutput128 net128 VGND VGND VPWR VPWR rdata[24] sky130_fd_sc_hd__buf_2
X_2482_ _0595_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__nor2_1
Xoutput117 net117 VGND VGND VPWR VPWR rdata[14] sky130_fd_sc_hd__buf_2
Xoutput139 net139 VGND VGND VPWR VPWR rdata[5] sky130_fd_sc_hd__buf_2
X_4221_ cordic_inst.cordic_inst.cos_out\[23\] _2184_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_91_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4152_ net260 _2123_ cordic_inst.cordic_inst.sin_out\[15\] VGND VGND VPWR VPWR _2124_
+ sky130_fd_sc_hd__a21oi_1
X_3103_ _1230_ _1403_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__o21ai_1
X_4083_ axi_controller.result_out\[6\] _2063_ net203 VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux2_1
X_3034_ cordic_inst.cordic_inst.x\[22\] _1336_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__nand2_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3936_ _1976_ _1978_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__nand2_1
X_3867_ axi_controller.write_addr_reg\[1\] axi_controller.write_addr_reg\[0\] _1949_
+ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__or3_1
X_3798_ _1896_ _1897_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__xnor2_1
X_2818_ cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.y\[6\] cordic_inst.cordic_inst.y\[7\]
+ cordic_inst.cordic_inst.y\[8\] net312 net302 VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__mux4_1
X_2749_ net184 _1058_ _1059_ net166 cordic_inst.cordic_inst.y\[7\] VGND VGND VPWR
+ VPWR _0537_ sky130_fd_sc_hd__a32o_1
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout322 net328 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__buf_2
X_4419_ net337 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__inv_2
Xfanout311 cordic_inst.cordic_inst.i\[0\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_2
Xfanout300 net301 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_2
Xfanout355 net34 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_2
Xfanout333 net349 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_2
Xfanout366 net369 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_2
Xfanout344 net348 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_4
Xfanout388 net389 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_2
Xfanout377 net382 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_2
Xfanout399 net401 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 araddr[25] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4770_ net363 _0497_ _0192_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_3721_ cordic_inst.deg_handler_inst.theta_norm\[16\] _1839_ net256 VGND VGND VPWR
+ VPWR _1841_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3652_ _1771_ net148 _1804_ net152 cordic_inst.deg_handler_inst.theta_abs\[14\] VGND
+ VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a32o_1
X_2603_ _0769_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__xnor2_1
X_3583_ net171 _1755_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__nor2_1
X_2534_ _0850_ _0854_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__or3b_1
X_2465_ _0789_ _0791_ _0793_ _0794_ net269 VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__o41a_1
X_4204_ net259 _2169_ cordic_inst.cordic_inst.sin_out\[21\] VGND VGND VPWR VPWR _2170_
+ sky130_fd_sc_hd__a21o_1
X_2396_ cordic_inst.cordic_inst.x\[3\] cordic_inst.cordic_inst.x\[4\] net312 VGND
+ VGND VPWR VPWR _0731_ sky130_fd_sc_hd__mux2_1
X_4135_ cordic_inst.cordic_inst.sin_out\[13\] net260 _2107_ net228 VGND VGND VPWR
+ VPWR _2109_ sky130_fd_sc_hd__a31o_1
XFILLER_68_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4066_ net226 _2048_ cordic_inst.cordic_inst.cos_out\[4\] VGND VGND VPWR VPWR _2049_
+ sky130_fd_sc_hd__a21oi_1
X_3017_ _1187_ _1319_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__xor2_1
XFILLER_51_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4968_ net108 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4899_ net379 _0052_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_3919_ axi_controller.read_addr_reg\[20\] net14 net197 VGND VGND VPWR VPWR _0286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout152 _1781_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
Xfanout163 net165 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_4
Xfanout174 _0627_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_4
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout196 net197 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_2
XFILLER_47_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout185 net186 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4822_ net394 _0549_ _0244_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_33_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4753_ net399 _0480_ _0175_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3704_ cordic_inst.deg_handler_inst.theta_norm\[10\] _1830_ VGND VGND VPWR VPWR _0009_
+ sky130_fd_sc_hd__xnor2_1
X_4684_ net409 _0411_ _0106_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3635_ cordic_inst.deg_handler_inst.theta_abs\[6\] _1762_ VGND VGND VPWR VPWR _1796_
+ sky130_fd_sc_hd__nand2_1
X_3566_ cordic_inst.cordic_inst.x\[13\] cordic_inst.cordic_inst.cos_out\[13\] net210
+ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_88_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3497_ _1527_ _1719_ net183 VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__o21ai_1
X_2517_ _0596_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__or2_1
X_2448_ net244 _0725_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__nand2_1
X_2379_ net222 _0711_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__nand2_1
X_4118_ net261 _2093_ cordic_inst.cordic_inst.sin_out\[11\] VGND VGND VPWR VPWR _2094_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_67_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4049_ cordic_inst.cordic_inst.sin_out\[1\] cordic_inst.cordic_inst.sin_out\[0\]
+ net262 VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_39_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3420_ net273 cordic_inst.cordic_inst.z\[25\] VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__xor2_2
X_3351_ _1579_ _1589_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__xor2_1
X_2302_ net265 net284 VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nand2_2
X_3282_ net237 net313 VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__or2_1
XFILLER_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4805_ net406 _0532_ _0227_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2997_ _1189_ _1190_ _1192_ net271 VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__o31a_1
X_4736_ net383 _0463_ _0158_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[29\] sky130_fd_sc_hd__dfrtp_1
X_4667_ net376 _0396_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[21\] sky130_fd_sc_hd__dfxtp_2
X_3618_ _1785_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__inv_2
X_4598_ net362 _0330_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[31\] sky130_fd_sc_hd__dfxtp_1
X_3549_ cordic_inst.cordic_inst.x\[30\] cordic_inst.cordic_inst.cos_out\[30\] net214
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_88_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2920_ net268 _1212_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__a21o_1
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2851_ cordic_inst.cordic_inst.y\[3\] cordic_inst.cordic_inst.y\[4\] net314 VGND
+ VGND VPWR VPWR _1154_ sky130_fd_sc_hd__mux2_1
X_2782_ cordic_inst.cordic_inst.y\[27\] cordic_inst.cordic_inst.y\[28\] net305 VGND
+ VGND VPWR VPWR _1085_ sky130_fd_sc_hd__mux2_1
X_4521_ net374 _0000_ _0087_ VGND VGND VPWR VPWR cordic_inst.state\[2\] sky130_fd_sc_hd__dfrtp_1
X_4452_ net322 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__inv_2
X_3403_ _1639_ _1641_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__nand2_1
X_4383_ net321 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
X_3334_ net287 _1499_ _1571_ _1572_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__a31o_1
X_3265_ net250 net206 VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _1271_ _1270_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__nand2b_1
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4719_ net390 _0446_ _0141_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3050_ cordic_inst.cordic_inst.x\[19\] _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__nor2_1
XFILLER_82_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3952_ axi_controller.write_addr_reg\[1\] net47 net190 VGND VGND VPWR VPWR _0300_
+ sky130_fd_sc_hd__mux2_1
X_3883_ axi_controller.reg_input_data\[8\] _1964_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__or2_1
X_2903_ net244 _1130_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__nand2_1
X_2834_ _1079_ _1133_ _1135_ _1132_ net241 net235 VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__mux4_2
X_4504_ net329 VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__inv_2
X_2765_ net264 net278 VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__and2_1
X_2696_ _0842_ _1022_ _0841_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__a21bo_1
X_4435_ net334 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__inv_2
X_4366_ net344 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
XFILLER_86_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3317_ _1554_ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__or2_1
X_4297_ axi_controller.reg_input_data\[20\] _2242_ VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__or2_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3248_ net273 _0708_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ cordic_inst.cordic_inst.x\[8\] net157 _1458_ net174 VGND VGND VPWR VPWR _0506_
+ sky130_fd_sc_hd__o22a_1
XFILLER_54_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2550_ _0599_ _0882_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__nor2_1
Xoutput129 net129 VGND VGND VPWR VPWR rdata[25] sky130_fd_sc_hd__buf_2
Xoutput118 net118 VGND VGND VPWR VPWR rdata[15] sky130_fd_sc_hd__buf_2
X_2481_ _0644_ _0805_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__xnor2_1
X_4220_ cordic_inst.cordic_inst.cos_out\[22\] _2173_ net223 VGND VGND VPWR VPWR _2184_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_91_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4151_ cordic_inst.cordic_inst.sin_out\[14\] cordic_inst.cordic_inst.sin_out\[13\]
+ _2107_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__or3_1
XFILLER_83_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3102_ _1002_ _1404_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__xor2_1
XFILLER_55_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4082_ net229 _2059_ _2061_ _2062_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__a22o_1
X_3033_ _1210_ _1219_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3935_ axi_controller.read_addr_reg\[3\] axi_controller.read_addr_reg\[4\] axi_controller.read_addr_reg\[5\]
+ _1977_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__and4bb_1
X_3866_ axi_controller.write_addr_reg\[2\] axi_controller.write_addr_reg\[7\] axi_controller.write_addr_reg\[6\]
+ axi_controller.write_addr_reg\[9\] VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__or4_1
X_3797_ axi_controller.reg_input_data\[24\] _1893_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__xnor2_1
X_2817_ cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.y\[6\] net312 VGND
+ VGND VPWR VPWR _1120_ sky130_fd_sc_hd__mux2_1
X_2748_ _0873_ _0914_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nand2b_1
X_2679_ _0976_ _0979_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__or2_1
X_4418_ net338 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__inv_2
Xfanout323 net325 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__buf_4
Xfanout301 cordic_inst.cordic_inst.i\[1\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_2
Xfanout312 net315 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout356 net357 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_2
Xfanout334 net336 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_4
X_4349_ net339 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
Xfanout345 net348 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_4
Xfanout389 net392 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout378 net379 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_2
Xfanout367 net368 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ cordic_inst.deg_handler_inst.theta_norm\[16\] _1840_ VGND VGND VPWR VPWR _0015_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_13_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3651_ cordic_inst.deg_handler_inst.theta_abs\[14\] _1770_ VGND VGND VPWR VPWR _1804_
+ sky130_fd_sc_hd__nand2_1
X_2602_ net153 _0758_ _0765_ net252 VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__a31o_1
X_3582_ net289 net182 _1580_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__and3_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2533_ _0858_ _0861_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__and2b_1
X_2464_ _0789_ _0791_ _0793_ net269 VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__o31ai_1
X_4203_ cordic_inst.cordic_inst.sin_out\[20\] cordic_inst.cordic_inst.sin_out\[19\]
+ _2151_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__or3_1
X_2395_ cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.x\[6\] cordic_inst.cordic_inst.x\[7\]
+ cordic_inst.cordic_inst.x\[8\] net312 net302 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__mux4_1
X_4134_ net260 _2107_ cordic_inst.cordic_inst.sin_out\[13\] VGND VGND VPWR VPWR _2108_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4065_ cordic_inst.cordic_inst.cos_out\[3\] cordic_inst.cordic_inst.cos_out\[2\]
+ cordic_inst.cordic_inst.cos_out\[1\] cordic_inst.cordic_inst.cos_out\[0\] VGND VGND
+ VPWR VPWR _2048_ sky130_fd_sc_hd__or4_2
X_3016_ _1180_ _1185_ net271 VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4898_ net377 _0051_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_3918_ axi_controller.read_addr_reg\[19\] net12 net195 VGND VGND VPWR VPWR _0285_
+ sky130_fd_sc_hd__mux2_1
X_3849_ net63 net62 net61 VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__nand3b_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout164 net165 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout197 net198 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_4
Xfanout175 _0627_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_2
XFILLER_47_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout186 _0626_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_2
XFILLER_47_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4821_ net394 _0548_ _0243_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_61_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4752_ net399 _0479_ _0174_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3703_ net255 _1829_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__nand2_1
X_4683_ net409 _0410_ _0105_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3634_ _1762_ net147 _1795_ net151 cordic_inst.deg_handler_inst.theta_abs\[5\] VGND
+ VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3565_ cordic_inst.cordic_inst.x\[14\] cordic_inst.cordic_inst.cos_out\[14\] net214
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3496_ _1518_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2516_ _0667_ _0845_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__xor2_1
X_2447_ _0771_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nor2_1
XFILLER_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2378_ _0609_ net222 VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and2_1
X_4117_ cordic_inst.cordic_inst.sin_out\[10\] _2086_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__or2_1
XFILLER_56_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4048_ axi_controller.result_out\[1\] _2033_ net204 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3350_ net274 _1582_ _1588_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__a21boi_1
X_2301_ net233 _0634_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a21oi_1
X_3281_ _1518_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__or2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4804_ net406 _0531_ _0226_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2996_ _1297_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__and2b_1
X_4735_ net383 _0462_ _0157_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[28\] sky130_fd_sc_hd__dfrtp_1
X_4666_ net376 _0395_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[20\] sky130_fd_sc_hd__dfxtp_1
X_4597_ net361 _0329_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[30\] sky130_fd_sc_hd__dfxtp_1
X_3617_ cordic_inst.deg_handler_inst.theta_abs\[23\] _1784_ _1779_ VGND VGND VPWR
+ VPWR _1785_ sky130_fd_sc_hd__a21o_1
X_3548_ net267 cordic_inst.cordic_inst.cos_out\[31\] net208 VGND VGND VPWR VPWR _0433_
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3479_ _1632_ _1647_ _1705_ _1641_ _1645_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__o311a_1
XFILLER_28_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2850_ net288 _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__and2_1
X_2781_ cordic_inst.cordic_inst.y\[23\] cordic_inst.cordic_inst.y\[24\] cordic_inst.cordic_inst.y\[25\]
+ cordic_inst.cordic_inst.y\[26\] net306 net297 VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_41_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4520_ net374 _0007_ _0086_ VGND VGND VPWR VPWR cordic_inst.state\[1\] sky130_fd_sc_hd__dfrtp_1
X_4451_ net322 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__inv_2
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3402_ cordic_inst.cordic_inst.z\[18\] _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__xor2_1
X_4382_ net323 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
X_3333_ net242 net302 net313 net293 VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__o211a_1
X_3264_ net287 net206 _1501_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3195_ cordic_inst.cordic_inst.x\[2\] net157 _1468_ net177 VGND VGND VPWR VPWR _0500_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2979_ _1254_ _1258_ _1278_ _1252_ _1249_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__a311o_1
X_4718_ net404 _0445_ _0140_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[11\] sky130_fd_sc_hd__dfrtp_1
X_4649_ net365 _0380_ net321 VGND VGND VPWR VPWR axi_controller.result_out\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_82_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3951_ axi_controller.write_addr_reg\[0\] net36 net190 VGND VGND VPWR VPWR _0299_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2902_ net244 _1163_ _1202_ _1203_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a211o_1
X_3882_ net104 _1963_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__nand2_2
X_2833_ _1079_ _1135_ net232 VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__mux2_1
X_2764_ _0600_ _1067_ _1066_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux2_1
X_4503_ net330 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2695_ _0835_ _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__nand2_1
X_4434_ net335 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__inv_2
X_4365_ net344 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
X_3316_ cordic_inst.cordic_inst.z\[7\] _1553_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__nor2_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4296_ net81 _2243_ _2247_ net350 VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o211a_1
X_3247_ _1484_ _1485_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__or2_1
X_3178_ _1290_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__and2_1
XFILLER_25_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput108 net108 VGND VGND VPWR VPWR arready sky130_fd_sc_hd__buf_2
Xoutput119 net119 VGND VGND VPWR VPWR rdata[16] sky130_fd_sc_hd__buf_2
X_2480_ cordic_inst.cordic_inst.y\[29\] _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_91_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4150_ cordic_inst.cordic_inst.cos_out\[15\] net224 _2120_ net318 VGND VGND VPWR
+ VPWR _2122_ sky130_fd_sc_hd__a31o_1
X_3101_ _1077_ _1226_ _1227_ net270 VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__o31a_1
X_4081_ cordic_inst.cordic_inst.sin_out\[6\] _2060_ net230 VGND VGND VPWR VPWR _2062_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_83_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3032_ cordic_inst.cordic_inst.x\[23\] _1334_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3934_ axi_controller.read_addr_reg\[1\] axi_controller.read_addr_reg\[0\] axi_controller.read_addr_reg\[7\]
+ axi_controller.read_addr_reg\[6\] VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__nor4_1
X_3865_ _1944_ _1945_ _1946_ _1947_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__or4_1
X_2816_ _1117_ _1118_ net291 VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__mux2_1
X_3796_ axi_controller.reg_input_data\[23\] _1890_ _1874_ VGND VGND VPWR VPWR _1896_
+ sky130_fd_sc_hd__o21ba_1
X_2747_ _0873_ _0874_ _0878_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__o211ai_1
X_2678_ net178 _0997_ _1009_ net158 cordic_inst.cordic_inst.y\[28\] VGND VGND VPWR
+ VPWR _0558_ sky130_fd_sc_hd__a32o_1
X_4417_ net337 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
Xfanout302 net304 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_4
Xfanout313 net315 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__buf_2
Xfanout346 net347 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__buf_4
Xfanout357 net358 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout324 net325 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_2
Xfanout335 net336 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_4
X_4348_ net337 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
Xfanout379 net382 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_2
Xfanout368 net369 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlymetal6s2s_1
X_4279_ net199 _2235_ _2230_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3650_ _1770_ _1790_ _1803_ net151 cordic_inst.deg_handler_inst.theta_abs\[13\] VGND
+ VGND VPWR VPWR _0057_ sky130_fd_sc_hd__a32o_1
X_2601_ _0926_ _0930_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__nand3b_1
X_3581_ cordic_inst.cordic_inst.start cordic_inst.state\[2\] _0620_ _0618_ VGND VGND
+ VPWR VPWR _0400_ sky130_fd_sc_hd__o211a_1
X_2532_ _0844_ _0864_ _0865_ _0832_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__o221a_1
X_4202_ cordic_inst.cordic_inst.cos_out\[21\] net225 _2166_ net318 VGND VGND VPWR
+ VPWR _2168_ sky130_fd_sc_hd__a31oi_1
X_2463_ net278 _0766_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nor2_1
X_2394_ cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.x\[6\] net312 VGND
+ VGND VPWR VPWR _0729_ sky130_fd_sc_hd__mux2_1
XFILLER_68_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4133_ cordic_inst.cordic_inst.sin_out\[12\] _2099_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__or2_1
XFILLER_56_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4064_ net262 _2045_ cordic_inst.cordic_inst.sin_out\[4\] VGND VGND VPWR VPWR _2047_
+ sky130_fd_sc_hd__a21oi_1
X_3015_ _1316_ _1317_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_54_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4897_ net381 _0050_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_3917_ axi_controller.read_addr_reg\[18\] net11 net195 VGND VGND VPWR VPWR _0284_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3848_ net350 _1931_ _1930_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a21o_1
X_3779_ axi_controller.reg_input_data\[20\] _1882_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout154 _2256_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xfanout165 net168 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout198 _1926_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
Xfanout187 _1929_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_4
Xfanout176 _0627_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4820_ net395 _0547_ _0242_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4751_ net400 _0478_ _0173_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3702_ cordic_inst.deg_handler_inst.theta_norm\[9\] _1827_ VGND VGND VPWR VPWR _1829_
+ sky130_fd_sc_hd__or2_1
X_4682_ net409 _0409_ _0104_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3633_ cordic_inst.deg_handler_inst.theta_abs\[5\] _1761_ VGND VGND VPWR VPWR _1795_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3564_ cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.cos_out\[15\] net210
+ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
X_3495_ _1520_ _1717_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__nor2_1
X_2515_ _0849_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__inv_2
X_2446_ _0672_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__nand2_1
X_2377_ net303 net314 VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__or2_1
XFILLER_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4116_ net203 _2092_ _2085_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4047_ _2030_ _2032_ net229 VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4949_ net398 _0578_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3280_ cordic_inst.cordic_inst.z\[14\] _1517_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__nor2_1
X_2300_ net265 net295 VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__and2_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4803_ net406 _0530_ _0225_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[0\] sky130_fd_sc_hd__dfrtp_1
X_2995_ cordic_inst.cordic_inst.x\[15\] _1296_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__nand2_1
X_4734_ net383 _0461_ _0156_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4665_ net376 _0394_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[19\] sky130_fd_sc_hd__dfxtp_2
X_3616_ _1782_ _1783_ _0617_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__o21ai_1
X_4596_ net361 _0328_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[29\] sky130_fd_sc_hd__dfxtp_1
X_3547_ cordic_inst.cordic_inst.angle\[0\] net172 net165 cordic_inst.cordic_inst.z\[0\]
+ _1754_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a221o_1
XFILLER_88_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3478_ _1629_ _1634_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__and2_1
X_2429_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__inv_2
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ cordic_inst.cordic_inst.y\[25\] cordic_inst.cordic_inst.y\[26\] net305 VGND
+ VGND VPWR VPWR _1083_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4450_ net322 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__inv_2
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4381_ net323 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
X_3401_ net251 _1508_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__xnor2_1
X_3332_ net313 _0705_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__nor2_1
X_3263_ net293 net303 net313 VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__nor3_1
X_3194_ _1274_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2978_ _1254_ _1258_ _1278_ _1252_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__a31o_1
X_4717_ net405 _0444_ _0139_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[10\] sky130_fd_sc_hd__dfrtp_1
X_4648_ net365 _0379_ net321 VGND VGND VPWR VPWR axi_controller.result_out\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4579_ net361 _0311_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3950_ axi_controller.done _1992_ net351 _0085_ _1918_ VGND VGND VPWR VPWR _0298_
+ sky130_fd_sc_hd__o2111a_1
X_2901_ net244 _1163_ _1068_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__a21o_1
XFILLER_50_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3881_ net104 _1963_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__and2_1
X_2832_ cordic_inst.cordic_inst.y\[24\] cordic_inst.cordic_inst.y\[25\] cordic_inst.cordic_inst.y\[26\]
+ cordic_inst.cordic_inst.y\[27\] net305 net296 VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__mux4_1
X_2763_ _0600_ net171 VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nor2_1
X_4502_ net330 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__inv_2
X_2694_ _0864_ _0973_ _0837_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a21o_1
X_4433_ net336 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__inv_2
X_4364_ net344 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
X_3315_ cordic_inst.cordic_inst.z\[7\] _1553_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__and2_1
X_4295_ axi_controller.reg_input_data\[19\] _2242_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__or2_1
X_3246_ _1481_ _1483_ cordic_inst.cordic_inst.z\[21\] VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__a21oi_1
X_3177_ _1284_ _1289_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__nand2_1
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput109 net109 VGND VGND VPWR VPWR awready sky130_fd_sc_hd__buf_2
XFILLER_49_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3100_ _1236_ _1238_ _1401_ _1234_ _1231_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__a311oi_1
X_4080_ cordic_inst.cordic_inst.sin_out\[6\] _2060_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__or2_1
XFILLER_83_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3031_ _1220_ _1333_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__xnor2_1
X_3933_ _1974_ _1975_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__nor2_1
X_3864_ axi_controller.write_addr_reg\[24\] axi_controller.write_addr_reg\[27\] axi_controller.write_addr_reg\[26\]
+ axi_controller.write_addr_reg\[28\] VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__or4b_1
X_2815_ cordic_inst.cordic_inst.y\[17\] cordic_inst.cordic_inst.y\[18\] cordic_inst.cordic_inst.y\[19\]
+ cordic_inst.cordic_inst.y\[20\] net308 net298 VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__mux4_1
X_3795_ _1891_ _1895_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2746_ _0876_ _0879_ _0913_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__or3b_1
X_2677_ _0821_ _0996_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__nand2_1
X_4416_ net337 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__inv_2
Xfanout303 net304 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_2
Xfanout314 net315 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__buf_2
Xfanout347 net348 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__buf_4
Xfanout325 net328 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
Xfanout336 net349 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_2
X_4347_ net337 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
XFILLER_59_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4278_ net316 _2231_ _2232_ _2233_ _2234_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__o32a_1
Xfanout358 net359 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout369 net414 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_2
XFILLER_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3229_ cordic_inst.cordic_inst.y\[4\] cordic_inst.cordic_inst.sin_out\[4\] net212
+ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2600_ _0933_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__nor2_1
X_3580_ cordic_inst.cordic_inst.done cordic_inst.cordic_inst.state\[0\] cordic_inst.cordic_inst.state\[1\]
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o21a_1
X_2531_ _0823_ _0828_ _0829_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a21o_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4201_ net225 _2166_ cordic_inst.cordic_inst.cos_out\[21\] VGND VGND VPWR VPWR _2167_
+ sky130_fd_sc_hd__a21o_1
X_2462_ net243 _0676_ net169 VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__a21o_1
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2393_ _0726_ _0727_ net295 VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__mux2_1
X_4132_ _2102_ _2106_ axi_controller.result_out\[12\] net201 VGND VGND VPWR VPWR _0366_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4063_ cordic_inst.cordic_inst.sin_out\[4\] net262 _2045_ VGND VGND VPWR VPWR _2046_
+ sky130_fd_sc_hd__and3_1
XFILLER_68_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3014_ cordic_inst.cordic_inst.x\[11\] _1315_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__nand2_1
XFILLER_36_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4965_ net371 _0594_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_1
X_3916_ axi_controller.read_addr_reg\[17\] net10 net195 VGND VGND VPWR VPWR _0283_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4896_ net381 _0049_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_3847_ axi_controller.state\[0\] net68 net107 _1920_ axi_controller.state\[2\] VGND
+ VGND VPWR VPWR _1931_ sky130_fd_sc_hd__a32o_1
X_3778_ _1874_ _1880_ axi_controller.reg_input_data\[19\] VGND VGND VPWR VPWR _1882_
+ sky130_fd_sc_hd__mux2_1
X_2729_ net181 _1043_ _1046_ net162 cordic_inst.cordic_inst.y\[14\] VGND VGND VPWR
+ VPWR _0544_ sky130_fd_sc_hd__a32o_1
XFILLER_3_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout155 _2256_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xfanout199 net205 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
Xfanout188 _1929_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
Xfanout177 _0627_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
Xfanout166 net168 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4750_ net400 _0477_ _0172_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3701_ cordic_inst.deg_handler_inst.theta_norm\[9\] _1828_ VGND VGND VPWR VPWR _0039_
+ sky130_fd_sc_hd__xnor2_1
X_4681_ net410 _0408_ _0103_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3632_ _1761_ net147 _1794_ net152 cordic_inst.deg_handler_inst.theta_abs\[4\] VGND
+ VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a32o_1
X_3563_ cordic_inst.cordic_inst.x\[16\] cordic_inst.cordic_inst.cos_out\[16\] net210
+ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
X_3494_ _1515_ _1627_ _1530_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__a21o_1
X_2514_ cordic_inst.cordic_inst.y\[19\] _0847_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__xor2_1
XFILLER_5_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2445_ _0776_ _0777_ _0779_ _0773_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4115_ net229 _2087_ _2088_ _2090_ _2091_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__o32a_1
X_2376_ net304 net312 VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nor2_2
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4046_ cordic_inst.cordic_inst.cos_out\[1\] _2031_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4948_ net398 _0577_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4879_ net388 axi_controller.reg_input_data\[11\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2994_ cordic_inst.cordic_inst.x\[15\] _1296_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__nor2_1
X_4802_ net369 _0529_ _0224_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4733_ net383 _0460_ _0155_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[26\] sky130_fd_sc_hd__dfrtp_1
X_4664_ net376 _0393_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[18\] sky130_fd_sc_hd__dfxtp_1
X_4595_ net362 _0327_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[28\] sky130_fd_sc_hd__dfxtp_1
X_3615_ cordic_inst.deg_handler_inst.theta_abs\[20\] cordic_inst.deg_handler_inst.theta_abs\[21\]
+ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__nand2_1
X_3546_ _1597_ _1753_ net183 VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__o21a_1
X_3477_ _1703_ _1704_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__nand2_1
X_2428_ _0760_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__or2_1
XFILLER_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2359_ cordic_inst.cordic_inst.x\[16\] cordic_inst.cordic_inst.x\[17\] cordic_inst.cordic_inst.x\[18\]
+ cordic_inst.cordic_inst.x\[19\] net308 net298 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__mux4_1
XFILLER_56_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4029_ axi_controller.reg_input_data\[2\] _2018_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__or2_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4380_ net323 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
X_3400_ _1637_ _1638_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__and2_1
X_3331_ _1568_ _1569_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__nor2_1
X_3262_ _1499_ _1500_ net287 VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__a21oi_1
X_3193_ _1269_ _1272_ _1273_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__nand3_1
XFILLER_66_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2977_ _1252_ _1253_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__or2_1
X_4716_ net405 _0443_ _0138_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[9\] sky130_fd_sc_hd__dfrtp_1
X_4647_ net367 _0378_ net323 VGND VGND VPWR VPWR axi_controller.result_out\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4578_ net370 _0310_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[11\] sky130_fd_sc_hd__dfxtp_1
X_3529_ cordic_inst.cordic_inst.angle\[6\] net172 net167 cordic_inst.cordic_inst.z\[6\]
+ _1742_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a221o_1
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2900_ net279 _1168_ _1069_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3880_ _0622_ _1962_ _1943_ _1922_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__and4bb_4
X_2831_ _1132_ _1133_ net291 VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__mux2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2762_ net184 _0718_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__nand2_1
X_4501_ net335 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__inv_2
X_2693_ cordic_inst.cordic_inst.y\[24\] net159 _1019_ _1020_ VGND VGND VPWR VPWR _0554_
+ sky130_fd_sc_hd__a22o_1
X_4432_ net336 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__inv_2
X_4363_ net344 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
X_3314_ net275 _1481_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__mux2_1
X_4294_ net80 _2243_ _2246_ net353 VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__o211a_1
X_3245_ cordic_inst.cordic_inst.z\[21\] _1481_ _1483_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__and3_1
XFILLER_39_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ cordic_inst.cordic_inst.x\[9\] net157 _1455_ _1456_ VGND VGND VPWR VPWR _0507_
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3030_ net215 _1090_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__or2_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3932_ axi_controller.read_addr_reg\[9\] axi_controller.read_addr_reg\[8\] axi_controller.read_addr_reg\[11\]
+ axi_controller.read_addr_reg\[10\] VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__or4_1
X_3863_ axi_controller.write_addr_reg\[29\] axi_controller.write_addr_reg\[30\] axi_controller.write_addr_reg\[31\]
+ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__nand3_1
X_2814_ cordic_inst.cordic_inst.y\[13\] cordic_inst.cordic_inst.y\[14\] cordic_inst.cordic_inst.y\[15\]
+ cordic_inst.cordic_inst.y\[16\] net308 net298 VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__mux4_1
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3794_ axi_controller.reg_input_data\[23\] _1880_ _1894_ VGND VGND VPWR VPWR _1895_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2745_ net181 _1037_ _1056_ net161 cordic_inst.cordic_inst.y\[8\] VGND VGND VPWR
+ VPWR _0538_ sky130_fd_sc_hd__a32o_1
X_2676_ cordic_inst.cordic_inst.y\[29\] net158 _1008_ net178 VGND VGND VPWR VPWR _0559_
+ sky130_fd_sc_hd__a22o_1
X_4415_ net338 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
Xfanout304 cordic_inst.cordic_inst.i\[1\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__buf_2
X_4346_ net253 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
Xfanout326 net328 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__buf_4
Xfanout337 net338 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_4
Xfanout315 cordic_inst.cordic_inst.i\[0\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_2
Xfanout348 net349 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_4
X_4277_ cordic_inst.cordic_inst.sin_out\[30\] net258 _2224_ net228 VGND VGND VPWR
+ VPWR _2234_ sky130_fd_sc_hd__a31o_1
Xfanout359 net364 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__buf_2
X_3228_ cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.sin_out\[5\] net211
+ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
X_3159_ _1302_ _1445_ _1299_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ _0835_ _0841_ _0842_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__a21bo_1
X_2461_ _0637_ _0761_ net280 VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__a21oi_1
X_4200_ cordic_inst.cordic_inst.cos_out\[20\] cordic_inst.cordic_inst.cos_out\[19\]
+ _2155_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__or3_1
X_2392_ cordic_inst.cordic_inst.x\[13\] cordic_inst.cordic_inst.x\[14\] cordic_inst.cordic_inst.x\[15\]
+ cordic_inst.cordic_inst.x\[16\] net309 net299 VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_79_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4131_ _2104_ _2105_ net201 VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__o21a_1
X_4062_ cordic_inst.cordic_inst.sin_out\[3\] cordic_inst.cordic_inst.sin_out\[2\]
+ cordic_inst.cordic_inst.sin_out\[1\] cordic_inst.cordic_inst.sin_out\[0\] VGND VGND
+ VPWR VPWR _2045_ sky130_fd_sc_hd__or4_2
X_3013_ cordic_inst.cordic_inst.x\[11\] _1315_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nor2_1
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4964_ net413 _0593_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_88_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3915_ axi_controller.read_addr_reg\[16\] net9 net195 VGND VGND VPWR VPWR _0282_
+ sky130_fd_sc_hd__mux2_1
X_4895_ net378 _0048_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3846_ net350 net107 axi_controller.state\[3\] VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__and3_1
X_3777_ axi_controller.reg_input_data\[19\] _1881_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__xor2_1
X_2728_ _0925_ _1042_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__nand2_1
X_2659_ _0984_ _0986_ _0989_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__nand4_1
X_4329_ net117 net192 net155 axi_controller.result_out\[14\] VGND VGND VPWR VPWR _0580_
+ sky130_fd_sc_hd__a22o_1
Xfanout156 _2256_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
Xfanout178 net186 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_4
Xfanout189 _1929_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3700_ net255 _1827_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__nand2_1
XFILLER_14_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4680_ net410 _0407_ _0102_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3631_ cordic_inst.deg_handler_inst.theta_abs\[4\] _1760_ VGND VGND VPWR VPWR _1794_
+ sky130_fd_sc_hd__nand2_1
X_3562_ cordic_inst.cordic_inst.x\[17\] cordic_inst.cordic_inst.cos_out\[17\] net209
+ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
X_2513_ cordic_inst.cordic_inst.y\[19\] _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nor2_1
X_3493_ cordic_inst.cordic_inst.angle\[16\] net173 net165 cordic_inst.cordic_inst.z\[16\]
+ _1716_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a221o_1
X_2444_ _0601_ _0636_ _0691_ _0686_ net240 net247 VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__mux4_2
X_2375_ cordic_inst.cordic_inst.x\[2\] cordic_inst.cordic_inst.x\[3\] net312 VGND
+ VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux2_1
X_4114_ cordic_inst.cordic_inst.cos_out\[10\] net226 _2089_ net319 VGND VGND VPWR
+ VPWR _2091_ sky130_fd_sc_hd__a31o_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4045_ cordic_inst.cordic_inst.cos_out\[0\] net227 VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4947_ net396 _0576_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4878_ net388 axi_controller.reg_input_data\[10\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3829_ cordic_inst.sign_handler_inst.done_d cordic_inst.cordic_inst.done VGND VGND
+ VPWR VPWR cordic_inst.sign_handler_inst.done_pulse sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_30_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2993_ _1198_ _1216_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__xnor2_1
X_4801_ net369 _0528_ _0223_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[30\] sky130_fd_sc_hd__dfrtp_2
X_4732_ net384 _0459_ _0154_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[25\] sky130_fd_sc_hd__dfrtp_1
X_4663_ net376 _0392_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[17\] sky130_fd_sc_hd__dfxtp_1
X_3614_ cordic_inst.deg_handler_inst.theta_abs\[18\] cordic_inst.deg_handler_inst.theta_abs\[19\]
+ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__nor2_1
X_4594_ net362 _0326_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[27\] sky130_fd_sc_hd__dfxtp_1
X_3545_ cordic_inst.cordic_inst.z\[0\] _1583_ _1584_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__and3_1
X_3476_ cordic_inst.cordic_inst.angle\[20\] net170 net164 cordic_inst.cordic_inst.z\[20\]
+ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__a22oi_1
X_2427_ net265 _0721_ _0724_ _0728_ net247 net240 VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__mux4_1
X_2358_ net247 _0692_ _0689_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2289_ axi_controller.read_addr_reg\[31\] VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__inv_2
XFILLER_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4028_ net82 _2019_ _2021_ net354 VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__o211a_1
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3330_ cordic_inst.cordic_inst.z\[5\] _1567_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__nor2_1
X_3261_ net303 net313 VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__nand2_1
XFILLER_85_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3192_ net184 _1277_ _1466_ net166 cordic_inst.cordic_inst.x\[3\] VGND VGND VPWR
+ VPWR _0501_ sky130_fd_sc_hd__a32o_1
XFILLER_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2976_ _1258_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__nand2_1
X_4715_ net405 _0442_ _0137_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[8\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_15_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4646_ net393 _0377_ net323 VGND VGND VPWR VPWR axi_controller.result_out\[23\] sky130_fd_sc_hd__dfrtp_1
X_4577_ net370 _0309_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3528_ _1563_ _1607_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__a21oi_1
X_3459_ cordic_inst.cordic_inst.angle\[24\] net171 net163 cordic_inst.cordic_inst.z\[24\]
+ _1690_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__a221o_1
XFILLER_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2830_ cordic_inst.cordic_inst.y\[20\] cordic_inst.cordic_inst.y\[21\] cordic_inst.cordic_inst.y\[22\]
+ cordic_inst.cordic_inst.y\[23\] net308 net298 VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_51_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2761_ net184 _0898_ _1065_ net166 cordic_inst.cordic_inst.y\[1\] VGND VGND VPWR
+ VPWR _0531_ sky130_fd_sc_hd__a32o_1
X_2692_ net174 _0979_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__nor2_1
X_4500_ net349 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__inv_2
X_4431_ net342 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__inv_2
XANTENNA_1 _2028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4362_ net344 VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
X_4293_ axi_controller.reg_input_data\[18\] _2242_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__or2_1
X_3313_ net287 _0707_ _1521_ _1510_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_60_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3244_ _1482_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__inv_2
XFILLER_39_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _1295_ _1439_ net175 VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__a21o_1
XFILLER_81_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2959_ _1169_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__xor2_1
X_4629_ net410 _0360_ net343 VGND VGND VPWR VPWR axi_controller.result_out\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3931_ axi_controller.read_addr_reg\[13\] axi_controller.read_addr_reg\[12\] axi_controller.read_addr_reg\[15\]
+ axi_controller.read_addr_reg\[14\] VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__or4_1
X_3862_ axi_controller.write_addr_reg\[16\] axi_controller.write_addr_reg\[19\] axi_controller.write_addr_reg\[18\]
+ axi_controller.write_addr_reg\[21\] VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__or4_1
X_2813_ net245 _1115_ _1110_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__o21ai_2
X_3793_ axi_controller.reg_input_data\[23\] _1892_ _1893_ VGND VGND VPWR VPWR _1894_
+ sky130_fd_sc_hd__o21a_1
X_2744_ _0915_ _0959_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nand2_1
X_2675_ _0998_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__xnor2_1
X_4414_ net338 VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__inv_2
Xfanout305 net306 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_4
X_4345_ cordic_inst.deg_handler_inst.theta_abs\[31\] VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
Xfanout316 net320 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_2
Xfanout327 net328 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_4
Xfanout338 net341 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__buf_2
X_4276_ net258 _2224_ cordic_inst.cordic_inst.sin_out\[30\] VGND VGND VPWR VPWR _2233_
+ sky130_fd_sc_hd__a21oi_1
Xfanout349 axi_controller.rst VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3227_ cordic_inst.cordic_inst.y\[6\] cordic_inst.cordic_inst.sin_out\[6\] net211
+ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux2_1
X_3158_ _1303_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nand2_1
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3089_ _1222_ _1391_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2460_ net243 _0759_ net169 VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21o_1
XFILLER_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4130_ cordic_inst.cordic_inst.cos_out\[12\] net225 _2103_ net318 VGND VGND VPWR
+ VPWR _2105_ sky130_fd_sc_hd__a31o_1
X_2391_ cordic_inst.cordic_inst.x\[9\] cordic_inst.cordic_inst.x\[10\] cordic_inst.cordic_inst.x\[11\]
+ cordic_inst.cordic_inst.x\[12\] net309 net299 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__mux4_1
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4061_ axi_controller.result_out\[4\] net204 VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__nor2_1
XFILLER_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3012_ _1098_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4963_ net412 _0592_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
X_3914_ axi_controller.read_addr_reg\[15\] net8 net198 VGND VGND VPWR VPWR _0281_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4894_ net372 _0047_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3845_ net350 _0622_ axi_controller.state\[3\] net190 VGND VGND VPWR VPWR _0004_
+ sky130_fd_sc_hd__a31o_1
X_3776_ _1874_ _1880_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__nand2_1
X_2727_ cordic_inst.cordic_inst.y\[15\] net162 _1045_ net181 VGND VGND VPWR VPWR _0545_
+ sky130_fd_sc_hd__a22o_1
X_2658_ cordic_inst.cordic_inst.y\[25\] _0988_ _0976_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a21o_1
X_2589_ cordic_inst.cordic_inst.y\[14\] _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__nand2_1
X_4328_ net118 net192 net155 axi_controller.result_out\[15\] VGND VGND VPWR VPWR _0579_
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4259_ cordic_inst.deg_handler_inst.kuadran\[0\] _2211_ VGND VGND VPWR VPWR _2218_
+ sky130_fd_sc_hd__nor2_1
Xfanout179 net186 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
Xfanout168 _0629_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
Xfanout157 cordic_inst.cordic_inst.next_state\[1\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3630_ _1760_ _1790_ _1793_ net152 cordic_inst.deg_handler_inst.theta_abs\[3\] VGND
+ VGND VPWR VPWR _0078_ sky130_fd_sc_hd__a32o_1
X_3561_ cordic_inst.cordic_inst.x\[18\] cordic_inst.cordic_inst.cos_out\[18\] net209
+ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
X_2512_ _0666_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3492_ _1629_ _1634_ _1715_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__o21a_1
X_2443_ _0776_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nor2_1
X_2374_ net288 net295 net302 VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nor3b_2
X_4113_ net226 _2089_ cordic_inst.cordic_inst.cos_out\[10\] VGND VGND VPWR VPWR _2090_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_67_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4044_ cordic_inst.cordic_inst.sin_out\[1\] _2029_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4946_ net396 _0575_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4877_ net388 axi_controller.reg_input_data\[9\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3828_ _0618_ _1918_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3759_ axi_controller.reg_input_data\[11\] axi_controller.reg_input_data\[10\] axi_controller.reg_input_data\[9\]
+ axi_controller.reg_input_data\[8\] VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__or4_1
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4800_ net369 _0527_ _0222_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_61_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2992_ _1293_ _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__nand2b_1
X_4731_ net384 _0458_ _0153_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[24\] sky130_fd_sc_hd__dfrtp_1
X_4662_ net376 _0391_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[16\] sky130_fd_sc_hd__dfxtp_1
X_3613_ cordic_inst.deg_handler_inst.theta_abs\[31\] _1780_ VGND VGND VPWR VPWR _1781_
+ sky130_fd_sc_hd__or2_1
X_4593_ net360 _0325_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[26\] sky130_fd_sc_hd__dfxtp_1
X_3544_ cordic_inst.cordic_inst.angle\[1\] net172 net165 cordic_inst.cordic_inst.z\[1\]
+ _1752_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__a221o_1
X_3475_ _1490_ _1650_ _1654_ _1702_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__a31o_1
X_2426_ net240 _0724_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nand2_1
XFILLER_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2357_ net266 _0634_ _0657_ _0654_ net233 net240 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__mux4_2
XFILLER_84_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2288_ axi_controller.state\[3\] VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__inv_2
XFILLER_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4027_ axi_controller.reg_input_data\[1\] _2018_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__or2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4929_ net373 _0029_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3260_ net293 net303 VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__nand2_1
X_3191_ _1266_ _1274_ _1276_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_77_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4714_ net405 _0441_ _0136_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[7\] sky130_fd_sc_hd__dfrtp_1
X_2975_ _1263_ _1277_ _1260_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a21o_1
X_4645_ net367 _0376_ net324 VGND VGND VPWR VPWR axi_controller.result_out\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4576_ net370 _0308_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[9\] sky130_fd_sc_hd__dfxtp_1
X_3527_ net176 _1608_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__or2_1
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3458_ _1689_ net182 _1658_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__and3b_1
X_3389_ _1625_ _1626_ _1529_ _1533_ _1535_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__a2111o_1
XFILLER_69_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2409_ _0694_ _0701_ net236 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2760_ _0896_ _0897_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nand2_1
X_2691_ _0974_ _0978_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__nand2_1
XFILLER_8_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4430_ net342 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__inv_2
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4361_ net343 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
X_3312_ _1550_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__inv_2
X_4292_ net79 _2243_ _2245_ net353 VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o211a_1
X_3243_ net273 _0714_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _1295_ _1439_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__nor2_1
XFILLER_81_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ _1148_ _1157_ _1164_ net276 VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__o31a_1
X_2889_ net263 _1127_ _1129_ _1119_ net243 net239 VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__mux4_2
X_4628_ net410 _0359_ net343 VGND VGND VPWR VPWR axi_controller.result_out\[5\] sky130_fd_sc_hd__dfrtp_1
X_4559_ net357 _0291_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3930_ axi_controller.read_addr_reg\[31\] net26 net197 VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3861_ axi_controller.write_addr_reg\[20\] axi_controller.write_addr_reg\[23\] axi_controller.write_addr_reg\[22\]
+ axi_controller.write_addr_reg\[25\] VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__or4_1
X_3792_ axi_controller.reg_input_data\[23\] _1892_ _1880_ VGND VGND VPWR VPWR _1893_
+ sky130_fd_sc_hd__a21oi_1
X_2812_ net263 _1074_ _1113_ _1111_ net232 net239 VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__mux4_2
X_2743_ net181 _1054_ _1055_ net161 cordic_inst.cordic_inst.y\[9\] VGND VGND VPWR
+ VPWR _0539_ sky130_fd_sc_hd__a32o_1
X_2674_ _0817_ _0997_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__and2b_1
X_4413_ net339 VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__inv_2
X_4344_ _2257_ net112 net194 VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux2_1
Xfanout317 net320 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout306 net307 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_4
Xfanout328 net349 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 net341 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__buf_4
X_4275_ net223 _2227_ cordic_inst.cordic_inst.cos_out\[30\] VGND VGND VPWR VPWR _2232_
+ sky130_fd_sc_hd__a21oi_1
X_3226_ cordic_inst.cordic_inst.y\[7\] cordic_inst.cordic_inst.sin_out\[7\] net211
+ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
X_3157_ _1326_ _1443_ _1307_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__o21a_1
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3088_ net215 _1212_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__or2_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2390_ _0721_ _0724_ net284 VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__mux2_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4060_ axi_controller.result_out\[3\] _2043_ net204 VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
XFILLER_76_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3011_ _1180_ _1185_ _1187_ net271 VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o31a_1
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4962_ net412 _0591_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3913_ axi_controller.read_addr_reg\[14\] net7 net198 VGND VGND VPWR VPWR _0280_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4893_ net371 _0046_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_3844_ axi_controller.state\[0\] net350 net68 _0622_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_62_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3775_ axi_controller.reg_input_data\[31\] _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__nand2_2
X_2726_ _0920_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__xnor2_1
X_2657_ _0979_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__nand2_1
X_2588_ _0779_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__xor2_2
XFILLER_86_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout147 _1790_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
X_4327_ net119 net192 net155 axi_controller.result_out\[16\] VGND VGND VPWR VPWR _0578_
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4258_ axi_controller.result_out\[27\] net199 _2216_ _2217_ VGND VGND VPWR VPWR _0381_
+ sky130_fd_sc_hd__o22a_1
Xfanout169 _0630_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_2
Xfanout158 net159 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_2
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3209_ cordic_inst.cordic_inst.y\[24\] cordic_inst.cordic_inst.sin_out\[24\] net208
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_1
X_4189_ cordic_inst.cordic_inst.cos_out\[19\] net225 _2155_ net318 VGND VGND VPWR
+ VPWR _2157_ sky130_fd_sc_hd__a31o_1
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3560_ cordic_inst.cordic_inst.x\[19\] cordic_inst.cordic_inst.cos_out\[19\] net209
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ _0667_ _0787_ net272 VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o21a_1
X_3491_ net176 _1705_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__nor2_1
X_2442_ net284 _0754_ _0637_ net278 VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__o211a_1
X_2373_ net289 net295 net304 net315 VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nor4b_1
X_4112_ cordic_inst.cordic_inst.cos_out\[9\] cordic_inst.cordic_inst.cos_out\[8\]
+ cordic_inst.cordic_inst.cos_out\[7\] _2068_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__or4_2
X_4043_ cordic_inst.cordic_inst.sin_out\[0\] net262 VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4945_ net395 _0574_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4876_ net388 axi_controller.reg_input_data\[8\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3827_ axi_controller.reg_done_flag axi_controller.start_pulse_reg VGND VGND VPWR
+ VPWR _1918_ sky130_fd_sc_hd__nand2b_1
XFILLER_20_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3758_ cordic_inst.deg_handler_inst.theta_norm\[30\] cordic_inst.deg_handler_inst.theta_norm\[29\]
+ _1861_ net253 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and4bb_1
X_2709_ _0850_ _0852_ _1030_ net175 VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__a31o_1
X_3689_ cordic_inst.deg_handler_inst.theta_norm\[4\] _1819_ net256 VGND VGND VPWR
+ VPWR _1821_ sky130_fd_sc_hd__o21ai_1
XFILLER_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ _1292_ cordic_inst.cordic_inst.x\[9\] VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__nand2b_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4730_ net386 _0457_ _0152_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[23\] sky130_fd_sc_hd__dfrtp_1
X_4661_ net385 cordic_inst.cordic_inst.done net339 VGND VGND VPWR VPWR cordic_inst.sign_handler_inst.done_d
+ sky130_fd_sc_hd__dfrtp_1
X_3612_ cordic_inst.deg_handler_inst.theta_abs\[22\] _1776_ _1779_ cordic_inst.deg_handler_inst.theta_abs\[23\]
+ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__a211oi_1
X_4592_ net360 _0324_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[25\] sky130_fd_sc_hd__dfxtp_1
X_3543_ _1597_ _1598_ _1751_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__a21oi_1
X_3474_ net182 _1691_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__nand2_1
X_2425_ net266 _0696_ _0698_ _0702_ net247 net242 VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__mux4_1
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2356_ net233 _0657_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2287_ axi_controller.write_addr_reg\[4\] VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__inv_2
XFILLER_84_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4026_ net71 _2019_ _2020_ net355 VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_35_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4928_ net373 _0028_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4859_ net384 _0068_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3190_ cordic_inst.cordic_inst.x\[4\] net157 _1465_ net177 VGND VGND VPWR VPWR _0502_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_77_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2974_ _1266_ _1274_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a21o_1
X_4713_ net405 _0440_ _0135_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[6\] sky130_fd_sc_hd__dfrtp_1
X_4644_ net393 _0375_ net329 VGND VGND VPWR VPWR axi_controller.result_out\[21\] sky130_fd_sc_hd__dfrtp_1
X_4575_ net361 _0307_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3526_ cordic_inst.cordic_inst.angle\[7\] net173 net167 cordic_inst.cordic_inst.z\[7\]
+ _1740_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__a221o_1
X_3457_ _1480_ _1655_ _1657_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__and3_1
X_3388_ _1625_ _1626_ _1535_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__a21o_1
XFILLER_69_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2408_ _0718_ _0735_ _0738_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nor4b_2
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2339_ cordic_inst.cordic_inst.x\[14\] cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.x\[16\]
+ cordic_inst.cordic_inst.x\[17\] net310 net300 VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4009_ axi_controller.reg_input_data\[25\] _2008_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2690_ net178 _1017_ _1018_ net159 cordic_inst.cordic_inst.y\[25\] VGND VGND VPWR
+ VPWR _0555_ sky130_fd_sc_hd__a32o_1
XANTENNA_3 net320 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4360_ net343 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
X_3311_ cordic_inst.cordic_inst.z\[9\] _1549_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__or2_1
X_4291_ axi_controller.reg_input_data\[17\] _2242_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__or2_1
X_3242_ net274 _0714_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__nand2_2
X_3173_ net181 _1441_ _1454_ net161 cordic_inst.cordic_inst.x\[10\] VGND VGND VPWR
+ VPWR _0508_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_1_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2957_ _1257_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__or2_1
X_2888_ net238 _1129_ _1070_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__a21boi_1
X_4627_ net410 _0358_ net344 VGND VGND VPWR VPWR axi_controller.result_out\[4\] sky130_fd_sc_hd__dfrtp_1
X_4558_ net359 _0290_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[24\] sky130_fd_sc_hd__dfxtp_1
X_3509_ cordic_inst.cordic_inst.angle\[12\] net173 net165 cordic_inst.cordic_inst.z\[12\]
+ _1728_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a221o_1
X_4489_ net346 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__inv_2
XFILLER_85_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3860_ axi_controller.state\[0\] axi_controller.state\[3\] VGND VGND VPWR VPWR _1943_
+ sky130_fd_sc_hd__or2_1
X_3791_ axi_controller.reg_input_data\[22\] axi_controller.reg_input_data\[21\] _1883_
+ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__or3_1
X_2811_ _1111_ _1113_ net291 VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__mux2_1
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2742_ _0957_ _1037_ _0955_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__a21o_1
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2673_ net178 _1000_ _1006_ net158 cordic_inst.cordic_inst.y\[30\] VGND VGND VPWR
+ VPWR _0560_ sky130_fd_sc_hd__a32o_1
X_4412_ net340 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__inv_2
X_4343_ axi_controller.reg_done_flag _1990_ _2254_ axi_controller.result_out\[0\]
+ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__a22o_1
Xfanout329 net333 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_4
Xfanout318 net319 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_4
X_4274_ cordic_inst.cordic_inst.cos_out\[30\] net223 _2227_ VGND VGND VPWR VPWR _2231_
+ sky130_fd_sc_hd__and3_1
Xfanout307 net311 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_4
X_3225_ cordic_inst.cordic_inst.y\[8\] cordic_inst.cordic_inst.sin_out\[8\] net213
+ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3156_ _1311_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__nor2_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3087_ _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__inv_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3989_ axi_controller.state\[0\] _1998_ _1996_ _1995_ VGND VGND VPWR VPWR _1999_
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3010_ _1304_ _1309_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__and3_1
XFILLER_64_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4961_ net411 _0590_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_1
X_3912_ axi_controller.read_addr_reg\[13\] net6 net196 VGND VGND VPWR VPWR _0279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4892_ net378 _0045_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3843_ _1926_ _1928_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3774_ _1876_ _1878_ axi_controller.reg_input_data\[24\] VGND VGND VPWR VPWR _1879_
+ sky130_fd_sc_hd__or3b_1
X_2725_ cordic_inst.cordic_inst.y\[14\] _0923_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__a21bo_1
X_2656_ _0984_ _0986_ _0989_ _0990_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__and4_1
X_2587_ _0771_ _0772_ _0778_ cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR _0922_
+ sky130_fd_sc_hd__o31ai_2
XFILLER_86_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4326_ net120 net192 net155 axi_controller.result_out\[17\] VGND VGND VPWR VPWR _0577_
+ sky130_fd_sc_hd__a22o_1
X_4257_ _2211_ _2212_ net199 VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__o21ai_1
Xfanout159 net162 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout148 _1790_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_2
X_3208_ cordic_inst.cordic_inst.y\[25\] cordic_inst.cordic_inst.sin_out\[25\] net207
+ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux2_1
X_4188_ net225 _2155_ cordic_inst.cordic_inst.cos_out\[19\] VGND VGND VPWR VPWR _2156_
+ sky130_fd_sc_hd__a21oi_1
X_3139_ _1332_ _1361_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__nand2_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2510_ net272 _0787_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__nand2_1
X_3490_ net183 _1712_ _1713_ _1714_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__a31o_1
XFILLER_5_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2441_ net282 _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nor2_1
X_2372_ net304 net313 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nand2b_2
X_4111_ net261 _2086_ cordic_inst.cordic_inst.sin_out\[10\] VGND VGND VPWR VPWR _2088_
+ sky130_fd_sc_hd__a21oi_1
X_4042_ axi_controller.result_out\[0\] _2028_ net205 VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
XFILLER_83_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4944_ net394 _0573_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4875_ net388 axi_controller.reg_input_data\[7\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3826_ net282 _0614_ _1917_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.next_state\[0\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3757_ cordic_inst.deg_handler_inst.theta_norm\[30\] _1863_ VGND VGND VPWR VPWR _0031_
+ sky130_fd_sc_hd__xor2_1
X_2708_ _0852_ _1030_ _0850_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_30_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3688_ cordic_inst.deg_handler_inst.theta_norm\[4\] _1820_ VGND VGND VPWR VPWR _0034_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2639_ _0844_ _0869_ _0968_ _0970_ _0867_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__o41a_1
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4309_ net194 _1990_ _2254_ _2255_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__o31ai_1
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2990_ cordic_inst.cordic_inst.x\[9\] _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__and2b_1
X_4660_ net406 _0390_ _0092_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[4\] sky130_fd_sc_hd__dfrtp_1
X_3611_ _1777_ _1778_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__or2_1
X_4591_ net360 _0323_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[24\] sky130_fd_sc_hd__dfxtp_1
X_3542_ net176 _1599_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__or2_1
X_3473_ net183 _1699_ _1700_ _1701_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a31o_1
XFILLER_69_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2424_ net239 _0698_ _0637_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__a21bo_1
X_2355_ net292 _0654_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__or2_1
XFILLER_69_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2286_ net107 VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__inv_2
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4025_ axi_controller.reg_input_data\[0\] _2018_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__or2_1
XFILLER_25_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4927_ net373 _0027_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_4858_ net384 _0067_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[22\] sky130_fd_sc_hd__dfxtp_1
X_3809_ _1905_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__inv_2
X_4789_ net397 _0516_ _0211_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_87_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2973_ _1263_ _1275_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__nand2_1
X_4712_ net403 _0439_ _0134_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[5\] sky130_fd_sc_hd__dfrtp_1
X_4643_ net394 _0374_ net329 VGND VGND VPWR VPWR axi_controller.result_out\[20\] sky130_fd_sc_hd__dfrtp_1
X_4574_ net370 _0306_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_3525_ _1556_ _1609_ _1739_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3456_ cordic_inst.cordic_inst.angle\[25\] net171 net163 cordic_inst.cordic_inst.z\[25\]
+ _1688_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__a221o_1
X_3387_ _1554_ _1610_ _1618_ _1622_ _1547_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__o2111ai_4
X_2407_ _0740_ _0741_ net281 _0664_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_4_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2338_ cordic_inst.cordic_inst.x\[10\] cordic_inst.cordic_inst.x\[11\] cordic_inst.cordic_inst.x\[12\]
+ cordic_inst.cordic_inst.x\[13\] net310 net300 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux4_1
X_2269_ net282 VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__inv_2
X_4008_ net87 _2009_ _2010_ net352 VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o211a_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3310_ net275 _1481_ _1548_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__mux2_1
X_4290_ net78 _2243_ _2244_ net353 VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__o211a_1
X_3241_ _1478_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__nand2_1
X_3172_ _1293_ _1440_ _1323_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2956_ cordic_inst.cordic_inst.x\[4\] _1256_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__nor2_1
X_2887_ net263 _1080_ _1174_ _1171_ net241 net244 VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__mux4_2
X_4626_ net412 _0357_ net347 VGND VGND VPWR VPWR axi_controller.result_out\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4557_ net359 _0289_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[23\] sky130_fd_sc_hd__dfxtp_1
X_3508_ _1727_ net183 _1627_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__and3b_1
X_4488_ net345 VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__inv_2
X_3439_ cordic_inst.cordic_inst.angle\[29\] net170 net159 cordic_inst.cordic_inst.z\[29\]
+ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__a22o_1
XFILLER_66_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3790_ _1874_ _1890_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__nor2_1
X_2810_ _1078_ _1112_ net231 VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__mux2_1
X_2741_ _0955_ _0957_ _1037_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nand3_1
X_2672_ _0812_ _0999_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__nand2_1
X_4411_ net340 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__inv_2
X_4342_ net123 net193 net154 axi_controller.result_out\[1\] VGND VGND VPWR VPWR _0593_
+ sky130_fd_sc_hd__a22o_1
X_4273_ axi_controller.result_out\[30\] net199 VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__nor2_1
Xfanout308 net311 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_4
Xfanout319 net320 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__buf_4
XFILLER_86_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3224_ cordic_inst.cordic_inst.y\[9\] cordic_inst.cordic_inst.sin_out\[9\] net213
+ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
.ends

