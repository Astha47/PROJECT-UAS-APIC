// DRAM Controller for LPDDR4 - Fixed version
module dram_controller #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 32,
    parameter AXI4_ID_WIDTH = 4,
    parameter LPDDR4_CAPACITY_GB = 4
)(
    // Clock and Reset
    input wire                     clk,
    input wire                     rst_n,
    
    // AXI4 Interface (slave interface to the interconnect)
    // Write Address Channel
    input  wire [AXI4_ID_WIDTH-1:0] S_AXI4_AWID,
    input  wire [ADDR_WIDTH-1:0]    S_AXI4_AWADDR,
    input  wire [7:0]               S_AXI4_AWLEN,
    input  wire [2:0]               S_AXI4_AWSIZE,
    input  wire [1:0]               S_AXI4_AWBURST,
    input  wire                     S_AXI4_AWVALID,
    output wire                     S_AXI4_AWREADY,
    
    // Write Data Channel
    input  wire [DATA_WIDTH-1:0]    S_AXI4_WDATA,
    input  wire [(DATA_WIDTH/8)-1:0] S_AXI4_WSTRB,
    input  wire                     S_AXI4_WLAST,
    input  wire                     S_AXI4_WVALID,
    output wire                     S_AXI4_WREADY,
    
    // Write Response Channel
    output wire [AXI4_ID_WIDTH-1:0] S_AXI4_BID,
    output wire [1:0]               S_AXI4_BRESP,
    output wire                     S_AXI4_BVALID,
    input  wire                     S_AXI4_BREADY,
    
    // Read Address Channel
    input  wire [AXI4_ID_WIDTH-1:0] S_AXI4_ARID,
    input  wire [ADDR_WIDTH-1:0]    S_AXI4_ARADDR,
    input  wire [7:0]               S_AXI4_ARLEN,
    input  wire [2:0]               S_AXI4_ARSIZE,
    input  wire [1:0]               S_AXI4_ARBURST,
    input  wire                     S_AXI4_ARVALID,
    output wire                     S_AXI4_ARREADY,
    
    // Read Data Channel
    output wire [AXI4_ID_WIDTH-1:0] S_AXI4_RID,
    output wire [DATA_WIDTH-1:0]    S_AXI4_RDATA,
    output wire [1:0]               S_AXI4_RRESP,
    output wire                     S_AXI4_RLAST,
    output wire                     S_AXI4_RVALID,
    input  wire                     S_AXI4_RREADY,
    
    // LPDDR4 Interface
    output wire                    lpddr4_ck_t,         // Clock (true)
    output wire                    lpddr4_ck_c,         // Clock (complement)
    output wire                    lpddr4_cke,          // Clock enable
    output wire                    lpddr4_reset_n,      // Reset
    output wire                    lpddr4_cs_n,         // Chip select
    output wire [5:0]              lpddr4_ca,           // Command/Address bus
    inout  wire [31:0]             lpddr4_dq,           // Data bus (32-bit for dual channel)
    inout  wire [3:0]              lpddr4_dqs_t,        // Data strobe (true)
    inout  wire [3:0]              lpddr4_dqs_c         // Data strobe (complement)
);

    // Internal parameters
    localparam ROW_BITS = 16;        // 16 bits for 4GB LPDDR4
    localparam COL_BITS = 10;        // 10 bits for column addressing
    localparam BANK_BITS = 3;        // 8 banks per bank group
    localparam BANKGROUP_BITS = 2;   // 4 bank groups
    
    // State machine for memory controller
    localparam IDLE = 4'd0,
               INIT = 4'd1,
               WRITE_ACT = 4'd2,
               WRITE_CAS = 4'd3,
               WRITE_DATA = 4'd4,
               WRITE_RESP = 4'd5,
               READ_ACT = 4'd6,
               READ_CAS = 4'd7,
               READ_DATA = 4'd8,
               PRECHARGE = 4'd9,
               REFRESH = 4'd10;
    
    reg [3:0] state, next_state;
    
    // Command encoding for LPDDR4
    localparam CMD_MRW     = 6'b000001, // Mode Register Write
               CMD_MRR     = 6'b000010, // Mode Register Read
               CMD_REFRESH = 6'b000100, // Refresh
               CMD_PRECHARGE = 6'b001000, // Precharge
               CMD_ACTIVATE = 6'b010000, // Activate
               CMD_WRITE   = 6'b100000, // Write
               CMD_READ    = 6'b100001, // Read
               CMD_NOP     = 6'b000000; // No Operation
    
    // AXI transaction tracking
    reg [AXI4_ID_WIDTH-1:0] active_id;
    reg [7:0]  active_len;
    reg [2:0]  active_size;
    reg [1:0]  active_burst;
    reg [ADDR_WIDTH-1:0] active_addr;
    
    // Address decomposition
    reg [ROW_BITS-1:0] row_addr;
    reg [COL_BITS-1:0] col_addr;
    reg [BANK_BITS-1:0] bank_addr;
    reg [BANKGROUP_BITS-1:0] bank_group;
    
    reg [7:0]  burst_counter;
    reg [15:0] refresh_counter;
    
    // LPDDR4 control signals
    reg        lpddr4_ck_reg;
    reg        lpddr4_cke_reg;
    reg        lpddr4_cs_n_reg;
    reg [5:0]  lpddr4_ca_reg;
    
    // Data path
    reg [31:0] lpddr4_dq_out;
    reg        lpddr4_dq_oe;  // Output enable for DQ bus
    reg [3:0]  lpddr4_dqs_out;
    reg        lpddr4_dqs_oe; // Output enable for DQS
    
    // Data buffers
    reg [DATA_WIDTH-1:0] read_data_buffer [0:15];  // Support up to 16 beats
    reg [DATA_WIDTH-1:0] write_data_buffer [0:15]; // Support up to 16 beats
    reg [(DATA_WIDTH/8)-1:0] write_strb_buffer [0:15];
    
    // Initialization sequence tracking
    reg [7:0]  init_state;
    reg [15:0] init_timer;
    reg        init_done;

    reg [3:0] state_counter; // For tracking state transitions during initialization
    
    // Timing parameters (in clock cycles)
    localparam tRCD = 6;  // ACT to CAS delay
    localparam tRP = 6;   // Precharge time
    localparam tRAS = 16; // ACT to PRE delay
    localparam tRC = 22;  // ACT to ACT delay
    localparam tRFC = 35; // Refresh cycle time
    localparam tREFI = 1950; // Refresh interval (avg)
    
    reg [7:0] timing_counter;
    
    // Assign physical interface signals
    assign lpddr4_ck_t = lpddr4_ck_reg;
    assign lpddr4_ck_c = ~lpddr4_ck_reg;
    assign lpddr4_cke = lpddr4_cke_reg;
    assign lpddr4_reset_n = rst_n;
    assign lpddr4_cs_n = lpddr4_cs_n_reg;
    assign lpddr4_ca = lpddr4_ca_reg;
    
    // Bidirectional data interface
    assign lpddr4_dq = lpddr4_dq_oe ? lpddr4_dq_out : 32'bz;
    assign lpddr4_dqs_t = lpddr4_dqs_oe ? lpddr4_dqs_out : 4'bz;
    assign lpddr4_dqs_c = lpddr4_dqs_oe ? ~lpddr4_dqs_out : 4'bz;
    
    // AXI interface assignments
    assign S_AXI4_AWREADY = (state == IDLE) && !refresh_counter[15] && init_done;
    assign S_AXI4_WREADY = (state == WRITE_DATA);

    // BUG
    assign S_AXI4_ARREADY =  (state == IDLE) && !refresh_counter[15] && init_done;
    
    assign S_AXI4_BID = active_id;
    assign S_AXI4_BRESP = 2'b00; // OKAY
    assign S_AXI4_BVALID = (state == WRITE_RESP);
    
    // Fixed AXI4 read data assignments
    assign S_AXI4_RID = active_id;
    assign S_AXI4_RDATA = read_data_buffer[burst_counter];
    assign S_AXI4_RRESP = 2'b00; // OKAY
    assign S_AXI4_RLAST = (state == READ_DATA) && (burst_counter == active_len);
    assign S_AXI4_RVALID = (state == READ_DATA) && (burst_counter <= active_len);
    
    // Address translation from AXI to LPDDR4
    always @(*) begin
        // Map the AXI address to LPDDR4 address components
        // This is a simple mapping example - adjust according to your memory layout
        row_addr = active_addr[ROW_BITS+COL_BITS+BANK_BITS+BANKGROUP_BITS-1:COL_BITS+BANK_BITS+BANKGROUP_BITS];
        col_addr = active_addr[COL_BITS+BANK_BITS+BANKGROUP_BITS-1:BANK_BITS+BANKGROUP_BITS];
        bank_addr = active_addr[BANK_BITS+BANKGROUP_BITS-1:BANKGROUP_BITS];
        bank_group = active_addr[BANKGROUP_BITS-1:0];
    end
    
    // Clock generation (simplified - in real design would be PLL/DLL controlled)
    always @(posedge clk) begin
        lpddr4_ck_reg <= ~lpddr4_ck_reg;
    end
    
    // Main state machine
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= INIT;
            state_counter <= 4'd0;
            init_state <= 8'd0;
            init_timer <= 16'd0;
            init_done <= 1'b0;
            lpddr4_cke_reg <= 1'b0;
            lpddr4_cs_n_reg <= 1'b1;
            lpddr4_ca_reg <= 6'b0;
            refresh_counter <= 16'd0;
            lpddr4_dq_oe <= 1'b0;
            lpddr4_dqs_oe <= 1'b0;
            burst_counter <= 8'd0;
            timing_counter <= 8'd0;
        end else begin
            state <= next_state;
            state_counter <= next_state;
            
            // Refresh counter
            if (refresh_counter < tREFI)
                refresh_counter <= refresh_counter + 1'b1;
                
            // Timing counter for command delays
            if (timing_counter > 0)
                timing_counter <= timing_counter - 1'b1;
            
            case (state)
                INIT: begin
                    if (!init_done) begin
                        $display("Time %t: DRAM_CTRL INIT: init_state=%d, init_timer=%d", $time, init_state, init_timer);
                        case (init_state)
                            8'd0: begin // Power-up wait
                                if (init_timer < 16'd200) begin
                                    init_timer <= init_timer + 1'b1;
                                    lpddr4_cke_reg <= 1'b0;
                                    lpddr4_cs_n_reg <= 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd1: begin // CKE high
                                lpddr4_cke_reg <= 1'b1;
                                lpddr4_cs_n_reg <= 1'b1;
                                if (init_timer < 16'd10) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd2: begin // Reset command
                                lpddr4_cs_n_reg <= 1'b0;
                                lpddr4_ca_reg <= CMD_MRW;
                                if (init_timer < 16'd5) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd3: begin // Mode Register 1 - Device Feature
                                lpddr4_cs_n_reg <= 1'b0;
                                lpddr4_ca_reg <= CMD_MRW;
                                if (init_timer < 16'd5) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd4: begin // Mode Register 2 - Device Feature 2
                                lpddr4_cs_n_reg <= 1'b0;
                                lpddr4_ca_reg <= CMD_MRW;
                                if (init_timer < 16'd5) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd5: begin // Mode Register 3 - I/O Configuration
                                lpddr4_cs_n_reg <= 1'b0;
                                lpddr4_ca_reg <= CMD_MRW;
                                if (init_timer < 16'd5) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd6: begin // ZQ Calibration Start
                                lpddr4_cs_n_reg <= 1'b0;
                                lpddr4_ca_reg <= CMD_MRW;
                                if (init_timer < 16'd10) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd7: begin // Wait for ZQ calibration completion
                                lpddr4_cs_n_reg <= 1'b1; // NOP
                                if (init_timer < 16'd50) begin // tZQINIT wait
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd8: begin // Additional mode register setup
                                lpddr4_cs_n_reg <= 1'b0;
                                lpddr4_ca_reg <= CMD_MRW;
                                if (init_timer < 16'd5) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd9: begin // Precharge all banks
                                lpddr4_cs_n_reg <= 1'b0;
                                lpddr4_ca_reg <= CMD_PRECHARGE;
                                if (init_timer < 16'd10) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_timer <= 16'd0;
                                    init_state <= init_state + 1'b1;
                                end
                            end
                            
                            8'd10: begin // Final initialization step
                                lpddr4_cs_n_reg <= 1'b1;
                                if (init_timer < 16'd50) begin
                                    init_timer <= init_timer + 1'b1;
                                end else begin
                                    init_done <= 1'b1;
                                end
                            end
                            
                            default: begin
                                // Skip to completion for any undefined states
                                init_state <= 8'd10;
                                init_timer <= 16'd0;
                            end
                        endcase
                    end
                end
                
                IDLE: begin
                    lpddr4_cs_n_reg <= 1'b1; // Default to NOP
                    lpddr4_dq_oe <= 1'b0;
                    lpddr4_dqs_oe <= 1'b0;
                    burst_counter <= 8'd0;
                    
                    if (refresh_counter >= tREFI) begin
                        refresh_counter <= 16'd0;
                    end else if (S_AXI4_AWVALID) begin
                        active_id <= S_AXI4_AWID;
                        active_addr <= S_AXI4_AWADDR;
                        active_len <= S_AXI4_AWLEN;
                        active_size <= S_AXI4_AWSIZE;
                        active_burst <= S_AXI4_AWBURST;
                    end else if (S_AXI4_ARVALID) begin
                        active_id <= S_AXI4_ARID;
                        active_addr <= S_AXI4_ARADDR;
                        active_len <= S_AXI4_ARLEN;
                        active_size <= S_AXI4_ARSIZE;
                        active_burst <= S_AXI4_ARBURST;
                    end
                end
                
                WRITE_ACT: begin
                    lpddr4_cs_n_reg <= 1'b0;
                    lpddr4_ca_reg <= CMD_ACTIVATE;
                    // In real implementation, row address would be sent here
                    timing_counter <= tRCD; // Set timing for ACT-to-CAS
                end
                
                WRITE_CAS: begin
                    if (timing_counter == 0) begin
                        lpddr4_cs_n_reg <= 1'b0;
                        lpddr4_ca_reg <= CMD_WRITE;
                        // Column address and bank information would be sent
                    end else begin
                        lpddr4_cs_n_reg <= 1'b1; // NOP while waiting
                    end
                end
                
                WRITE_DATA: begin
                    if (S_AXI4_WVALID) begin
                        // Store data for current beat
                        write_data_buffer[burst_counter] <= S_AXI4_WDATA;
                        write_strb_buffer[burst_counter] <= S_AXI4_WSTRB;
                        
                        // Prepare data for LPDDR4
                        lpddr4_dq_oe <= 1'b1;
                        lpddr4_dqs_oe <= 1'b1;
                        lpddr4_dq_out <= S_AXI4_WDATA;
                        lpddr4_dqs_out <= 4'b1010; // Toggle DQS for data valid
                        
                        if (S_AXI4_WLAST || burst_counter == active_len) begin
                            // Last beat
                        end else begin
                            burst_counter <= burst_counter + 1'b1;
                        end
                    end
                end
                
                WRITE_RESP: begin
                    lpddr4_cs_n_reg <= 1'b1; // NOP
                    lpddr4_dq_oe <= 1'b0;
                    lpddr4_dqs_oe <= 1'b0;
                end
                
                READ_ACT: begin
                    lpddr4_cs_n_reg <= 1'b0;
                    lpddr4_ca_reg <= CMD_ACTIVATE;
                    // Row address would be sent
                    timing_counter <= tRCD; // Set timing for ACT-to-CAS
                end
                
                READ_CAS: begin
                    if (timing_counter == 0) begin
                        lpddr4_cs_n_reg <= 1'b0;
                        lpddr4_ca_reg <= CMD_READ;
                        $display("Time %t: DRAM_CTRL READ_CAS: Issuing READ command. active_addr=0x%h, active_len=%d", $time, active_addr, active_len);
                        // Column address would be sent
                        timing_counter <= 8; // CAS latency for read data
                    end else begin
                        lpddr4_cs_n_reg <= 1'b1; // NOP while waiting
                    end
                end
                
                READ_DATA: begin
                    // Fixed read data logic for proper AXI4 compliance
                    if (timing_counter == 0) begin
                        // Simulate read data being available after CAS latency
                        read_data_buffer[burst_counter] <= lpddr4_dq;
                        $display("Time %t: DRAM_CTRL READ_DATA: burst_cnt=%d, active_len=%d, S_AXI4_RREADY=%b, S_AXI4_RVALID_OUT=%b, lpddr4_dq=0x%h",
                                 $time, burst_counter, active_len, S_AXI4_RREADY, S_AXI4_RVALID, lpddr4_dq);
                        
                        // Increment burst counter when data is accepted by master
                        if (S_AXI4_RVALID && S_AXI4_RREADY && burst_counter <= active_len) begin
                            $display("Time %t: DRAM_CTRL READ_DATA: Handshake OK. burst_counter %d -> %d.", $time, burst_counter, burst_counter + 1);
                            burst_counter <= burst_counter + 1'b1;
                        end else if (burst_counter < active_len) begin
                            timing_counter <= 2; // Small delay between beats
                        end
                    end else if (timing_counter > 0) begin
                        timing_counter <= timing_counter - 1'b1;
                    end
                end
                
                PRECHARGE: begin
                    lpddr4_cs_n_reg <= 1'b0;
                    lpddr4_ca_reg <= CMD_PRECHARGE;
                    timing_counter <= tRP;
                end
                
                REFRESH: begin
                    lpddr4_cs_n_reg <= 1'b0;
                    lpddr4_ca_reg <= CMD_REFRESH;
                    timing_counter <= tRFC;
                end
            endcase
        end
    end
    
    // Next state logic
    always @(*) begin
        next_state = state;
        
        case (state)
            INIT: begin
                if (init_done) next_state = IDLE;
            end
            
            IDLE: begin
                if (refresh_counter >= tREFI) begin
                    next_state = REFRESH;
                end else if (S_AXI4_AWVALID && init_done) begin
                    next_state = WRITE_ACT;
                end else if (S_AXI4_ARVALID && init_done) begin
                    next_state = READ_ACT;
                end
            end
            
            WRITE_ACT: begin
                if (timing_counter == 0) next_state = WRITE_CAS;
            end
            
            WRITE_CAS: begin
                next_state = WRITE_DATA;
            end
            
            WRITE_DATA: begin
                if (S_AXI4_WLAST && S_AXI4_WVALID) next_state = WRITE_RESP;
            end
            
            WRITE_RESP: begin
                if (S_AXI4_BREADY) next_state = PRECHARGE;
            end
            
            READ_ACT: begin
                if (timing_counter == 0) next_state = READ_CAS;
            end
            
            READ_CAS: begin
                if (timing_counter == 0) begin
                    $display("Time %t: DRAM_CTRL READ_CAS: Next State -> READ_DATA. CAS latency met.", $time);
                    next_state = READ_DATA;
                end
            end
            
            READ_DATA: begin
                // If burst_counter has incremented past active_len, all data has been sent and acknowledged by master
                if (burst_counter > active_len) begin
                    $display("Time %t: DRAM_CTRL READ_DATA: Next State -> PRECHARGE. Read complete. burst_cnt=%d, active_len=%d", $time, burst_counter, active_len);
                    next_state = PRECHARGE;
                end
            end
            
            PRECHARGE: begin
                if (timing_counter == 0) next_state = IDLE;
            end
            
            REFRESH: begin
                if (timing_counter == 0) next_state = IDLE;
            end
        endcase
    end

endmodule
