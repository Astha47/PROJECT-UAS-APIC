* NGSPICE file created from cordic_system.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

.subckt cordic_system VGND VPWR aclk araddr[0] araddr[10] araddr[11] araddr[12] araddr[13]
+ araddr[14] araddr[15] araddr[16] araddr[17] araddr[18] araddr[19] araddr[1] araddr[20]
+ araddr[21] araddr[22] araddr[23] araddr[24] araddr[25] araddr[26] araddr[27] araddr[28]
+ araddr[29] araddr[2] araddr[30] araddr[31] araddr[3] araddr[4] araddr[5] araddr[6]
+ araddr[7] araddr[8] araddr[9] aresetn arready arvalid awaddr[0] awaddr[10] awaddr[11]
+ awaddr[12] awaddr[13] awaddr[14] awaddr[15] awaddr[16] awaddr[17] awaddr[18] awaddr[19]
+ awaddr[1] awaddr[20] awaddr[21] awaddr[22] awaddr[23] awaddr[24] awaddr[25] awaddr[26]
+ awaddr[27] awaddr[28] awaddr[29] awaddr[2] awaddr[30] awaddr[31] awaddr[3] awaddr[4]
+ awaddr[5] awaddr[6] awaddr[7] awaddr[8] awaddr[9] awready awvalid bready bresp[0]
+ bresp[1] bvalid rdata[0] rdata[10] rdata[11] rdata[12] rdata[13] rdata[14] rdata[15]
+ rdata[16] rdata[17] rdata[18] rdata[19] rdata[1] rdata[20] rdata[21] rdata[22] rdata[23]
+ rdata[24] rdata[25] rdata[26] rdata[27] rdata[28] rdata[29] rdata[2] rdata[30] rdata[31]
+ rdata[3] rdata[4] rdata[5] rdata[6] rdata[7] rdata[8] rdata[9] rready rresp[0] rresp[1]
+ rvalid wdata[0] wdata[10] wdata[11] wdata[12] wdata[13] wdata[14] wdata[15] wdata[16]
+ wdata[17] wdata[18] wdata[19] wdata[1] wdata[20] wdata[21] wdata[22] wdata[23] wdata[24]
+ wdata[25] wdata[26] wdata[27] wdata[28] wdata[29] wdata[2] wdata[30] wdata[31] wdata[3]
+ wdata[4] wdata[5] wdata[6] wdata[7] wdata[8] wdata[9] wready wstrb[0] wstrb[1] wstrb[2]
+ wstrb[3] wvalid
X_3155_ _1318_ _1441_ _1329_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__o21a_1
XFILLER_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3086_ _1387_ _1388_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__and2_1
XFILLER_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3988_ _1939_ _1941_ _1997_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__or3_1
X_2939_ _1103_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__xnor2_1
X_4609_ net357 _0341_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4960_ net399 _0589_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4891_ net358 _0044_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_3911_ axi_controller.read_addr_reg\[12\] net5 net198 VGND VGND VPWR VPWR _0278_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3842_ net145 net70 net194 VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__a21oi_1
X_3773_ axi_controller.reg_input_data\[30\] axi_controller.reg_input_data\[29\] _1877_
+ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__nand3_1
X_2724_ _0925_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__or2_1
X_2655_ cordic_inst.cordic_inst.y\[25\] _0988_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nand2_1
X_2586_ net250 _0770_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__nor2_1
X_4325_ net121 net192 net156 axi_controller.result_out\[18\] VGND VGND VPWR VPWR _0576_
+ sky130_fd_sc_hd__a22o_1
X_4256_ net313 _2214_ _2215_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__and3_1
Xfanout149 _1790_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4187_ cordic_inst.cordic_inst.cos_out\[18\] _2147_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__or2_1
X_3207_ cordic_inst.cordic_inst.y\[26\] cordic_inst.cordic_inst.sin_out\[26\] net209
+ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
X_3138_ net183 _1421_ _1429_ net165 cordic_inst.cordic_inst.x\[20\] VGND VGND VPWR
+ VPWR _0518_ sky130_fd_sc_hd__a32o_1
XFILLER_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3069_ cordic_inst.cordic_inst.x\[23\] _1334_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2440_ _0719_ _0722_ _0727_ _0720_ net285 net235 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__mux4_1
X_2371_ net241 net302 VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__nand2_1
X_4110_ cordic_inst.cordic_inst.sin_out\[10\] net258 _2086_ VGND VGND VPWR VPWR _2087_
+ sky130_fd_sc_hd__and3_1
X_4041_ cordic_inst.cordic_inst.cos_out\[0\] cordic_inst.cordic_inst.sin_out\[0\]
+ net316 VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__mux2_2
X_4943_ net394 _0572_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
X_4874_ net365 axi_controller.reg_input_data\[6\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3825_ cordic_inst.cordic_inst.start cordic_inst.cordic_inst.state\[1\] cordic_inst.cordic_inst.state\[0\]
+ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__o21ba_1
XFILLER_20_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3756_ cordic_inst.deg_handler_inst.theta_norm\[29\] cordic_inst.deg_handler_inst.theta_norm\[28\]
+ _1859_ net254 VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__o31a_1
X_2707_ _0854_ _0858_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__or3_1
X_3687_ net252 _1819_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__nand2_1
X_2638_ _0869_ _0968_ _0970_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__or3_1
X_2569_ _0889_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nor2_1
X_4308_ axi_controller.state\[0\] axi_controller.state\[1\] _0621_ net144 VGND VGND
+ VPWR VPWR _2255_ sky130_fd_sc_hd__or4b_1
X_4239_ cordic_inst.cordic_inst.sin_out\[25\] net257 _2199_ net231 VGND VGND VPWR
+ VPWR _2201_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_2_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3610_ cordic_inst.deg_handler_inst.theta_abs\[24\] cordic_inst.deg_handler_inst.theta_abs\[25\]
+ cordic_inst.deg_handler_inst.theta_abs\[26\] cordic_inst.deg_handler_inst.theta_abs\[27\]
+ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__or4_1
X_4590_ net382 _0322_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[23\] sky130_fd_sc_hd__dfxtp_1
X_3541_ net182 _1601_ _1749_ _1750_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a31o_1
X_3472_ cordic_inst.cordic_inst.angle\[21\] net173 net162 cordic_inst.cordic_inst.z\[21\]
+ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__a22o_1
X_2423_ _0684_ _0693_ _0750_ _0756_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__and4_1
X_2354_ net284 _0685_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__a21o_1
X_2285_ net349 VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__inv_2
X_4024_ net103 _1963_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__nand2_2
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4926_ net372 _0026_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4857_ net378 _0066_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[21\] sky130_fd_sc_hd__dfxtp_1
X_3808_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1900_
+ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__and3_1
X_4788_ net404 _0515_ _0210_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[17\] sky130_fd_sc_hd__dfrtp_2
X_3739_ cordic_inst.deg_handler_inst.theta_norm\[23\] cordic_inst.deg_handler_inst.theta_norm\[22\]
+ _1849_ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_7_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2972_ cordic_inst.cordic_inst.x\[3\] _1262_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__or2_1
X_4711_ net379 _0438_ _0133_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[4\] sky130_fd_sc_hd__dfrtp_1
X_4642_ net403 _0373_ net340 VGND VGND VPWR VPWR axi_controller.result_out\[19\] sky130_fd_sc_hd__dfrtp_1
X_4573_ net364 _0305_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3524_ net175 _1610_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__or2_1
X_3455_ _1686_ _1687_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__nor2_1
X_2406_ _0679_ net218 _0739_ net284 VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__a22o_1
XFILLER_39_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3386_ _1540_ _1546_ _1621_ _1624_ _1539_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__o311a_1
X_2337_ net278 _0670_ _0671_ _0631_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o31a_1
X_2268_ cordic_inst.cordic_inst.cos_out\[26\] VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__inv_2
X_4007_ axi_controller.reg_input_data\[24\] _2008_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__or2_1
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4909_ net360 _0039_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3240_ net248 cordic_inst.cordic_inst.z\[24\] VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__or2_1
X_3171_ net178 _1452_ _1453_ cordic_inst.cordic_inst.next_state\[1\] cordic_inst.cordic_inst.x\[11\]
+ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__o32a_1
XFILLER_19_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2955_ _1257_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__inv_2
X_2886_ _1180_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__or2_1
XFILLER_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4625_ net398 _0356_ net339 VGND VGND VPWR VPWR axi_controller.result_out\[2\] sky130_fd_sc_hd__dfrtp_1
X_4556_ net355 _0288_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[22\] sky130_fd_sc_hd__dfxtp_1
X_3507_ _1535_ _1625_ _1626_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__and3_1
X_4487_ net329 VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__inv_2
X_3438_ _1475_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__xnor2_1
X_3369_ _1568_ _1606_ _1563_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__o21ba_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2740_ cordic_inst.cordic_inst.y\[10\] net166 _1052_ _1053_ VGND VGND VPWR VPWR _0540_
+ sky130_fd_sc_hd__a22o_1
X_2671_ _1004_ _1005_ net263 net164 VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4410_ net328 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__inv_2
X_4341_ net134 net191 net155 axi_controller.result_out\[2\] VGND VGND VPWR VPWR _0592_
+ sky130_fd_sc_hd__a22o_1
Xfanout309 net312 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_2
X_4272_ axi_controller.result_out\[29\] _2229_ net200 VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__mux2_1
X_3223_ cordic_inst.cordic_inst.y\[10\] cordic_inst.cordic_inst.sin_out\[10\] net211
+ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3154_ _1293_ _1323_ _1440_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__or3_1
X_3085_ cordic_inst.cordic_inst.x\[26\] _1386_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__or2_1
XFILLER_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3987_ net61 net62 net63 VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__or3b_1
XFILLER_11_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2938_ _1116_ _1131_ _1178_ net251 VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__a31o_1
X_2869_ net219 _1139_ _1143_ net221 VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__a22o_1
X_4608_ net351 _0340_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[26\] sky130_fd_sc_hd__dfxtp_1
X_4539_ net362 _0271_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4890_ net358 _0043_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_3910_ axi_controller.read_addr_reg\[11\] net4 net195 VGND VGND VPWR VPWR _0277_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3841_ axi_controller.state\[1\] net349 VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__nand2_1
X_3772_ axi_controller.reg_input_data\[28\] axi_controller.reg_input_data\[27\] axi_controller.reg_input_data\[26\]
+ axi_controller.reg_input_data\[25\] VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__and4_1
XFILLER_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2723_ _0965_ _1041_ _0933_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__a21o_1
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2654_ cordic_inst.cordic_inst.y\[25\] _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__or2_1
X_2585_ cordic_inst.cordic_inst.y\[15\] _0917_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__xnor2_1
X_4324_ net122 net192 _2256_ axi_controller.result_out\[19\] VGND VGND VPWR VPWR _0575_
+ sky130_fd_sc_hd__a22o_1
X_4255_ cordic_inst.cordic_inst.sin_out\[27\] net256 _2213_ VGND VGND VPWR VPWR _2215_
+ sky130_fd_sc_hd__nand3_1
X_4186_ net230 _2152_ _2153_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__or3_1
X_3206_ cordic_inst.cordic_inst.y\[27\] cordic_inst.cordic_inst.sin_out\[27\] net209
+ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
X_3137_ _1343_ _1375_ _1420_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__nand3_1
XFILLER_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3068_ cordic_inst.cordic_inst.x\[23\] _1334_ _1337_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2370_ net288 net294 VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nor2_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4040_ net100 _2019_ _2027_ net350 VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o211a_1
XFILLER_37_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4942_ net393 _0571_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4873_ net365 axi_controller.reg_input_data\[5\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3824_ _1874_ _1915_ _1916_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a21bo_1
X_3755_ cordic_inst.deg_handler_inst.theta_norm\[29\] _1862_ VGND VGND VPWR VPWR _0029_
+ sky130_fd_sc_hd__xnor2_1
X_3686_ cordic_inst.deg_handler_inst.theta_norm\[0\] cordic_inst.deg_handler_inst.theta_norm\[1\]
+ cordic_inst.deg_handler_inst.theta_norm\[3\] cordic_inst.deg_handler_inst.theta_norm\[2\]
+ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__or4_1
X_2706_ _0860_ _0861_ _0972_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__inv_2
X_2568_ cordic_inst.cordic_inst.y\[3\] _0888_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nor2_1
X_4307_ _1989_ _2253_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__nor2_1
X_2499_ _0793_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__xnor2_1
X_4238_ net257 _2199_ cordic_inst.cordic_inst.sin_out\[25\] VGND VGND VPWR VPWR _2200_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4169_ _2137_ _2138_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__or2_1
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ cordic_inst.cordic_inst.angle\[2\] net172 net160 cordic_inst.cordic_inst.z\[2\]
+ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__a22o_1
X_3471_ _1488_ _1691_ _1486_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__a21o_1
X_2422_ _0750_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and2_1
X_2353_ _0673_ net219 _0687_ net221 net277 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a221o_1
X_2284_ cordic_inst.state\[1\] VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__inv_2
X_4023_ net103 _1963_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__and2_1
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4925_ net372 _0025_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_4856_ net378 _0065_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[20\] sky130_fd_sc_hd__dfxtp_1
X_3807_ axi_controller.reg_input_data\[26\] _1904_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4787_ net404 _0514_ _0209_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[16\] sky130_fd_sc_hd__dfrtp_4
X_3738_ cordic_inst.deg_handler_inst.theta_norm\[23\] _1851_ VGND VGND VPWR VPWR _0023_
+ sky130_fd_sc_hd__xnor2_1
X_3669_ _0617_ _1783_ _1808_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_7_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2971_ _1269_ _1272_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__a21o_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4710_ net379 _0437_ _0132_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[3\] sky130_fd_sc_hd__dfrtp_1
X_4641_ net403 _0372_ net340 VGND VGND VPWR VPWR axi_controller.result_out\[18\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_12_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4572_ net369 _0304_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3523_ cordic_inst.cordic_inst.angle\[8\] net171 net160 cordic_inst.cordic_inst.z\[8\]
+ _1738_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__a221o_1
X_3454_ _1478_ _1658_ _1659_ net176 VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__a31o_1
X_2405_ net216 _0729_ _0731_ _0713_ net275 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__a221o_1
X_3385_ _1538_ _1544_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__nand2_1
X_2336_ net240 _0650_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nor2_1
X_2267_ net270 VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__inv_2
X_4006_ net106 _1963_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__nand2_2
XFILLER_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4908_ net366 _0038_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_4839_ net367 _0078_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3170_ _1318_ _1321_ _1441_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__and3b_1
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2954_ cordic_inst.cordic_inst.x\[4\] _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__and2_1
X_2885_ _1098_ _1185_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__or3_1
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4624_ net399 _0355_ net336 VGND VGND VPWR VPWR axi_controller.result_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_4555_ net355 _0287_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[21\] sky130_fd_sc_hd__dfxtp_1
X_3506_ net179 _1724_ _1725_ _1726_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a31o_1
X_4486_ net322 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__inv_2
X_3437_ net249 cordic_inst.cordic_inst.z\[28\] _1667_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__a21oi_1
X_3368_ _1568_ _1606_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__nor2_1
X_2319_ cordic_inst.cordic_inst.x\[22\] cordic_inst.cordic_inst.x\[23\] cordic_inst.cordic_inst.x\[24\]
+ cordic_inst.cordic_inst.x\[25\] net307 net301 VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux4_1
X_3299_ cordic_inst.cordic_inst.z\[11\] _1537_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__or2_1
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2670_ _0810_ _1000_ _1003_ net176 VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a31o_1
XFILLER_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4340_ net137 net191 net155 axi_controller.result_out\[3\] VGND VGND VPWR VPWR _0591_
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4271_ net313 _2224_ _2225_ _2228_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__a31o_1
X_3222_ cordic_inst.cordic_inst.y\[11\] cordic_inst.cordic_inst.sin_out\[11\] net210
+ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
X_3153_ _1287_ _1290_ _1294_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__and3_1
X_3084_ cordic_inst.cordic_inst.x\[26\] _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__nand2_1
XFILLER_23_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3986_ net107 net103 _1922_ _1943_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__nand4_1
X_2937_ _1236_ _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__and2_1
X_4607_ net352 _0339_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[25\] sky130_fd_sc_hd__dfxtp_2
X_2868_ _1132_ _1140_ net234 VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2799_ net283 _1099_ _1101_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__a21oi_1
X_4538_ net362 _0270_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_4469_ net338 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__inv_2
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3840_ net68 net35 axi_controller.state\[0\] net349 VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__and4b_1
X_3771_ axi_controller.reg_input_data\[22\] _1875_ axi_controller.reg_input_data\[23\]
+ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2722_ _0963_ _1039_ _0930_ _0939_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__o211ai_2
X_2653_ _0802_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__xnor2_1
X_2584_ cordic_inst.cordic_inst.y\[15\] _0917_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__nor2_1
X_4323_ net124 net193 _2256_ axi_controller.result_out\[20\] VGND VGND VPWR VPWR _0574_
+ sky130_fd_sc_hd__a22o_1
X_4254_ net256 _2213_ cordic_inst.cordic_inst.sin_out\[27\] VGND VGND VPWR VPWR _2214_
+ sky130_fd_sc_hd__a21o_1
X_4185_ net261 _2151_ cordic_inst.cordic_inst.sin_out\[19\] VGND VGND VPWR VPWR _2153_
+ sky130_fd_sc_hd__a21oi_1
X_3205_ cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.sin_out\[28\] net207
+ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
X_3136_ _1427_ _1428_ cordic_inst.cordic_inst.x\[21\] net165 VGND VGND VPWR VPWR _0519_
+ sky130_fd_sc_hd__a2bb2o_1
X_3067_ _1335_ _1339_ _1346_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__or4_1
XFILLER_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3969_ axi_controller.write_addr_reg\[18\] net45 net190 VGND VGND VPWR VPWR _0317_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_0_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4941_ net392 _0570_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_1
XFILLER_18_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4872_ net365 axi_controller.reg_input_data\[4\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3823_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1872_
+ _1903_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__or4_1
XFILLER_33_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3754_ cordic_inst.deg_handler_inst.theta_norm\[28\] _1859_ net254 VGND VGND VPWR
+ VPWR _1862_ sky130_fd_sc_hd__o21ai_1
X_3685_ cordic_inst.deg_handler_inst.theta_norm\[3\] _1818_ VGND VGND VPWR VPWR _0033_
+ sky130_fd_sc_hd__xor2_1
X_2705_ net183 _1021_ _1028_ net167 cordic_inst.cordic_inst.y\[20\] VGND VGND VPWR
+ VPWR _0550_ sky130_fd_sc_hd__a32o_1
X_2636_ _0968_ _0970_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_42_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2567_ _0899_ _0900_ _0892_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a21o_1
X_4306_ _1976_ _2252_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__nand2_1
X_2498_ net271 _0789_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__nand2_1
X_4237_ cordic_inst.cordic_inst.sin_out\[24\] _2191_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4168_ cordic_inst.cordic_inst.sin_out\[17\] net260 _2136_ net229 VGND VGND VPWR
+ VPWR _2138_ sky130_fd_sc_hd__a31o_1
X_4099_ _2076_ _2077_ net203 _2074_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__o211a_1
X_3119_ net181 _1413_ _1416_ net163 cordic_inst.cordic_inst.x\[26\] VGND VGND VPWR
+ VPWR _0524_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_41_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3470_ _1486_ _1488_ _1691_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__nand3_1
X_2421_ net244 _0755_ _0753_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__o21ai_2
X_2352_ cordic_inst.cordic_inst.x\[6\] cordic_inst.cordic_inst.x\[7\] cordic_inst.cordic_inst.x\[8\]
+ cordic_inst.cordic_inst.x\[9\] net309 net297 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__mux4_1
X_2283_ axi_controller.state\[1\] VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__inv_2
X_4022_ net95 _2009_ _2017_ net346 VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o211a_1
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4924_ net374 _0024_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_4855_ net374 _0063_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3806_ _1903_ _1899_ axi_controller.reg_input_data\[25\] VGND VGND VPWR VPWR _1904_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4786_ net401 _0513_ _0208_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3737_ cordic_inst.deg_handler_inst.theta_norm\[22\] _1849_ net254 VGND VGND VPWR
+ VPWR _1851_ sky130_fd_sc_hd__o21ai_1
X_3668_ cordic_inst.deg_handler_inst.theta_abs\[21\] net152 net149 _1813_ VGND VGND
+ VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
X_3599_ cordic_inst.deg_handler_inst.theta_abs\[10\] _1766_ VGND VGND VPWR VPWR _1767_
+ sky130_fd_sc_hd__or2_1
X_2619_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout290 net292 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2970_ cordic_inst.cordic_inst.x\[2\] _1265_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4640_ net407 _0371_ net343 VGND VGND VPWR VPWR axi_controller.result_out\[17\] sky130_fd_sc_hd__dfrtp_1
X_4571_ net369 _0303_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3522_ _1611_ _1618_ _1737_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__o21a_1
X_3453_ _1478_ _1658_ _1659_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__a21oi_1
X_2404_ _0668_ _0681_ net236 VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__mux2_1
X_3384_ _1616_ _1619_ _1620_ _1550_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__o31a_1
X_2335_ net285 _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__nor2_1
X_2266_ cordic_inst.cordic_inst.x\[0\] VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__inv_2
XFILLER_38_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4005_ net106 _1963_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__and2_1
XFILLER_38_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4907_ net366 _0037_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_4838_ net379 _0075_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4769_ net384 _0496_ _0191_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_45_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2953_ _1177_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2884_ net262 _1161_ _1162_ _1158_ net243 net240 VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__mux4_1
X_4623_ net381 _0354_ net317 VGND VGND VPWR VPWR axi_controller.result_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_4554_ net355 _0286_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[20\] sky130_fd_sc_hd__dfxtp_1
X_3505_ cordic_inst.cordic_inst.angle\[13\] net172 net159 cordic_inst.cordic_inst.z\[13\]
+ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__a22o_1
X_4485_ net321 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__inv_2
X_3436_ cordic_inst.cordic_inst.z\[30\] net158 _1673_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__o21a_1
X_3367_ _1575_ _1605_ _1570_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__a21boi_1
X_2318_ cordic_inst.cordic_inst.x\[18\] cordic_inst.cordic_inst.x\[19\] cordic_inst.cordic_inst.x\[20\]
+ cordic_inst.cordic_inst.x\[21\] net311 net300 VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux4_1
X_3298_ net266 _1504_ _1536_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__mux2_1
XFILLER_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput100 wdata[7] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ net313 _2226_ _2227_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__nor3b_1
X_3221_ cordic_inst.cordic_inst.y\[12\] cordic_inst.cordic_inst.sin_out\[12\] net210
+ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
X_3152_ _1287_ _1290_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__nand2_1
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3083_ _1213_ _1223_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3985_ _0624_ _1994_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__nor2_1
X_2936_ cordic_inst.cordic_inst.x\[28\] _1235_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__or2_1
X_2867_ _1148_ _1157_ _1164_ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__or4b_1
X_4606_ net352 _0338_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[24\] sky130_fd_sc_hd__dfxtp_1
X_2798_ net218 _1095_ _1100_ net221 net277 VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__a221o_1
X_4537_ net362 _0269_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_4468_ net335 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__inv_2
X_3419_ _1655_ _1657_ _1480_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__a21o_1
X_4399_ net317 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_46_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3770_ axi_controller.reg_input_data\[19\] axi_controller.reg_input_data\[18\] axi_controller.reg_input_data\[21\]
+ axi_controller.reg_input_data\[20\] VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__a211o_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2721_ _0963_ _1039_ _0939_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__o21a_1
X_2652_ net170 _0796_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__nor2_1
X_2583_ cordic_inst.cordic_inst.y\[15\] _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nand2_1
X_4322_ net125 net193 _2256_ axi_controller.result_out\[21\] VGND VGND VPWR VPWR _0573_
+ sky130_fd_sc_hd__a22o_1
X_4253_ cordic_inst.cordic_inst.sin_out\[26\] cordic_inst.cordic_inst.sin_out\[25\]
+ _2199_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__or3_1
X_3204_ cordic_inst.cordic_inst.y\[29\] cordic_inst.cordic_inst.sin_out\[29\] net207
+ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux2_1
X_4184_ cordic_inst.cordic_inst.sin_out\[19\] net261 _2151_ VGND VGND VPWR VPWR _2152_
+ sky130_fd_sc_hd__and3_1
X_3135_ _1341_ _1348_ _1421_ net177 VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__a31o_1
X_3066_ _1341_ _1347_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__and2_1
X_3968_ axi_controller.write_addr_reg\[17\] net44 net190 VGND VGND VPWR VPWR _0316_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2919_ net269 _1211_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__a21o_1
X_3899_ axi_controller.read_addr_reg\[0\] net2 net197 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
XFILLER_2_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4940_ net393 _0569_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4871_ net368 axi_controller.reg_input_data\[3\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3822_ _1880_ _1914_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3753_ cordic_inst.deg_handler_inst.theta_norm\[28\] _1859_ VGND VGND VPWR VPWR _1861_
+ sky130_fd_sc_hd__nor2_1
X_3684_ cordic_inst.deg_handler_inst.theta_norm\[0\] cordic_inst.deg_handler_inst.theta_norm\[1\]
+ cordic_inst.deg_handler_inst.theta_norm\[2\] net252 VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__o31a_1
X_2704_ _0837_ _0864_ _0973_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__nand3_1
X_2635_ _0860_ _0969_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__nand2_1
X_2566_ _0899_ _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4305_ axi_controller.read_addr_reg\[5\] _1977_ axi_controller.read_addr_reg\[3\]
+ axi_controller.read_addr_reg\[4\] VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__and4b_1
X_2497_ _0825_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nand2_1
X_4236_ net223 _2196_ cordic_inst.cordic_inst.cos_out\[25\] VGND VGND VPWR VPWR _2198_
+ sky130_fd_sc_hd__a21oi_1
X_4167_ net260 _2136_ cordic_inst.cordic_inst.sin_out\[17\] VGND VGND VPWR VPWR _2137_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3118_ _1390_ _1412_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__nand2_1
X_4098_ cordic_inst.cordic_inst.sin_out\[8\] net258 _2075_ net228 VGND VGND VPWR VPWR
+ _2077_ sky130_fd_sc_hd__a31o_1
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3049_ _1203_ _1351_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2420_ net265 _0722_ _0723_ _0720_ net240 net235 VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__mux4_2
X_2351_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__inv_2
X_2282_ cordic_inst.state\[0\] VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__inv_2
X_4021_ axi_controller.reg_input_data\[31\] _2008_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__or2_1
XFILLER_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4923_ net373 _0023_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4854_ net374 _0062_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[18\] sky130_fd_sc_hd__dfxtp_1
X_3805_ _1901_ _1903_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__xnor2_1
X_4785_ net397 _0512_ _0207_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[14\] sky130_fd_sc_hd__dfrtp_4
X_3736_ cordic_inst.deg_handler_inst.theta_norm\[22\] _1850_ VGND VGND VPWR VPWR _0022_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3667_ _1783_ _1808_ _1812_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__o21ai_1
X_3598_ cordic_inst.deg_handler_inst.theta_abs\[9\] _1765_ VGND VGND VPWR VPWR _1766_
+ sky130_fd_sc_hd__or2_1
X_2618_ cordic_inst.cordic_inst.y\[9\] _0951_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__nor2_1
X_2549_ _0599_ _0882_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4219_ cordic_inst.cordic_inst.sin_out\[23\] net257 _2180_ _2182_ VGND VGND VPWR
+ VPWR _2183_ sky130_fd_sc_hd__a31o_1
XFILLER_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout291 net293 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_4
Xfanout280 net282 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__buf_2
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ net370 _0302_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3521_ net176 _1619_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__nor2_1
XFILLER_7_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3452_ net180 _1680_ _1684_ _1685_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a31o_1
X_2403_ net243 _0659_ _0736_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__o22a_1
X_3383_ _1551_ _1620_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__nor2_1
X_2334_ _0660_ _0668_ net236 VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux2_1
X_2265_ cordic_inst.cordic_inst.x\[5\] VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__inv_2
X_4004_ net146 _1943_ _2002_ _2007_ net350 VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o221a_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4906_ net367 _0036_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4837_ net379 _0064_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4768_ net384 _0495_ _0190_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_3719_ net253 _1839_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__nand2_1
X_4699_ net393 _0426_ _0121_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2952_ net270 _1170_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2883_ net241 _1162_ _1070_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__a21bo_1
X_4622_ net363 _0353_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[7\] sky130_fd_sc_hd__dfxtp_1
X_4553_ net364 _0285_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[19\] sky130_fd_sc_hd__dfxtp_1
X_3504_ _1514_ _1627_ _1533_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__a21o_1
X_4484_ net324 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__inv_2
X_3435_ cordic_inst.cordic_inst.angle\[30\] net176 _1670_ _1672_ net162 VGND VGND
+ VPWR VPWR _1673_ sky130_fd_sc_hd__a221o_1
X_3366_ _1591_ _1602_ _1604_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__o21ai_1
X_3297_ net294 net302 _0706_ net288 _0713_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__a221o_1
X_2317_ net278 _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__nor2_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 wdata[8] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3220_ cordic_inst.cordic_inst.y\[13\] cordic_inst.cordic_inst.sin_out\[13\] net213
+ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__mux2_1
X_3151_ net184 _1430_ _1438_ net167 cordic_inst.cordic_inst.x\[16\] VGND VGND VPWR
+ VPWR _0514_ sky130_fd_sc_hd__a32o_1
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3082_ cordic_inst.cordic_inst.x\[27\] _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_33_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3984_ _1993_ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__inv_2
XFILLER_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ cordic_inst.cordic_inst.x\[29\] _1233_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nand2_1
X_2866_ _1165_ _1166_ _1168_ net275 VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__a2bb2o_1
X_4605_ net371 _0337_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2797_ cordic_inst.cordic_inst.y\[7\] cordic_inst.cordic_inst.y\[8\] cordic_inst.cordic_inst.y\[9\]
+ cordic_inst.cordic_inst.y\[10\] net308 net297 VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__mux4_1
X_4536_ net351 _0268_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_4467_ net337 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__inv_2
X_3418_ net248 cordic_inst.cordic_inst.z\[23\] _1491_ _1656_ VGND VGND VPWR VPWR _1657_
+ sky130_fd_sc_hd__a211oi_1
X_4398_ net320 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__inv_2
X_3349_ net267 _1587_ _1585_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2720_ _0947_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__nor2_1
X_2651_ cordic_inst.cordic_inst.y\[26\] _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__xor2_1
X_2582_ _0672_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__xnor2_2
X_4321_ net126 net193 net157 axi_controller.result_out\[22\] VGND VGND VPWR VPWR _0572_
+ sky130_fd_sc_hd__a22o_1
X_4252_ cordic_inst.cordic_inst.cos_out\[27\] _2210_ net313 VGND VGND VPWR VPWR _2212_
+ sky130_fd_sc_hd__a21o_1
X_3203_ cordic_inst.cordic_inst.y\[30\] cordic_inst.cordic_inst.sin_out\[30\] net209
+ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__mux2_1
X_4183_ cordic_inst.cordic_inst.sin_out\[18\] _2143_ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__or2_1
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3134_ _1341_ _1421_ _1348_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__a21oi_1
X_3065_ _1349_ _1359_ _1362_ _1367_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__nor4_1
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3967_ axi_controller.write_addr_reg\[16\] net43 net190 VGND VGND VPWR VPWR _0315_
+ sky130_fd_sc_hd__mux2_1
X_2918_ net270 _1090_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__a21o_1
X_3898_ net77 _1965_ _1973_ net347 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__o211a_1
X_2849_ _1117_ _1122_ net235 VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__mux2_1
X_4519_ net380 _0006_ _0085_ VGND VGND VPWR VPWR cordic_inst.state\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_46_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4870_ net368 axi_controller.reg_input_data\[2\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3821_ _1878_ _1898_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__nor2_1
X_3752_ cordic_inst.deg_handler_inst.theta_norm\[28\] _1860_ VGND VGND VPWR VPWR _0028_
+ sky130_fd_sc_hd__xnor2_1
X_3683_ cordic_inst.deg_handler_inst.theta_norm\[2\] _1817_ VGND VGND VPWR VPWR _0030_
+ sky130_fd_sc_hd__xnor2_1
X_2703_ cordic_inst.cordic_inst.y\[21\] net165 _1027_ net183 VGND VGND VPWR VPWR _0551_
+ sky130_fd_sc_hd__a22o_1
X_2634_ cordic_inst.cordic_inst.y\[16\] _0859_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__or2_1
X_2565_ cordic_inst.cordic_inst.y\[2\] _0891_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__xor2_1
X_4304_ net86 _2243_ _2251_ net346 VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o211a_1
X_2496_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__inv_2
X_4235_ cordic_inst.cordic_inst.cos_out\[25\] net223 _2196_ VGND VGND VPWR VPWR _2197_
+ sky130_fd_sc_hd__and3_1
X_4166_ cordic_inst.cordic_inst.sin_out\[16\] _2128_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3117_ cordic_inst.cordic_inst.x\[27\] net163 _1415_ net176 VGND VGND VPWR VPWR _0525_
+ sky130_fd_sc_hd__o2bb2ai_1
X_4097_ net258 _2075_ cordic_inst.cordic_inst.sin_out\[8\] VGND VGND VPWR VPWR _2076_
+ sky130_fd_sc_hd__a21oi_1
X_3048_ _1195_ _1198_ _1202_ _1204_ net273 VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__o41a_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2350_ _0653_ _0674_ net235 VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux2_1
X_2281_ cordic_inst.deg_handler_inst.theta_abs\[22\] VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__inv_2
XFILLER_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4020_ net94 _2009_ _2016_ net347 VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o211a_1
XFILLER_38_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4922_ net373 _0022_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_4853_ net374 _0061_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3804_ _1874_ _1902_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__or2_1
X_4784_ net401 _0511_ _0206_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[13\] sky130_fd_sc_hd__dfrtp_4
X_3735_ net254 _1849_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__nand2_1
X_3666_ _0616_ _1808_ cordic_inst.deg_handler_inst.theta_abs\[21\] VGND VGND VPWR
+ VPWR _1812_ sky130_fd_sc_hd__o21bai_1
X_2617_ cordic_inst.cordic_inst.y\[9\] _0951_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__nand2_1
X_3597_ cordic_inst.deg_handler_inst.theta_abs\[8\] _1764_ VGND VGND VPWR VPWR _1765_
+ sky130_fd_sc_hd__or2_1
X_2548_ _0599_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4218_ net316 _2181_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__nand2_1
X_2479_ _0806_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4149_ net227 _2120_ cordic_inst.cordic_inst.cos_out\[15\] VGND VGND VPWR VPWR _2121_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout270 net273 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_4
Xfanout292 net293 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_2
Xfanout281 net282 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_1
XFILLER_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3520_ net182 _1734_ _1735_ _1736_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__a31o_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3451_ cordic_inst.cordic_inst.angle\[26\] net173 net161 cordic_inst.cordic_inst.z\[26\]
+ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__a22o_1
X_2402_ net284 _0675_ net218 _0687_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__a22o_1
X_3382_ _1550_ _1616_ _1620_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__a21oi_1
X_2333_ cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.x\[16\] cordic_inst.cordic_inst.x\[17\]
+ cordic_inst.cordic_inst.x\[18\] net311 net299 VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__mux4_1
X_2264_ net264 VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__inv_2
X_4003_ net68 _0622_ _0624_ _1923_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__a22o_1
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4905_ net366 _0035_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_4836_ net379 _0053_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4767_ net385 _0494_ _0189_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_3718_ cordic_inst.deg_handler_inst.theta_norm\[15\] _1837_ VGND VGND VPWR VPWR _1839_
+ sky130_fd_sc_hd__or2_1
X_4698_ net392 _0425_ _0120_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3649_ cordic_inst.deg_handler_inst.theta_abs\[13\] _1769_ VGND VGND VPWR VPWR _1803_
+ sky130_fd_sc_hd__nand2_1
XFILLER_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2951_ _1253_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2882_ _1182_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or2_1
X_4621_ net363 _0352_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_4552_ net355 _0284_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[18\] sky130_fd_sc_hd__dfxtp_1
X_3503_ _1514_ _1533_ _1627_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__nand3_1
X_4483_ net317 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__inv_2
X_3434_ _1474_ _1669_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__or2_1
X_3365_ _1575_ _1603_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__and2_1
X_3296_ _1514_ _1534_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__nand2_1
X_2316_ net239 _0650_ _0637_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__a21boi_1
XFILLER_26_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4819_ net403 _0546_ _0241_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput102 wdata[9] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3150_ _1332_ _1361_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__or2_1
X_3081_ _1224_ _1383_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3983_ axi_controller.write_addr_reg\[3\] axi_controller.write_addr_reg\[4\] _1953_
+ axi_controller.write_addr_reg\[5\] VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__or4b_1
XFILLER_16_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2934_ cordic_inst.cordic_inst.x\[29\] _1233_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__and2_1
X_2865_ net285 _1094_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4604_ net370 _0336_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
X_2796_ _1093_ _1096_ net235 VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux2_1
X_4535_ net362 _0267_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_4466_ net337 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__inv_2
X_3417_ _1495_ _1497_ _1654_ _1496_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__o22ai_1
X_4397_ net319 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
X_3348_ _1564_ _1586_ _1577_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__a21o_1
X_3279_ cordic_inst.cordic_inst.z\[14\] _1517_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__and2_1
XFILLER_38_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2650_ _0797_ _0803_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__xor2_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2581_ _0770_ _0780_ net251 VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a21oi_1
X_4320_ net127 net193 net157 axi_controller.result_out\[23\] VGND VGND VPWR VPWR _0571_
+ sky130_fd_sc_hd__a22o_1
X_4251_ cordic_inst.cordic_inst.cos_out\[27\] _2210_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__nor2_1
X_3202_ net263 cordic_inst.cordic_inst.sin_out\[31\] net207 VGND VGND VPWR VPWR _0497_
+ sky130_fd_sc_hd__mux2_1
X_4182_ _2146_ _2150_ axi_controller.result_out\[18\] net204 VGND VGND VPWR VPWR _0372_
+ sky130_fd_sc_hd__o2bb2a_1
X_3133_ net183 _1423_ _1426_ net165 cordic_inst.cordic_inst.x\[22\] VGND VGND VPWR
+ VPWR _0520_ sky130_fd_sc_hd__a32o_1
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3064_ _1365_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_19_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3966_ axi_controller.write_addr_reg\[15\] net42 net188 VGND VGND VPWR VPWR _0314_
+ sky130_fd_sc_hd__mux2_1
X_2917_ net270 _1210_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__a21o_1
X_3897_ axi_controller.reg_input_data\[15\] _1964_ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__or2_1
XFILLER_31_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2848_ _1149_ _1150_ net283 VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__mux2_1
X_2779_ net242 _1081_ net215 VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__a21o_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4518_ net318 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__inv_2
X_4449_ net325 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__inv_2
XFILLER_37_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ axi_controller.reg_input_data\[30\] _1913_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__xor2_1
X_3751_ net254 _1859_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__nand2_1
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2702_ _0843_ _1022_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__xnor2_1
X_3682_ cordic_inst.deg_handler_inst.theta_norm\[0\] cordic_inst.deg_handler_inst.theta_norm\[1\]
+ net252 VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__o21ai_1
X_2633_ _0961_ _0966_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__and3_1
X_2564_ _0896_ _0897_ _0895_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__o21ai_1
X_4303_ axi_controller.reg_input_data\[23\] _2242_ VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__or2_1
X_2495_ cordic_inst.cordic_inst.y\[23\] _0827_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__xnor2_1
X_4234_ cordic_inst.cordic_inst.cos_out\[24\] _2188_ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__or2_1
X_4165_ axi_controller.result_out\[16\] _2135_ net204 VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
X_3116_ _1385_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_2_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4096_ cordic_inst.cordic_inst.sin_out\[7\] _2065_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__or2_1
X_3047_ net273 _1202_ _1217_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3949_ _0619_ _1991_ axi_controller.reg_done_flag VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__o21a_1
XFILLER_3_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2280_ cordic_inst.deg_handler_inst.theta_abs\[20\] VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4921_ net373 _0021_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_4852_ net374 _0060_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[16\] sky130_fd_sc_hd__dfxtp_1
X_3803_ axi_controller.reg_input_data\[23\] _1890_ axi_controller.reg_input_data\[24\]
+ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__o21a_1
XFILLER_21_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4783_ net400 _0510_ _0205_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3734_ cordic_inst.deg_handler_inst.theta_norm\[21\] _1847_ VGND VGND VPWR VPWR _1849_
+ sky130_fd_sc_hd__or2_1
X_3665_ cordic_inst.deg_handler_inst.theta_abs\[20\] net152 net149 _1811_ VGND VGND
+ VPWR VPWR _0065_ sky130_fd_sc_hd__a22o_1
X_2616_ _0762_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__xnor2_1
X_3596_ cordic_inst.deg_handler_inst.theta_abs\[7\] _1763_ VGND VGND VPWR VPWR _1764_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_7_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2547_ _0756_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__xnor2_1
X_2478_ net170 _0807_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__nor2_1
X_4217_ net257 _2180_ cordic_inst.cordic_inst.sin_out\[23\] VGND VGND VPWR VPWR _2181_
+ sky130_fd_sc_hd__a21o_1
XFILLER_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4148_ cordic_inst.cordic_inst.cos_out\[14\] cordic_inst.cordic_inst.cos_out\[13\]
+ _2111_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__or3_1
X_4079_ cordic_inst.cordic_inst.sin_out\[5\] cordic_inst.cordic_inst.sin_out\[4\]
+ _2045_ net259 VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_26_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout282 net287 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_2
Xfanout271 net273 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__buf_2
Xfanout260 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_2
XFILLER_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout293 cordic_inst.cordic_inst.i\[2\] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3450_ _1661_ _1663_ _1679_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__or3_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2401_ _0703_ net216 _0710_ _0713_ net275 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__a221o_1
X_3381_ cordic_inst.cordic_inst.z\[9\] _1549_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__and2_1
X_2332_ net245 _0659_ net170 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__a21o_1
X_2263_ cordic_inst.cordic_inst.y\[0\] VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__inv_2
X_4002_ _1921_ _2006_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nor2_1
XFILLER_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4904_ net366 _0034_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4835_ net383 _0008_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.isNegative
+ sky130_fd_sc_hd__dfxtp_2
X_4766_ net385 _0493_ _0188_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_3717_ cordic_inst.deg_handler_inst.theta_norm\[15\] _1838_ VGND VGND VPWR VPWR _0014_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4697_ net392 _0424_ _0119_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_3648_ _1769_ net147 _1802_ net151 cordic_inst.deg_handler_inst.theta_abs\[12\] VGND
+ VGND VPWR VPWR _0056_ sky130_fd_sc_hd__a32o_1
X_3579_ cordic_inst.cordic_inst.x\[0\] cordic_inst.cordic_inst.cos_out\[0\] net208
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2950_ _0602_ _1251_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__nor2_1
XFILLER_15_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2881_ net262 _1134_ _1136_ _1141_ net242 net239 VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__mux4_2
X_4620_ net363 _0351_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4551_ net362 _0283_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3502_ cordic_inst.cordic_inst.angle\[14\] net172 net159 cordic_inst.cordic_inst.z\[14\]
+ _1723_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a221o_1
X_4482_ net324 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__inv_2
X_3433_ net268 net158 _1671_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o21a_1
X_3364_ cordic_inst.cordic_inst.z\[4\] _1574_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__or2_1
X_3295_ cordic_inst.cordic_inst.z\[12\] _1513_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__or2_1
X_2315_ _0646_ _0649_ net291 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux2_1
XFILLER_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4818_ net406 _0545_ _0240_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_5_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ net400 _0476_ _0171_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput103 wstrb[0] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_1
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3080_ net215 _1214_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__or2_1
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3982_ axi_controller.write_addr_reg\[31\] net60 net189 VGND VGND VPWR VPWR _0330_
+ sky130_fd_sc_hd__mux2_1
X_2933_ cordic_inst.cordic_inst.x\[28\] _1235_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2864_ net233 _1087_ _1071_ net238 VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a211o_1
XFILLER_31_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2795_ cordic_inst.cordic_inst.y\[31\] _1091_ _1094_ _1097_ net240 net243 VGND VGND
+ VPWR VPWR _1098_ sky130_fd_sc_hd__mux4_1
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4603_ net382 _0335_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
X_4534_ net362 _0266_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_4465_ net337 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__inv_2
X_3416_ _1532_ _1628_ _1649_ _1496_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__a211o_1
X_4396_ net319 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_2
X_3347_ net241 net302 net288 VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__o21a_1
X_3278_ net267 _1481_ _1516_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__mux2_1
XFILLER_39_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2580_ _0873_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nor2_1
X_4250_ cordic_inst.deg_handler_inst.kuadran\[0\] _2204_ VGND VGND VPWR VPWR _2210_
+ sky130_fd_sc_hd__nor2_1
X_3201_ cordic_inst.cordic_inst.state\[1\] cordic_inst.cordic_inst.state\[0\] VGND
+ VGND VPWR VPWR _1472_ sky130_fd_sc_hd__nand2_1
X_4181_ _2148_ _2149_ net204 VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__o21a_1
X_3132_ _1339_ _1422_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__nand2_1
X_3063_ cordic_inst.cordic_inst.x\[17\] _1364_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__and2_1
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3965_ axi_controller.write_addr_reg\[14\] net41 net188 VGND VGND VPWR VPWR _0313_
+ sky130_fd_sc_hd__mux2_1
X_3896_ net76 _1965_ _1972_ net347 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__o211a_1
X_2916_ net270 _1209_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__a21o_1
X_2847_ net262 _1085_ _1086_ _1083_ net233 net232 VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__mux4_2
XFILLER_12_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2778_ net241 _1080_ _1070_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__a21bo_1
X_4517_ net325 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__inv_2
X_4448_ net326 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__inv_2
X_4379_ net332 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
XFILLER_37_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_36_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3750_ cordic_inst.deg_handler_inst.theta_norm\[27\] _1857_ VGND VGND VPWR VPWR _1859_
+ sky130_fd_sc_hd__or2_1
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2701_ cordic_inst.cordic_inst.y\[22\] net165 _1026_ net183 VGND VGND VPWR VPWR _0552_
+ sky130_fd_sc_hd__a22o_1
X_3681_ cordic_inst.deg_handler_inst.theta_norm\[1\] _1816_ VGND VGND VPWR VPWR _0019_
+ sky130_fd_sc_hd__xnor2_1
X_2632_ _0926_ _0933_ _0965_ _0964_ _0936_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__o32a_1
X_2563_ _0896_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__or2_1
X_4302_ net85 _2243_ _2250_ net348 VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o211a_1
X_4233_ net201 _2195_ _2187_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21oi_1
X_2494_ cordic_inst.cordic_inst.y\[23\] _0827_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__nor2_1
X_4164_ _2133_ _2134_ _2131_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__o21ai_1
X_4095_ cordic_inst.cordic_inst.cos_out\[8\] _2072_ _2073_ VGND VGND VPWR VPWR _2074_
+ sky130_fd_sc_hd__a21o_1
X_3115_ _1387_ _1413_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3046_ _1335_ _1339_ _1343_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__or4_1
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3948_ net70 _1990_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__nand2_1
X_3879_ net107 axi_controller.state\[3\] _1961_ _1942_ axi_controller.state\[0\] VGND
+ VGND VPWR VPWR _1962_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_29_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4920_ net373 _0020_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4851_ net360 _0059_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[15\] sky130_fd_sc_hd__dfxtp_1
X_3802_ axi_controller.reg_input_data\[25\] _1899_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__xnor2_1
X_4782_ net400 _0509_ _0204_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[11\] sky130_fd_sc_hd__dfrtp_2
X_3733_ cordic_inst.deg_handler_inst.theta_norm\[21\] _1848_ VGND VGND VPWR VPWR _0021_
+ sky130_fd_sc_hd__xnor2_1
X_3664_ _0616_ _1808_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__xnor2_1
X_2615_ net271 _0760_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a21oi_1
X_3595_ cordic_inst.deg_handler_inst.theta_abs\[6\] _1762_ VGND VGND VPWR VPWR _1763_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_7_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2546_ _0743_ _0750_ net250 VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__a21o_1
X_2477_ _0810_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nand2_1
X_4216_ cordic_inst.cordic_inst.sin_out\[22\] _2176_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__or2_1
X_4147_ axi_controller.result_out\[14\] _2119_ net204 VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux2_1
X_4078_ cordic_inst.cordic_inst.cos_out\[6\] _2058_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__xor2_1
X_3029_ _1328_ _1331_ _1325_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__nand3b_2
XTAP_TAPCELL_ROW_26_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout250 net251 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_2
Xfanout261 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_4
Xfanout272 net273 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__buf_2
Xfanout283 net287 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_2
XFILLER_19_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout294 net296 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__buf_2
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2400_ net243 _0725_ _0734_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__o21a_1
X_3380_ _1611_ _1618_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__and2_1
X_2331_ net170 _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nor2_1
X_2262_ cordic_inst.cordic_inst.y\[5\] VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__inv_2
X_4001_ net111 _0610_ axi_controller.state\[2\] VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__a21oi_1
X_4903_ net371 _0033_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4834_ net386 _0561_ _0256_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[31\] sky130_fd_sc_hd__dfrtp_1
X_4765_ net384 _0492_ _0187_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_3716_ net253 _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4696_ net394 _0423_ _0118_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3647_ cordic_inst.deg_handler_inst.theta_abs\[12\] _1768_ VGND VGND VPWR VPWR _1802_
+ sky130_fd_sc_hd__nand2_1
X_3578_ cordic_inst.cordic_inst.x\[1\] cordic_inst.cordic_inst.cos_out\[1\] net208
+ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2529_ _0850_ _0854_ _0862_ _0863_ _0848_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__o32a_1
XFILLER_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ net239 _1136_ _1070_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a21bo_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4550_ net362 _0282_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3501_ _1520_ _1717_ _1722_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__a21boi_1
X_4481_ net324 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__inv_2
X_3432_ _0614_ cordic_inst.cordic_inst.angle\[31\] _1473_ _1670_ net162 VGND VGND
+ VPWR VPWR _1671_ sky130_fd_sc_hd__a221o_1
X_3363_ _1594_ _1601_ _1592_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__a21oi_1
X_3294_ _1506_ _1530_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__or2_1
X_2314_ cordic_inst.cordic_inst.x\[27\] cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.x\[29\]
+ cordic_inst.cordic_inst.x\[30\] net305 net296 VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux4_1
XFILLER_26_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4817_ net406 _0544_ _0239_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[14\] sky130_fd_sc_hd__dfrtp_4
X_4748_ net400 _0475_ _0170_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4679_ net396 _0406_ _0101_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput104 wstrb[1] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_1
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3981_ axi_controller.write_addr_reg\[30\] net59 net189 VGND VGND VPWR VPWR _0329_
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2932_ _1082_ _1225_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_33_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2863_ net283 _1097_ _1100_ net218 VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a22o_1
X_4602_ net370 _0334_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
X_2794_ _1095_ _1096_ net290 VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__mux2_1
X_4533_ net357 _0265_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4464_ net335 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__inv_2
X_3415_ _1637_ _1653_ _1652_ _1642_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__o2bb2a_1
X_4395_ net319 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
X_3346_ _1583_ _1584_ net248 VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__a21oi_1
X_3277_ net220 _0712_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__nand2_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3200_ _0603_ _1471_ _1470_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
X_4180_ cordic_inst.cordic_inst.cos_out\[18\] net226 _2147_ net315 VGND VGND VPWR
+ VPWR _2149_ sky130_fd_sc_hd__a31o_1
X_3131_ _1424_ _1425_ cordic_inst.cordic_inst.x\[23\] net169 VGND VGND VPWR VPWR _0521_
+ sky130_fd_sc_hd__a2bb2o_1
X_3062_ cordic_inst.cordic_inst.x\[17\] _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__nor2_1
XFILLER_36_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3964_ axi_controller.write_addr_reg\[13\] net40 net187 VGND VGND VPWR VPWR _0312_
+ sky130_fd_sc_hd__mux2_1
X_3895_ axi_controller.reg_input_data\[14\] _1964_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__or2_1
X_2915_ _1195_ _1198_ _1205_ net270 VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__o31a_1
X_2846_ _1118_ _1125_ net290 VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__mux2_1
X_2777_ net237 _1079_ _1071_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__a21o_1
X_4516_ net328 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__inv_2
X_4447_ net326 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__inv_2
X_4378_ net340 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
X_3329_ cordic_inst.cordic_inst.z\[5\] _1567_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__and2_1
XFILLER_27_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ _0825_ _1023_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__xor2_1
X_3680_ cordic_inst.deg_handler_inst.theta_norm\[0\] net255 VGND VGND VPWR VPWR _1816_
+ sky130_fd_sc_hd__nand2_1
X_2631_ _0918_ _0924_ _0919_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a21o_1
X_2562_ cordic_inst.cordic_inst.y\[1\] _0894_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__xnor2_1
X_4301_ axi_controller.reg_input_data\[22\] _2242_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__or2_1
X_4232_ _2189_ _2190_ _2194_ net231 VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__o22a_1
X_2493_ cordic_inst.cordic_inst.y\[23\] _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__nand2_1
X_4163_ cordic_inst.cordic_inst.cos_out\[16\] net226 _2132_ net315 VGND VGND VPWR
+ VPWR _2134_ sky130_fd_sc_hd__a31o_1
X_4094_ cordic_inst.cordic_inst.cos_out\[8\] _2072_ net228 VGND VGND VPWR VPWR _2073_
+ sky130_fd_sc_hd__o21ai_1
X_3114_ _1390_ _1412_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3045_ _1346_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__nand2b_1
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3947_ _1979_ _1989_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3878_ _0623_ _1950_ _1954_ _1960_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__or4_1
X_2829_ cordic_inst.cordic_inst.y\[16\] cordic_inst.cordic_inst.y\[17\] cordic_inst.cordic_inst.y\[18\]
+ cordic_inst.cordic_inst.y\[19\] net310 net299 VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_29_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ net359 _0058_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[14\] sky130_fd_sc_hd__dfxtp_1
X_3801_ _1899_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__inv_2
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4781_ net400 _0508_ _0203_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[10\] sky130_fd_sc_hd__dfrtp_2
X_3732_ net254 _1847_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__nand2_1
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3663_ cordic_inst.deg_handler_inst.theta_abs\[19\] net152 net149 _1810_ VGND VGND
+ VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
X_2614_ net154 _0758_ net250 VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__a21oi_1
X_3594_ cordic_inst.deg_handler_inst.theta_abs\[5\] _1761_ VGND VGND VPWR VPWR _1762_
+ sky130_fd_sc_hd__or2_1
X_2545_ net250 _0743_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nor2_1
X_2476_ cordic_inst.cordic_inst.y\[30\] _0809_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__or2_1
X_4215_ axi_controller.result_out\[22\] _2179_ net201 VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_1
XFILLER_18_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4146_ _2116_ _2118_ net229 VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__mux2_1
XFILLER_29_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4077_ cordic_inst.cordic_inst.cos_out\[5\] cordic_inst.cordic_inst.cos_out\[4\]
+ _2048_ net225 VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__o31a_1
X_3028_ _1329_ _1330_ _1313_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_26_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout240 _0607_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_4
Xfanout273 cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_4
Xfanout251 _0604_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_2
Xfanout262 cordic_inst.cordic_inst.y\[31\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout284 net287 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_2
Xfanout295 net296 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__buf_2
XFILLER_46_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2330_ net278 _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__nor2_1
X_2261_ cordic_inst.cordic_inst.y\[8\] VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__inv_2
X_4000_ _0621_ _2005_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nor2_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4902_ net371 _0030_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4833_ net384 _0560_ _0255_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[30\] sky130_fd_sc_hd__dfrtp_2
X_4764_ net393 _0491_ _0186_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3715_ cordic_inst.deg_handler_inst.theta_norm\[14\] cordic_inst.deg_handler_inst.theta_norm\[13\]
+ _1834_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_31_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4695_ net403 _0422_ _0117_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_3646_ _1768_ net147 _1801_ net150 cordic_inst.deg_handler_inst.theta_abs\[11\] VGND
+ VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a32o_1
X_3577_ cordic_inst.cordic_inst.x\[2\] cordic_inst.cordic_inst.cos_out\[2\] net208
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
X_2528_ cordic_inst.cordic_inst.y\[19\] _0847_ _0851_ _0596_ VGND VGND VPWR VPWR _0863_
+ sky130_fd_sc_hd__o2bb2a_1
X_2459_ net245 _0692_ _0630_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a21o_1
X_4129_ net225 _2103_ cordic_inst.cordic_inst.cos_out\[12\] VGND VGND VPWR VPWR _2104_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3500_ net175 _1718_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__nor2_1
XFILLER_7_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ net325 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__inv_2
X_3431_ _1474_ _1669_ net176 VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__a21oi_1
X_3362_ _1596_ _1599_ _1600_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__o21ai_1
X_2313_ cordic_inst.cordic_inst.x\[29\] cordic_inst.cordic_inst.x\[30\] net305 VGND
+ VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux2_1
X_3293_ _1515_ _1529_ _1530_ _1531_ _1526_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__o311a_1
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4816_ net405 _0543_ _0238_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[13\] sky130_fd_sc_hd__dfrtp_4
X_4747_ net400 _0474_ _0169_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4678_ net389 _0405_ _0100_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3629_ cordic_inst.deg_handler_inst.theta_abs\[3\] _1759_ VGND VGND VPWR VPWR _1793_
+ sky130_fd_sc_hd__nand2_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput105 wstrb[2] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ axi_controller.write_addr_reg\[29\] net57 net189 VGND VGND VPWR VPWR _0328_
+ sky130_fd_sc_hd__mux2_1
X_2931_ cordic_inst.cordic_inst.x\[29\] _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__nor2_1
XFILLER_31_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2862_ net216 _1120_ _1154_ _0713_ net276 VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a221o_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4601_ net370 _0333_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_1
X_2793_ cordic_inst.cordic_inst.y\[15\] cordic_inst.cordic_inst.y\[16\] cordic_inst.cordic_inst.y\[17\]
+ cordic_inst.cordic_inst.y\[18\] net310 net299 VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux4_1
X_4532_ net353 _0264_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[14\] sky130_fd_sc_hd__dfxtp_1
X_4463_ net335 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__inv_2
X_3414_ cordic_inst.cordic_inst.z\[19\] _1636_ _1640_ cordic_inst.cordic_inst.z\[18\]
+ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4394_ net317 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
X_3345_ _1511_ _0707_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__nand2b_1
X_3276_ _1506_ _1514_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__and2b_1
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3130_ _1335_ _1337_ _1423_ net177 VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__a31o_1
X_3061_ _1200_ _1363_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3963_ axi_controller.write_addr_reg\[12\] net39 net188 VGND VGND VPWR VPWR _0311_
+ sky130_fd_sc_hd__mux2_1
X_3894_ net75 _1965_ _1971_ net346 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__o211a_1
X_2914_ _1195_ _1198_ net271 VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__o21a_1
X_2845_ _1138_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__and2_1
XFILLER_31_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2776_ cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.y\[29\] cordic_inst.cordic_inst.y\[30\]
+ net263 net304 net295 VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__mux4_2
X_4515_ net326 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__inv_2
X_4446_ net327 VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__inv_2
X_4377_ net340 VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
X_3328_ net266 _1481_ _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__mux2_1
X_3259_ net237 net232 VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__nor2_1
XFILLER_27_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2630_ cordic_inst.cordic_inst.y\[13\] _0932_ _0928_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a21oi_1
XFILLER_40_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2561_ cordic_inst.cordic_inst.y\[0\] _0718_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__nand2_1
XFILLER_5_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4300_ net84 _2243_ _2249_ net348 VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o211a_1
X_2492_ _0800_ _0826_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__xnor2_1
X_4231_ _2192_ _2193_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__or2_1
X_4162_ net226 _2132_ cordic_inst.cordic_inst.cos_out\[16\] VGND VGND VPWR VPWR _2133_
+ sky130_fd_sc_hd__a21oi_1
X_4093_ cordic_inst.cordic_inst.cos_out\[7\] _2068_ net225 VGND VGND VPWR VPWR _2072_
+ sky130_fd_sc_hd__o21a_1
X_3113_ _1382_ _1397_ _1394_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__a21o_1
XFILLER_28_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3044_ cordic_inst.cordic_inst.x\[21\] _1345_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__nand2_1
XFILLER_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3946_ axi_controller.read_addr_reg\[17\] _1980_ _1988_ axi_controller.read_addr_reg\[2\]
+ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__or4b_1
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3877_ axi_controller.write_addr_reg\[5\] _1959_ axi_controller.write_addr_reg\[3\]
+ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_21_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2828_ net243 _1130_ _1124_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__o21ai_2
X_2759_ net183 _0901_ _1064_ net165 cordic_inst.cordic_inst.y\[2\] VGND VGND VPWR
+ VPWR _0532_ sky130_fd_sc_hd__a32o_1
X_4429_ net336 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
Xfanout400 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3800_ _1880_ _1898_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__or2_1
X_4780_ net397 _0507_ _0202_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3731_ cordic_inst.deg_handler_inst.theta_norm\[20\] cordic_inst.deg_handler_inst.theta_norm\[19\]
+ _1844_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__or3_1
XFILLER_14_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3662_ _1808_ _1809_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__nor2_1
X_2613_ _0940_ _0941_ _0947_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__or3_1
X_3593_ cordic_inst.deg_handler_inst.theta_abs\[4\] _1760_ VGND VGND VPWR VPWR _1761_
+ sky130_fd_sc_hd__or2_1
X_2544_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__inv_2
X_2475_ cordic_inst.cordic_inst.y\[30\] _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nand2_1
X_4214_ net316 _2177_ _2178_ _2174_ _2175_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__a32o_1
X_4145_ cordic_inst.cordic_inst.cos_out\[14\] _2117_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__xor2_1
XFILLER_18_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4076_ axi_controller.result_out\[5\] _2057_ net202 VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
XFILLER_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3027_ _1287_ _1294_ _1318_ _1323_ _1293_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_26_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3929_ axi_controller.read_addr_reg\[30\] net25 net195 VGND VGND VPWR VPWR _0296_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout241 _0607_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_2
Xfanout230 net231 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_2
Xfanout252 net253 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_2
Xfanout274 net279 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_4
Xfanout263 cordic_inst.cordic_inst.y\[31\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_4
Xfanout296 cordic_inst.cordic_inst.i\[1\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_2
Xfanout285 net287 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_4
XFILLER_43_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2260_ cordic_inst.cordic_inst.y\[10\] VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__inv_2
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4901_ net367 _0019_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4832_ net384 _0559_ _0254_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[29\] sky130_fd_sc_hd__dfrtp_4
X_4763_ net393 _0490_ _0185_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3714_ cordic_inst.deg_handler_inst.theta_norm\[14\] _1836_ VGND VGND VPWR VPWR _0013_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4694_ net403 _0421_ _0116_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3645_ cordic_inst.deg_handler_inst.theta_abs\[11\] _1767_ VGND VGND VPWR VPWR _1801_
+ sky130_fd_sc_hd__nand2_1
X_3576_ cordic_inst.cordic_inst.x\[3\] cordic_inst.cordic_inst.cos_out\[3\] net208
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_1
X_2527_ _0860_ _0861_ _0858_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__a21o_1
X_2458_ net278 _0749_ _0631_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__o21ai_2
X_2389_ net264 _0647_ _0648_ _0645_ net233 net232 VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__mux4_2
X_4128_ cordic_inst.cordic_inst.cos_out\[11\] cordic_inst.cordic_inst.cos_out\[10\]
+ _2089_ VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__or3_1
X_4059_ _2040_ _2042_ net230 VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__mux2_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap216 _0709_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
X_3430_ _1476_ _1477_ _1666_ _1668_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__o31ai_1
X_3361_ cordic_inst.cordic_inst.z\[2\] _1593_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__xor2_1
X_2312_ cordic_inst.cordic_inst.x\[27\] cordic_inst.cordic_inst.x\[28\] net304 VGND
+ VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3292_ _1518_ _1525_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__nand2_1
XFILLER_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4815_ net405 _0542_ _0237_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[12\] sky130_fd_sc_hd__dfrtp_2
X_4746_ net399 _0473_ _0168_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4677_ net389 _0404_ _0099_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3628_ _1759_ net148 _1792_ net150 cordic_inst.deg_handler_inst.theta_abs\[2\] VGND
+ VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a32o_1
X_3559_ cordic_inst.cordic_inst.x\[20\] cordic_inst.cordic_inst.cos_out\[20\] net214
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
Xinput106 wstrb[3] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2930_ _1226_ _1232_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2861_ _1159_ _1160_ _1163_ net243 VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__o22a_1
X_4600_ net365 _0332_ VGND VGND VPWR VPWR axi_controller.mode sky130_fd_sc_hd__dfxtp_2
X_2792_ cordic_inst.cordic_inst.y\[11\] cordic_inst.cordic_inst.y\[12\] cordic_inst.cordic_inst.y\[13\]
+ cordic_inst.cordic_inst.y\[14\] net310 net299 VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux4_1
X_4531_ net353 _0263_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4462_ net334 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__inv_2
X_3413_ _1651_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__inv_2
X_4393_ net317 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
X_3344_ net288 _1509_ net206 net280 VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__a211o_1
X_3275_ cordic_inst.cordic_inst.z\[12\] _1513_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__nand2_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4729_ net375 _0456_ _0151_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3060_ net250 _1201_ _1217_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__o21bai_1
XFILLER_23_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3962_ axi_controller.write_addr_reg\[11\] net38 net187 VGND VGND VPWR VPWR _0310_
+ sky130_fd_sc_hd__mux2_1
X_3893_ axi_controller.reg_input_data\[13\] _1964_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__or2_1
X_2913_ net271 _1195_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__and2_1
X_2844_ net286 _1141_ _1145_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__a211o_1
X_2775_ cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.y\[29\] net306 VGND
+ VGND VPWR VPWR _1078_ sky130_fd_sc_hd__mux2_1
X_4514_ net326 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__inv_2
X_4445_ net331 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__inv_2
X_4376_ net340 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
X_3327_ _1564_ _1565_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__and2_1
X_3258_ _1485_ _1488_ _1484_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__o21ba_1
X_3189_ _1278_ _1464_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__and2_1
XFILLER_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2560_ cordic_inst.cordic_inst.y\[1\] _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__nand2_1
X_2491_ _0630_ _0652_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__nor2_1
X_4230_ cordic_inst.cordic_inst.sin_out\[24\] net257 _2191_ VGND VGND VPWR VPWR _2193_
+ sky130_fd_sc_hd__and3_1
X_4161_ cordic_inst.cordic_inst.cos_out\[15\] cordic_inst.cordic_inst.cos_out\[14\]
+ cordic_inst.cordic_inst.cos_out\[13\] _2111_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__or4_2
X_4092_ net202 _2071_ _2064_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a21oi_1
X_3112_ net181 _1401_ _1411_ net163 cordic_inst.cordic_inst.x\[28\] VGND VGND VPWR
+ VPWR _0526_ sky130_fd_sc_hd__a32o_1
X_3043_ cordic_inst.cordic_inst.x\[21\] _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__nor2_1
XFILLER_36_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3945_ _0625_ _1982_ _1984_ _1985_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__or4_1
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3876_ _1955_ _1956_ _1957_ _1958_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2827_ net262 _1126_ _1128_ _1125_ net239 net233 VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux4_2
X_2758_ _0899_ _0900_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__or2_1
X_4428_ net334 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__inv_2
X_2689_ _0989_ _0990_ _1010_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a21o_1
Xfanout401 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__buf_2
X_4359_ net329 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3730_ cordic_inst.deg_handler_inst.theta_norm\[20\] _1846_ VGND VGND VPWR VPWR _0020_
+ sky130_fd_sc_hd__xnor2_1
X_3661_ cordic_inst.deg_handler_inst.theta_abs\[18\] cordic_inst.deg_handler_inst.theta_abs\[19\]
+ _1787_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__and3_1
X_2612_ _0945_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__or2_1
X_3592_ cordic_inst.deg_handler_inst.theta_abs\[3\] _1759_ VGND VGND VPWR VPWR _1760_
+ sky130_fd_sc_hd__or2_1
X_2543_ cordic_inst.cordic_inst.y\[6\] _0875_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__nand2_1
X_2474_ _0639_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__xnor2_1
X_4213_ cordic_inst.cordic_inst.sin_out\[22\] net257 _2176_ VGND VGND VPWR VPWR _2178_
+ sky130_fd_sc_hd__nand3_1
X_4144_ cordic_inst.cordic_inst.cos_out\[13\] _2111_ net227 VGND VGND VPWR VPWR _2117_
+ sky130_fd_sc_hd__o21a_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4075_ net314 _2053_ _2055_ _2056_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__a22o_1
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3026_ _1317_ _1321_ _1316_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_26_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3928_ axi_controller.read_addr_reg\[29\] net23 net195 VGND VGND VPWR VPWR _0295_
+ sky130_fd_sc_hd__mux2_1
X_3859_ _1932_ _1939_ _1941_ net107 net68 VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_6_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout220 _0680_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
Xfanout231 _0612_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_2
Xfanout253 net255 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_2
Xfanout242 _0606_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_4
Xfanout264 net265 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_2
Xfanout286 net287 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_2
Xfanout297 net300 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__buf_2
Xfanout275 net276 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_2
XFILLER_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4900_ net367 cordic_inst.deg_handler_inst.theta_norm\[0\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4831_ net384 _0558_ _0253_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[28\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4762_ net392 _0489_ _0184_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3713_ cordic_inst.deg_handler_inst.theta_norm\[13\] _1834_ net253 VGND VGND VPWR
+ VPWR _1836_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_31_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4693_ net404 _0420_ _0115_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_3644_ _1767_ net147 _1800_ net150 cordic_inst.deg_handler_inst.theta_abs\[10\] VGND
+ VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3575_ cordic_inst.cordic_inst.x\[4\] cordic_inst.cordic_inst.cos_out\[4\] net211
+ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux2_1
X_2526_ cordic_inst.cordic_inst.y\[17\] _0857_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nand2_1
X_2457_ _0631_ _0790_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__nand2_1
XFILLER_29_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2388_ net232 _0648_ _0633_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a21o_1
XFILLER_29_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4127_ net228 _2100_ _2101_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__or3_1
X_4058_ cordic_inst.cordic_inst.cos_out\[3\] _2041_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__xor2_1
X_3009_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap217 _0708_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
Xmax_cap206 _1502_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_1
X_3360_ _1597_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_27_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2311_ cordic_inst.cordic_inst.x\[23\] cordic_inst.cordic_inst.x\[24\] cordic_inst.cordic_inst.x\[25\]
+ cordic_inst.cordic_inst.x\[26\] net307 net301 VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux4_1
X_3291_ cordic_inst.cordic_inst.z\[13\] _1505_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__nor2_1
XFILLER_38_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4814_ net405 _0541_ _0236_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[11\] sky130_fd_sc_hd__dfrtp_2
X_4745_ net396 _0472_ _0167_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4676_ net391 _0403_ _0098_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3627_ cordic_inst.deg_handler_inst.theta_abs\[2\] _1758_ VGND VGND VPWR VPWR _1792_
+ sky130_fd_sc_hd__nand2_1
X_3558_ cordic_inst.cordic_inst.x\[21\] cordic_inst.cordic_inst.cos_out\[21\] net214
+ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2509_ _0832_ _0837_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__or3_1
Xinput107 wvalid VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
X_3489_ cordic_inst.cordic_inst.angle\[17\] net172 net159 cordic_inst.cordic_inst.z\[17\]
+ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2860_ _1161_ _1162_ net283 VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__mux2_1
XFILLER_31_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2791_ _1084_ _1093_ net235 VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__mux2_1
X_4530_ net353 _0262_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4461_ net334 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__inv_2
X_3412_ _1632_ _1647_ _1645_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__o21a_1
X_4392_ net317 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
X_3343_ net281 _1577_ _1580_ _1511_ _1522_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__o32a_1
X_3274_ net267 _1507_ _1512_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__mux2_1
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2989_ _1182_ _1291_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4728_ net378 _0455_ _0150_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[21\] sky130_fd_sc_hd__dfrtp_1
X_4659_ net377 _0389_ _0091_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3961_ axi_controller.write_addr_reg\[10\] net37 net187 VGND VGND VPWR VPWR _0309_
+ sky130_fd_sc_hd__mux2_1
X_2912_ net272 _1189_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__nand2_1
X_3892_ net74 _1965_ _1970_ net347 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o211a_1
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2843_ cordic_inst.cordic_inst.y\[0\] net221 _0711_ _1143_ net219 VGND VGND VPWR
+ VPWR _1146_ sky130_fd_sc_hd__a32o_1
XFILLER_31_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2774_ net242 _1076_ net215 VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__a21o_1
X_4513_ net327 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__inv_2
X_4444_ net331 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__inv_2
X_4375_ net341 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
X_3326_ _1498_ _1558_ _0706_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__o21ai_1
X_3257_ _1486_ _1490_ _1495_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__or3_1
X_3188_ _1260_ _1263_ _1277_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__nand3_1
XFILLER_26_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2490_ _0823_ _0824_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__and2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4160_ cordic_inst.cordic_inst.sin_out\[16\] net260 _2128_ _2130_ VGND VGND VPWR
+ VPWR _2131_ sky130_fd_sc_hd__a31o_1
X_3111_ _1240_ _1396_ _1398_ _1400_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__or4_1
X_4091_ net229 _2066_ _2067_ _2069_ _2070_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__o32a_1
X_3042_ _1207_ _1344_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3944_ axi_controller.read_addr_reg\[25\] _1981_ _1983_ _1986_ VGND VGND VPWR VPWR
+ _1987_ sky130_fd_sc_hd__nor4_1
X_3875_ axi_controller.write_addr_reg\[17\] axi_controller.write_addr_reg\[16\] axi_controller.write_addr_reg\[19\]
+ axi_controller.write_addr_reg\[18\] VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__or4_1
X_2826_ net237 _1128_ _1071_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_21_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2757_ net185 _0905_ _1063_ net168 cordic_inst.cordic_inst.y\[3\] VGND VGND VPWR
+ VPWR _0533_ sky130_fd_sc_hd__a32o_1
X_2688_ _0989_ _0990_ _1010_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__nand3_1
X_4427_ net334 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__inv_2
Xfanout402 net408 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_2
X_4358_ net329 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
X_4289_ axi_controller.reg_input_data\[16\] _2242_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__or2_1
X_3309_ net288 _0706_ _0712_ net222 _0705_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_1_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3660_ cordic_inst.deg_handler_inst.theta_abs\[18\] _1787_ cordic_inst.deg_handler_inst.theta_abs\[19\]
+ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__a21oi_2
X_2611_ _0597_ _0944_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__and2_1
X_3591_ cordic_inst.deg_handler_inst.theta_abs\[0\] cordic_inst.deg_handler_inst.theta_abs\[1\]
+ cordic_inst.deg_handler_inst.theta_abs\[2\] VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__or3_1
X_2542_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__inv_2
X_4212_ net257 _2176_ cordic_inst.cordic_inst.sin_out\[22\] VGND VGND VPWR VPWR _2177_
+ sky130_fd_sc_hd__a21o_1
X_2473_ net269 _0807_ _0806_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a21oi_1
X_4143_ cordic_inst.cordic_inst.sin_out\[14\] _2115_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__xor2_1
X_4074_ cordic_inst.cordic_inst.cos_out\[5\] _2054_ net314 VGND VGND VPWR VPWR _2056_
+ sky130_fd_sc_hd__a21oi_1
X_3025_ _1304_ _1307_ _1326_ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3927_ axi_controller.read_addr_reg\[28\] net22 net197 VGND VGND VPWR VPWR _0294_
+ sky130_fd_sc_hd__mux2_1
X_3858_ net47 net36 _1933_ _1940_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__or4_1
X_3789_ axi_controller.reg_input_data\[20\] axi_controller.reg_input_data\[19\] axi_controller.reg_input_data\[22\]
+ axi_controller.reg_input_data\[21\] VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__o211a_1
X_2809_ cordic_inst.cordic_inst.y\[26\] cordic_inst.cordic_inst.y\[27\] net306 VGND
+ VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout210 net211 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_4
Xfanout221 net222 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_2
Xfanout232 _0609_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_4
Xfanout254 net255 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_2
Xfanout243 net247 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_4
Xfanout265 cordic_inst.cordic_inst.x\[31\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_4
Xfanout287 cordic_inst.cordic_inst.i\[3\] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_2
Xfanout298 net300 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_1
Xfanout276 net279 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4830_ net393 _0557_ _0252_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[27\] sky130_fd_sc_hd__dfrtp_4
X_4761_ net394 _0488_ _0183_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_3712_ cordic_inst.deg_handler_inst.theta_norm\[13\] _1835_ VGND VGND VPWR VPWR _0012_
+ sky130_fd_sc_hd__xnor2_1
X_4692_ net405 _0419_ _0114_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_3643_ cordic_inst.deg_handler_inst.theta_abs\[10\] _1766_ VGND VGND VPWR VPWR _1800_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3574_ cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.cos_out\[5\] net211
+ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux2_1
X_2525_ cordic_inst.cordic_inst.y\[16\] _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__nand2_1
X_2456_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__inv_2
X_4126_ net259 _2099_ cordic_inst.cordic_inst.sin_out\[12\] VGND VGND VPWR VPWR _2101_
+ sky130_fd_sc_hd__a21oi_1
X_2387_ _0645_ _0647_ net301 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux2_1
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4057_ cordic_inst.cordic_inst.cos_out\[2\] cordic_inst.cordic_inst.cos_out\[1\]
+ cordic_inst.cordic_inst.cos_out\[0\] net223 VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__o31a_1
X_3008_ cordic_inst.cordic_inst.x\[12\] _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4959_ net398 _0588_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_1
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3290_ _1528_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__inv_2
X_2310_ cordic_inst.cordic_inst.x\[25\] cordic_inst.cordic_inst.x\[26\] net307 VGND
+ VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux2_1
XFILLER_26_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4813_ net405 _0540_ _0235_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_34_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4744_ net396 _0471_ _0166_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4675_ net389 _0402_ _0097_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3626_ _1758_ net148 _1791_ net151 cordic_inst.deg_handler_inst.theta_abs\[1\] VGND
+ VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a32o_1
X_3557_ cordic_inst.cordic_inst.x\[22\] cordic_inst.cordic_inst.cos_out\[22\] net208
+ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
X_2508_ _0841_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3488_ _1632_ _1648_ _1705_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__or3_1
X_2439_ net286 _0754_ _0637_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__o21a_1
X_4109_ cordic_inst.cordic_inst.sin_out\[9\] cordic_inst.cordic_inst.sin_out\[8\]
+ cordic_inst.cordic_inst.sin_out\[7\] _2065_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__or4_1
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_44_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2790_ cordic_inst.cordic_inst.y\[19\] cordic_inst.cordic_inst.y\[20\] cordic_inst.cordic_inst.y\[21\]
+ cordic_inst.cordic_inst.y\[22\] net307 net300 VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__mux4_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4460_ net329 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__inv_2
X_3411_ _1532_ _1628_ _1649_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__a21o_1
X_4391_ net317 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
X_3342_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__inv_2
X_3273_ _1510_ _1511_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__nand2b_1
XFILLER_38_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2988_ _1180_ _1184_ net272 VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__o21ai_1
X_4727_ net377 _0454_ _0149_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[20\] sky130_fd_sc_hd__dfrtp_1
X_4658_ net377 _0388_ _0090_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[2\] sky130_fd_sc_hd__dfrtp_1
X_3609_ cordic_inst.deg_handler_inst.theta_abs\[28\] cordic_inst.deg_handler_inst.theta_abs\[29\]
+ cordic_inst.deg_handler_inst.theta_abs\[30\] cordic_inst.deg_handler_inst.theta_abs\[31\]
+ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__or4_1
Xinput90 wdata[27] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
X_4589_ net382 _0321_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3960_ axi_controller.write_addr_reg\[9\] net67 net187 VGND VGND VPWR VPWR _0308_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2911_ _1070_ _1092_ net274 VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__a21oi_1
X_3891_ axi_controller.reg_input_data\[12\] _1964_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__or2_1
X_2842_ cordic_inst.cordic_inst.y\[1\] net217 _0709_ _1144_ net275 VGND VGND VPWR
+ VPWR _1145_ sky130_fd_sc_hd__a221o_1
X_2773_ net241 _1075_ _1070_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__a21bo_1
X_4512_ net327 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__inv_2
X_4443_ net333 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__inv_2
X_4374_ net341 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
X_3325_ net281 _0707_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__or2_1
X_3256_ _1491_ _1492_ _1494_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__or3b_1
X_3187_ cordic_inst.cordic_inst.x\[5\] net158 _1462_ _1463_ VGND VGND VPWR VPWR _0503_
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ net179 _1409_ _1410_ net163 cordic_inst.cordic_inst.x\[29\] VGND VGND VPWR
+ VPWR _0527_ sky130_fd_sc_hd__a32o_1
X_4090_ cordic_inst.cordic_inst.cos_out\[7\] net225 _2068_ net314 VGND VGND VPWR VPWR
+ _2070_ sky130_fd_sc_hd__a31o_1
X_3041_ net251 _1208_ _1218_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__o21bai_1
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3943_ axi_controller.read_addr_reg\[20\] axi_controller.read_addr_reg\[23\] axi_controller.read_addr_reg\[22\]
+ _1984_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__or4_1
X_3874_ axi_controller.write_addr_reg\[25\] axi_controller.write_addr_reg\[24\] axi_controller.write_addr_reg\[27\]
+ axi_controller.write_addr_reg\[26\] VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__or4_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2825_ net232 _1086_ _1072_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_21_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2756_ _0902_ _0904_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__or2_1
X_2687_ cordic_inst.cordic_inst.y\[26\] net169 _1015_ _1016_ VGND VGND VPWR VPWR _0556_
+ sky130_fd_sc_hd__a22o_1
X_4426_ net334 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__inv_2
Xfanout403 net404 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_2
X_4357_ net322 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
X_4288_ net105 _1963_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__nand2_2
X_3308_ _1540_ _1546_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__nor2_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3239_ net248 cordic_inst.cordic_inst.z\[24\] VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__nand2_1
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2610_ _0597_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__nor2_1
X_3590_ cordic_inst.deg_handler_inst.theta_abs\[0\] cordic_inst.deg_handler_inst.theta_abs\[1\]
+ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__or2_1
X_2541_ cordic_inst.cordic_inst.y\[6\] _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nor2_1
X_2472_ net274 _0774_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__nor2_1
X_4211_ cordic_inst.cordic_inst.sin_out\[21\] _2169_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__or2_1
X_4142_ cordic_inst.cordic_inst.sin_out\[13\] _2107_ net261 VGND VGND VPWR VPWR _2115_
+ sky130_fd_sc_hd__o21a_1
X_4073_ cordic_inst.cordic_inst.cos_out\[5\] _2054_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__or2_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3024_ _1298_ _1302_ _1297_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3926_ axi_controller.read_addr_reg\[27\] net21 net195 VGND VGND VPWR VPWR _0293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3857_ net39 net42 net41 _1934_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__or4_1
X_3788_ axi_controller.reg_input_data\[22\] _1889_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__xnor2_1
X_2808_ cordic_inst.cordic_inst.y\[22\] cordic_inst.cordic_inst.y\[23\] cordic_inst.cordic_inst.y\[24\]
+ cordic_inst.cordic_inst.y\[25\] net307 net301 VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__mux4_1
X_2739_ net177 _1039_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout211 net213 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_4
X_4409_ net321 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
Xfanout222 _0678_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_2
Xfanout200 net201 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
Xfanout255 cordic_inst.deg_handler_inst.theta_norm\[31\] VGND VGND VPWR VPWR net255
+ sky130_fd_sc_hd__clkbuf_2
Xfanout233 net234 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 net246 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_4
Xfanout266 net267 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_2
Xfanout288 net289 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_2
Xfanout277 net279 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_2
Xfanout299 net300 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_2
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4760_ net395 _0487_ _0182_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3711_ net253 _1834_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__nand2_1
X_4691_ net405 _0418_ _0113_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3642_ _1766_ net148 _1799_ net150 cordic_inst.deg_handler_inst.theta_abs\[9\] VGND
+ VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3573_ cordic_inst.cordic_inst.x\[6\] cordic_inst.cordic_inst.cos_out\[6\] net210
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
X_2524_ _0785_ _0855_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__xor2_1
X_2455_ net245 _0755_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__nand2_1
X_2386_ _0719_ _0720_ net290 VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux2_1
X_4125_ cordic_inst.cordic_inst.sin_out\[12\] net258 _2099_ VGND VGND VPWR VPWR _2100_
+ sky130_fd_sc_hd__and3_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4056_ cordic_inst.cordic_inst.sin_out\[3\] _2039_ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__xor2_1
X_3007_ _1190_ _1215_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__xor2_2
XFILLER_25_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4958_ net399 _0587_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_1
X_4889_ net358 _0042_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_3909_ axi_controller.read_addr_reg\[10\] net3 net196 VGND VGND VPWR VPWR _0276_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4812_ net401 _0539_ _0234_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[9\] sky130_fd_sc_hd__dfrtp_4
X_4743_ net396 _0470_ _0165_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4674_ net375 _0401_ _0096_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.done sky130_fd_sc_hd__dfrtp_1
X_3625_ cordic_inst.deg_handler_inst.theta_abs\[0\] cordic_inst.deg_handler_inst.theta_abs\[1\]
+ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__nand2_1
XFILLER_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3556_ cordic_inst.cordic_inst.x\[23\] cordic_inst.cordic_inst.cos_out\[23\] net208
+ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
X_2507_ cordic_inst.cordic_inst.y\[21\] _0840_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__or2_1
X_3487_ _1632_ _1705_ _1648_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__o21ai_1
X_2438_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__inv_2
X_2369_ cordic_inst.cordic_inst.x\[4\] cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.x\[6\]
+ cordic_inst.cordic_inst.x\[7\] net311 net300 VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__mux4_1
X_4108_ axi_controller.result_out\[10\] net203 VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__nor2_1
X_4039_ axi_controller.reg_input_data\[7\] _2018_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__or2_1
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3410_ _1647_ _1642_ _1634_ _1645_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__or4bb_1
X_4390_ net317 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
X_3341_ net293 net295 net306 VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__and3_1
X_3272_ net289 net294 net280 VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2987_ _1244_ _1247_ _1282_ _1289_ _1243_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a311o_1
X_4726_ net377 _0453_ _0148_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[19\] sky130_fd_sc_hd__dfrtp_1
X_4657_ net377 _0387_ _0089_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[1\] sky130_fd_sc_hd__dfrtp_1
X_3608_ cordic_inst.deg_handler_inst.theta_abs\[19\] cordic_inst.deg_handler_inst.theta_abs\[20\]
+ _1775_ cordic_inst.deg_handler_inst.theta_abs\[21\] VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__a31o_1
Xinput91 wdata[28] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
Xinput80 wdata[18] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
X_4588_ net380 _0320_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3539_ _1596_ _1599_ _1600_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__or3_1
XFILLER_45_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2910_ net242 _1186_ net215 VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__a21o_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3890_ net73 _1965_ _1969_ net347 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__o211a_1
X_2841_ cordic_inst.cordic_inst.y\[2\] cordic_inst.cordic_inst.y\[3\] net311 VGND
+ VGND VPWR VPWR _1144_ sky130_fd_sc_hd__mux2_1
XFILLER_12_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2772_ net237 _1074_ _1071_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__a21o_1
X_4511_ net331 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__inv_2
X_4442_ net333 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__inv_2
X_4373_ net342 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
X_3324_ _1561_ _1562_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__or2_1
X_3255_ net268 cordic_inst.cordic_inst.z\[23\] VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__xnor2_1
X_3186_ _1279_ _1280_ net177 VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__a21o_1
XFILLER_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4709_ net379 _0436_ _0131_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3040_ _1341_ _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__nand2_1
XFILLER_24_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3942_ axi_controller.read_addr_reg\[20\] axi_controller.read_addr_reg\[23\] axi_controller.read_addr_reg\[22\]
+ axi_controller.read_addr_reg\[25\] VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__or4_1
X_3873_ axi_controller.write_addr_reg\[28\] axi_controller.write_addr_reg\[29\] axi_controller.write_addr_reg\[30\]
+ axi_controller.write_addr_reg\[31\] VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__nand4_1
X_2824_ _1125_ _1126_ net291 VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__mux2_1
X_2755_ net185 _0909_ _1062_ net168 cordic_inst.cordic_inst.y\[4\] VGND VGND VPWR
+ VPWR _0534_ sky130_fd_sc_hd__a32o_1
X_2686_ net176 _1012_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__nor2_1
X_4425_ net329 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
X_4356_ net318 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
Xfanout404 net408 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_2
X_3307_ _1544_ _1545_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__nand2b_1
X_4287_ net105 _1963_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__and2_1
X_3238_ net268 cordic_inst.cordic_inst.z\[28\] VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__xor2_1
XFILLER_39_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _1321_ _1441_ _1318_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__a21boi_1
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2540_ _0693_ _0870_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2471_ _0644_ _0805_ net269 VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__o21a_1
X_4210_ cordic_inst.cordic_inst.cos_out\[22\] net224 _2173_ net316 VGND VGND VPWR
+ VPWR _2175_ sky130_fd_sc_hd__a31oi_1
X_4141_ axi_controller.result_out\[13\] _2114_ net204 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux2_1
X_4072_ cordic_inst.cordic_inst.cos_out\[4\] _2048_ net225 VGND VGND VPWR VPWR _2054_
+ sky130_fd_sc_hd__o21a_1
X_3023_ cordic_inst.cordic_inst.x\[13\] _1306_ _1310_ cordic_inst.cordic_inst.x\[12\]
+ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__a22o_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3925_ axi_controller.read_addr_reg\[26\] net20 net197 VGND VGND VPWR VPWR _0292_
+ sky130_fd_sc_hd__mux2_1
X_3856_ _1935_ _1936_ _1937_ _1938_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__or4b_1
X_3787_ axi_controller.reg_input_data\[21\] _1880_ _1883_ _1887_ VGND VGND VPWR VPWR
+ _1889_ sky130_fd_sc_hd__o31a_1
X_2807_ net283 _1106_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a21o_1
XFILLER_3_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2738_ _0947_ _1038_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__nand2_1
X_4408_ net320 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
X_2669_ _0810_ _1000_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__a21oi_1
Xfanout201 cordic_inst.sign_handler_inst.done_pulse VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout223 _0613_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_4
Xfanout212 net213 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_4
X_4339_ net138 net191 net155 axi_controller.result_out\[4\] VGND VGND VPWR VPWR _0590_
+ sky130_fd_sc_hd__a22o_1
Xfanout234 net236 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_4
Xfanout245 net246 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout256 net257 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_2
Xfanout267 cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__buf_2
Xfanout289 net293 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout278 net279 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3710_ cordic_inst.deg_handler_inst.theta_norm\[12\] _1832_ VGND VGND VPWR VPWR _1834_
+ sky130_fd_sc_hd__or2_1
X_4690_ net405 _0417_ _0112_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3641_ cordic_inst.deg_handler_inst.theta_abs\[9\] _1765_ VGND VGND VPWR VPWR _1799_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3572_ cordic_inst.cordic_inst.x\[7\] cordic_inst.cordic_inst.cos_out\[7\] net210
+ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux2_1
X_2523_ cordic_inst.cordic_inst.y\[17\] _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__nor2_1
X_2454_ _0771_ _0781_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__or3_2
X_2385_ cordic_inst.cordic_inst.x\[21\] cordic_inst.cordic_inst.x\[22\] cordic_inst.cordic_inst.x\[23\]
+ cordic_inst.cordic_inst.x\[24\] net312 net301 VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux4_1
X_4124_ cordic_inst.cordic_inst.sin_out\[11\] cordic_inst.cordic_inst.sin_out\[10\]
+ _2086_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__or3_1
Xinput1 aclk VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_4055_ cordic_inst.cordic_inst.sin_out\[2\] cordic_inst.cordic_inst.sin_out\[1\]
+ cordic_inst.cordic_inst.sin_out\[0\] net261 VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__o31a_1
X_3006_ _1307_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__and2_1
X_4957_ net402 _0586_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_1
X_3908_ axi_controller.read_addr_reg\[9\] net33 net195 VGND VGND VPWR VPWR _0275_
+ sky130_fd_sc_hd__mux2_1
X_4888_ net358 _0041_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3839_ _1924_ _1925_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__or2_1
XFILLER_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4811_ net401 _0538_ _0233_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[8\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_16_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4742_ net391 _0469_ _0164_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4673_ net381 _0400_ _0095_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.start sky130_fd_sc_hd__dfrtp_1
X_3624_ net149 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
X_3555_ cordic_inst.cordic_inst.x\[24\] cordic_inst.cordic_inst.cos_out\[24\] net209
+ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
X_3486_ cordic_inst.cordic_inst.angle\[18\] net172 net159 cordic_inst.cordic_inst.z\[18\]
+ _1711_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__a221o_1
X_2506_ cordic_inst.cordic_inst.y\[21\] _0840_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nand2_1
X_2437_ net264 _0642_ _0747_ _0744_ net240 net245 VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__mux4_2
X_2368_ cordic_inst.cordic_inst.x\[4\] cordic_inst.cordic_inst.x\[5\] net312 VGND
+ VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux2_1
X_4107_ axi_controller.result_out\[9\] _2084_ net202 VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__mux2_1
X_2299_ _0609_ _0632_ _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__a21o_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4038_ net99 _2019_ _2026_ net350 VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__o211a_1
XFILLER_37_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3340_ net281 _1521_ _1578_ net220 _1500_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__a32o_1
XFILLER_3_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3271_ net222 _0707_ _1509_ net220 VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__a22o_1
XFILLER_38_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2986_ _1287_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__nand2_1
X_4725_ net374 _0452_ _0147_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[18\] sky130_fd_sc_hd__dfrtp_1
X_4656_ net377 _0386_ _0088_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[0\] sky130_fd_sc_hd__dfrtp_1
Xinput70 rready VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
X_4587_ net380 _0319_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[20\] sky130_fd_sc_hd__dfxtp_1
X_3607_ _0615_ _1774_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__nand2_1
Xinput81 wdata[19] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
Xinput92 wdata[29] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
X_3538_ net175 _1602_ _1747_ _1748_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__o31ai_1
XFILLER_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3469_ cordic_inst.cordic_inst.angle\[22\] net173 net161 cordic_inst.cordic_inst.z\[22\]
+ _1698_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a221o_1
XFILLER_17_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2840_ cordic_inst.cordic_inst.y\[4\] cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.y\[6\]
+ cordic_inst.cordic_inst.y\[7\] net308 net297 VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__mux4_2
X_2771_ net232 _1073_ _1072_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__a21o_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4510_ net331 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__inv_2
X_4441_ net333 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4372_ net341 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
X_3323_ cordic_inst.cordic_inst.z\[6\] _1560_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__nor2_1
X_3254_ _1491_ _1492_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__or2_1
X_3185_ _1279_ _1280_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__nor2_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2969_ _1270_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__nand2b_1
X_4708_ net379 _0435_ _0130_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4639_ net407 _0370_ net343 VGND VGND VPWR VPWR axi_controller.result_out\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3941_ axi_controller.read_addr_reg\[24\] axi_controller.read_addr_reg\[27\] axi_controller.read_addr_reg\[26\]
+ axi_controller.read_addr_reg\[28\] VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__or4b_1
X_3872_ axi_controller.write_addr_reg\[21\] axi_controller.write_addr_reg\[20\] axi_controller.write_addr_reg\[23\]
+ axi_controller.write_addr_reg\[22\] VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__or4_1
X_2823_ _1083_ _1085_ net295 VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__mux2_1
XFILLER_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2754_ _0906_ _0907_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__or2_1
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2685_ _0986_ _1011_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__or2_1
X_4424_ net330 VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__inv_2
X_4355_ net323 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout405 net406 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_2
X_3306_ cordic_inst.cordic_inst.z\[10\] _1543_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__or2_1
X_4286_ _2240_ _2241_ axi_controller.result_out\[31\] net200 VGND VGND VPWR VPWR _0385_
+ sky130_fd_sc_hd__o2bb2a_1
X_3237_ _1475_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__inv_2
X_3168_ cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.next_state\[1\] _1451_
+ net178 VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_1_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3099_ _1236_ _1238_ _1401_ _1234_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_40_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2470_ net270 _0798_ _0804_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a21o_1
X_4140_ _2112_ _2113_ _2110_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__o21ai_1
X_4071_ cordic_inst.cordic_inst.sin_out\[5\] _2052_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__xnor2_1
X_3022_ _1290_ _1295_ _1313_ _1324_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__or4bb_1
X_3924_ axi_controller.read_addr_reg\[25\] net19 net197 VGND VGND VPWR VPWR _0291_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3855_ net56 net57 net59 net60 VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__and4_1
X_3786_ _1887_ _1888_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and2_1
X_2806_ net218 _1107_ _1108_ net221 net277 VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a221o_1
X_2737_ net184 _1050_ _1051_ net166 cordic_inst.cordic_inst.y\[11\] VGND VGND VPWR
+ VPWR _0541_ sky130_fd_sc_hd__a32o_1
X_2668_ _1001_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__xor2_1
X_4407_ net320 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout202 net203 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__buf_2
Xfanout213 net214 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_2
X_2599_ cordic_inst.cordic_inst.y\[13\] _0932_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__and2_1
Xfanout224 _0613_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
X_4338_ net139 net191 net155 axi_controller.result_out\[5\] VGND VGND VPWR VPWR _0589_
+ sky130_fd_sc_hd__a22o_1
Xfanout235 net236 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net247 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
Xfanout268 cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__buf_4
Xfanout279 cordic_inst.cordic_inst.i\[4\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_2
X_4269_ cordic_inst.cordic_inst.cos_out\[28\] net223 _2218_ cordic_inst.cordic_inst.cos_out\[29\]
+ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__a211o_1
Xfanout257 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_2
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _1765_ net148 _1798_ net150 cordic_inst.deg_handler_inst.theta_abs\[8\] VGND
+ VGND VPWR VPWR _0083_ sky130_fd_sc_hd__a32o_1
X_3571_ cordic_inst.cordic_inst.x\[8\] cordic_inst.cordic_inst.cos_out\[8\] net210
+ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2522_ _0784_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2453_ _0665_ _0667_ _0786_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__or3b_1
X_2384_ cordic_inst.cordic_inst.x\[17\] cordic_inst.cordic_inst.x\[18\] cordic_inst.cordic_inst.x\[19\]
+ cordic_inst.cordic_inst.x\[20\] net310 net299 VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__mux4_1
X_4123_ axi_controller.result_out\[11\] _2098_ net203 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
X_4054_ axi_controller.result_out\[2\] _2038_ net203 VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
Xinput2 araddr[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_3005_ cordic_inst.cordic_inst.x\[13\] _1306_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__nand2_1
XFILLER_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4956_ net402 _0585_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_1
X_4887_ net358 _0040_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_3907_ axi_controller.read_addr_reg\[8\] net32 net195 VGND VGND VPWR VPWR _0274_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3838_ net145 axi_controller.state\[1\] net70 _1921_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_30_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3769_ axi_controller.reg_input_data\[24\] _1873_ axi_controller.reg_input_data\[31\]
+ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__o21bai_2
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ net397 _0537_ _0232_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4741_ net391 _0468_ _0163_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4672_ net377 net158 _0094_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3623_ _1785_ _1789_ _1780_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__a21oi_1
X_3554_ cordic_inst.cordic_inst.x\[25\] cordic_inst.cordic_inst.cos_out\[25\] net207
+ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
X_3485_ _1706_ _1710_ net179 VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__and3b_1
X_2505_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__inv_2
X_2436_ net154 _0758_ _0765_ _0769_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__nand4_2
X_2367_ _0700_ _0701_ net292 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__mux2_1
XFILLER_29_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4106_ _2083_ _2082_ _2080_ net228 VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__a2bb2o_1
X_2298_ net264 net295 VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__and2_1
X_4037_ axi_controller.reg_input_data\[6\] _2018_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4939_ net387 _0568_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_1
XFILLER_20_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3270_ net294 net303 VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__xor2_1
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2985_ cordic_inst.cordic_inst.x\[8\] _1286_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__or2_1
X_4724_ net374 _0451_ _0146_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[17\] sky130_fd_sc_hd__dfrtp_1
X_4655_ net381 net200 net317 VGND VGND VPWR VPWR axi_controller.done sky130_fd_sc_hd__dfrtp_1
Xinput60 awaddr[31] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
Xinput82 wdata[1] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
Xinput71 wdata[0] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
X_4586_ net380 _0318_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[19\] sky130_fd_sc_hd__dfxtp_1
X_3606_ cordic_inst.deg_handler_inst.theta_abs\[17\] _1773_ VGND VGND VPWR VPWR _1774_
+ sky130_fd_sc_hd__nand2_1
Xinput93 wdata[2] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
X_3537_ cordic_inst.cordic_inst.angle\[3\] net171 net160 cordic_inst.cordic_inst.z\[3\]
+ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__a22oi_1
X_3468_ _1693_ _1697_ net180 VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__and3b_1
X_3399_ cordic_inst.cordic_inst.z\[19\] _1636_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__nand2_1
X_2419_ net233 _0723_ _0635_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2770_ cordic_inst.cordic_inst.y\[30\] net263 net306 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__mux2_1
X_4440_ net340 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__inv_2
X_4371_ net341 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
X_3322_ cordic_inst.cordic_inst.z\[6\] _1560_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__and2_1
X_3253_ net248 cordic_inst.cordic_inst.z\[22\] VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__nor2_1
X_3184_ net183 _1461_ net158 cordic_inst.cordic_inst.x\[6\] VGND VGND VPWR VPWR _0504_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2968_ cordic_inst.cordic_inst.x\[1\] _1268_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__xor2_1
X_4707_ net379 _0434_ _0129_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[0\] sky130_fd_sc_hd__dfrtp_1
X_2899_ _1199_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nand2_1
X_4638_ net406 _0369_ net342 VGND VGND VPWR VPWR axi_controller.result_out\[15\] sky130_fd_sc_hd__dfrtp_1
X_4569_ net364 _0301_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3940_ _0625_ _1982_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__or2_1
X_3871_ axi_controller.write_addr_reg\[12\] axi_controller.write_addr_reg\[15\] axi_controller.write_addr_reg\[14\]
+ _1951_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__or4_1
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2822_ cordic_inst.cordic_inst.y\[21\] cordic_inst.cordic_inst.y\[22\] cordic_inst.cordic_inst.y\[23\]
+ cordic_inst.cordic_inst.y\[24\] net307 net301 VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__mux4_1
XFILLER_32_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2753_ cordic_inst.cordic_inst.y\[5\] net168 _1061_ net185 VGND VGND VPWR VPWR _0535_
+ sky130_fd_sc_hd__a22o_1
X_2684_ cordic_inst.cordic_inst.y\[27\] net163 _1014_ net181 VGND VGND VPWR VPWR _0557_
+ sky130_fd_sc_hd__a22o_1
X_4423_ net330 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__inv_2
X_4354_ net322 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
X_3305_ cordic_inst.cordic_inst.z\[10\] _1543_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__and2_1
Xfanout406 net407 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_2
X_4285_ net313 _2236_ _2237_ net200 VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__o31a_1
X_3236_ net268 cordic_inst.cordic_inst.z\[29\] VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3167_ _1312_ _1442_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3098_ _1396_ _1398_ _1400_ _1240_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__o31ai_4
XFILLER_35_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4070_ cordic_inst.cordic_inst.sin_out\[4\] _2045_ net259 VGND VGND VPWR VPWR _2052_
+ sky130_fd_sc_hd__o21ai_1
X_3021_ _1318_ _1323_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__nor2_1
XFILLER_37_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3923_ axi_controller.read_addr_reg\[24\] net18 net195 VGND VGND VPWR VPWR _0290_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3854_ net53 net52 net55 net54 VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__or4_1
X_2805_ cordic_inst.cordic_inst.y\[6\] cordic_inst.cordic_inst.y\[7\] cordic_inst.cordic_inst.y\[8\]
+ cordic_inst.cordic_inst.y\[9\] net308 net297 VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__mux4_1
X_3785_ _1884_ _1885_ _1886_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__or3_1
X_2736_ _0942_ _0945_ _1039_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__or3_1
X_2667_ net263 net265 VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__xnor2_2
X_4406_ net320 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
Xfanout214 _1472_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout203 net204 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_2
X_2598_ cordic_inst.cordic_inst.y\[13\] _0932_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nor2_1
X_4337_ net140 net191 net155 axi_controller.result_out\[6\] VGND VGND VPWR VPWR _0588_
+ sky130_fd_sc_hd__a22o_1
Xfanout225 net226 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
Xfanout247 _0606_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
Xfanout236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
Xfanout258 net259 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 cordic_inst.cordic_inst.z\[31\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__buf_2
X_4268_ cordic_inst.cordic_inst.cos_out\[28\] cordic_inst.cordic_inst.cos_out\[27\]
+ _2210_ net223 cordic_inst.cordic_inst.cos_out\[29\] VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__o311a_1
X_3219_ cordic_inst.cordic_inst.y\[14\] cordic_inst.cordic_inst.sin_out\[14\] net212
+ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
X_4199_ _2162_ _2165_ axi_controller.result_out\[20\] net205 VGND VGND VPWR VPWR _0374_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3570_ cordic_inst.cordic_inst.x\[9\] cordic_inst.cordic_inst.cos_out\[9\] net210
+ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521_ _0782_ _0785_ net251 VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a21o_1
X_2452_ _0782_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nand2_1
X_2383_ net247 _0699_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4122_ _2094_ _2095_ _2097_ net314 VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__o22ai_1
X_4053_ _2035_ _2037_ net230 VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__mux2_1
XFILLER_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3004_ cordic_inst.cordic_inst.x\[13\] _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__or2_1
Xinput3 araddr[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4955_ net402 _0584_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3906_ axi_controller.read_addr_reg\[7\] net31 net198 VGND VGND VPWR VPWR _0273_
+ sky130_fd_sc_hd__mux2_1
X_4886_ net357 axi_controller.reg_input_data\[18\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_3837_ net35 _1922_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__nor2_1
X_3768_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1871_
+ _1872_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2719_ _0955_ _1037_ _0962_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o21a_1
X_3699_ cordic_inst.deg_handler_inst.theta_norm\[8\] cordic_inst.deg_handler_inst.theta_norm\[7\]
+ _1824_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ net391 _0467_ _0162_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4671_ net375 cordic_inst.cordic_inst.next_state\[0\] _0093_ VGND VGND VPWR VPWR
+ cordic_inst.cordic_inst.state\[0\] sky130_fd_sc_hd__dfrtp_1
X_3622_ _1779_ _1783_ _1787_ _1788_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__or4_1
X_3553_ cordic_inst.cordic_inst.x\[26\] cordic_inst.cordic_inst.cos_out\[26\] net207
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux2_1
X_3484_ _1648_ _1705_ _1651_ _1641_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__a211o_1
X_2504_ _0792_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__xnor2_1
X_2435_ net154 _0758_ _0765_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__and4_1
X_4105_ cordic_inst.cordic_inst.sin_out\[9\] net258 _2081_ net228 VGND VGND VPWR VPWR
+ _2083_ sky130_fd_sc_hd__a31o_1
X_2366_ cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.x\[13\] cordic_inst.cordic_inst.x\[14\]
+ cordic_inst.cordic_inst.x\[15\] net309 net297 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux4_1
X_2297_ cordic_inst.cordic_inst.x\[30\] net265 net304 VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux2_1
X_4036_ net98 _2019_ _2025_ net350 VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o211a_1
XFILLER_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4938_ net384 _0567_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_1
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4869_ net368 axi_controller.reg_input_data\[1\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2984_ cordic_inst.cordic_inst.x\[8\] _1286_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4723_ net374 _0450_ _0145_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[16\] sky130_fd_sc_hd__dfrtp_1
X_4654_ net382 _0385_ net325 VGND VGND VPWR VPWR axi_controller.result_out\[31\] sky130_fd_sc_hd__dfrtp_1
Xinput50 awaddr[22] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 awaddr[3] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
X_4585_ net380 _0317_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[18\] sky130_fd_sc_hd__dfxtp_1
Xinput72 wdata[10] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
X_3605_ cordic_inst.deg_handler_inst.theta_abs\[16\] _1772_ VGND VGND VPWR VPWR _1773_
+ sky130_fd_sc_hd__or2_1
Xinput94 wdata[30] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xinput83 wdata[20] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
X_3536_ _1592_ _1594_ _1601_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__and3_1
X_3467_ _1493_ _1692_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__nand2_1
X_3398_ cordic_inst.cordic_inst.z\[19\] _1636_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__or2_1
X_2418_ net285 _0751_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a21o_1
X_2349_ net277 _0651_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a21o_1
X_4019_ axi_controller.reg_input_data\[30\] _2008_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__or2_1
XFILLER_38_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4370_ net337 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
X_3321_ net266 _1504_ _1559_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__mux2_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3252_ net248 cordic_inst.cordic_inst.z\[22\] VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__and2_1
X_3183_ _1249_ _1281_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2967_ _0603_ _1138_ _1147_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__and3_1
X_2898_ net246 _1137_ net215 VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__a21oi_4
X_4706_ net379 _0433_ _0128_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_4637_ net406 _0368_ net342 VGND VGND VPWR VPWR axi_controller.result_out\[14\] sky130_fd_sc_hd__dfrtp_1
X_4568_ net364 _0300_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_3519_ cordic_inst.cordic_inst.angle\[9\] net171 net160 cordic_inst.cordic_inst.z\[9\]
+ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__a22o_1
X_4499_ net341 VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__inv_2
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3870_ _1948_ _1950_ _1951_ _1952_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_42_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2821_ net283 _1119_ _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a21o_1
X_2752_ _0910_ _0912_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__xor2_1
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4422_ net329 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__inv_2
X_2683_ _0984_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__xnor2_1
X_4353_ net323 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
X_3304_ _1481_ net266 _1542_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__mux2_1
Xfanout407 net408 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_2
X_4284_ cordic_inst.cordic_inst.sin_out\[31\] _2238_ _2239_ VGND VGND VPWR VPWR _2240_
+ sky130_fd_sc_hd__o21ai_1
X_3235_ net268 cordic_inst.cordic_inst.z\[30\] VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__xnor2_1
X_3166_ cordic_inst.cordic_inst.x\[13\] net168 _1450_ net185 VGND VGND VPWR VPWR _0511_
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3097_ cordic_inst.cordic_inst.x\[27\] _1384_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_40_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3999_ net108 _0610_ _1924_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3020_ _1321_ _1322_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nand2_1
XFILLER_17_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3922_ axi_controller.read_addr_reg\[23\] net17 net197 VGND VGND VPWR VPWR _0289_
+ sky130_fd_sc_hd__mux2_1
X_3853_ net44 net43 net46 net45 VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__or4_1
XFILLER_32_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2804_ cordic_inst.cordic_inst.y\[10\] cordic_inst.cordic_inst.y\[11\] cordic_inst.cordic_inst.y\[12\]
+ cordic_inst.cordic_inst.y\[13\] net308 net297 VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__mux4_1
X_3784_ axi_controller.reg_input_data\[21\] _1886_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__nand2_1
X_2735_ _0945_ _1039_ _0942_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__o21ai_1
X_2666_ _0639_ _0806_ _0807_ net269 VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__o31a_1
X_4405_ net320 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__inv_2
X_4336_ net141 net191 net155 axi_controller.result_out\[7\] VGND VGND VPWR VPWR _0587_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout204 net205 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_4
X_2597_ _0778_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__xnor2_1
Xfanout237 _0608_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_2
Xfanout215 _1068_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net227 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_4
Xfanout248 net249 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_2
Xfanout259 cordic_inst.deg_handler_inst.isNegative VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
X_4267_ cordic_inst.cordic_inst.sin_out\[29\] net256 _2221_ VGND VGND VPWR VPWR _2225_
+ sky130_fd_sc_hd__nand3_1
X_4198_ net314 _2164_ net205 VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__o21a_1
X_3218_ cordic_inst.cordic_inst.y\[15\] cordic_inst.cordic_inst.sin_out\[15\] net213
+ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_1
X_3149_ cordic_inst.cordic_inst.x\[17\] net166 _1437_ net184 VGND VGND VPWR VPWR _0515_
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2520_ net251 _0782_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__or2_1
XFILLER_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2451_ _0783_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and2_1
X_2382_ net284 _0702_ _0715_ _0716_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__a211o_1
X_4121_ cordic_inst.cordic_inst.cos_out\[11\] _2096_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__xnor2_1
X_4052_ cordic_inst.cordic_inst.cos_out\[2\] _2036_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__xor2_1
Xinput4 araddr[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_3003_ _1192_ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4954_ net402 _0583_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_1
X_3905_ axi_controller.read_addr_reg\[6\] net30 net198 VGND VGND VPWR VPWR _0272_
+ sky130_fd_sc_hd__mux2_1
X_4885_ net357 axi_controller.reg_input_data\[17\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_3836_ net68 net35 VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__nor2_1
X_3767_ axi_controller.reg_input_data\[30\] axi_controller.reg_input_data\[29\] axi_controller.reg_input_data\[28\]
+ axi_controller.reg_input_data\[27\] VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ _0915_ _0959_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__or2_1
X_3698_ cordic_inst.deg_handler_inst.theta_norm\[8\] _1826_ VGND VGND VPWR VPWR _0038_
+ sky130_fd_sc_hd__xnor2_1
X_2649_ _0982_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__and2b_1
X_4319_ net128 net193 net157 axi_controller.result_out\[24\] VGND VGND VPWR VPWR _0570_
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4670_ net371 _0399_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
X_3621_ _0615_ cordic_inst.deg_handler_inst.theta_abs\[19\] cordic_inst.deg_handler_inst.theta_abs\[22\]
+ cordic_inst.deg_handler_inst.theta_abs\[23\] VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__or4b_1
X_3552_ cordic_inst.cordic_inst.x\[27\] cordic_inst.cordic_inst.cos_out\[27\] net207
+ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
X_2503_ _0789_ _0793_ net271 VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__o21a_1
X_3483_ cordic_inst.cordic_inst.angle\[19\] net173 net162 cordic_inst.cordic_inst.z\[19\]
+ _1709_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a221o_1
X_2434_ net278 _0766_ _0767_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a22o_1
X_2365_ cordic_inst.cordic_inst.x\[8\] cordic_inst.cordic_inst.x\[9\] cordic_inst.cordic_inst.x\[10\]
+ cordic_inst.cordic_inst.x\[11\] net309 net298 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__mux4_1
X_4104_ net258 _2081_ cordic_inst.cordic_inst.sin_out\[9\] VGND VGND VPWR VPWR _2082_
+ sky130_fd_sc_hd__a21oi_1
X_2296_ net264 net278 VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nand2_1
X_4035_ axi_controller.reg_input_data\[5\] _2018_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__or2_1
XFILLER_37_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4937_ net385 _0566_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_1
X_4868_ net368 axi_controller.reg_input_data\[0\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3819_ _1912_ _1910_ axi_controller.reg_input_data\[29\] VGND VGND VPWR VPWR _1913_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4799_ net386 _0526_ _0221_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[28\] sky130_fd_sc_hd__dfrtp_2
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2983_ _1184_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__xor2_1
XFILLER_21_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4722_ net360 _0449_ _0144_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[15\] sky130_fd_sc_hd__dfrtp_1
Xinput40 awaddr[13] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
X_4653_ net381 _0384_ net317 VGND VGND VPWR VPWR axi_controller.result_out\[30\] sky130_fd_sc_hd__dfrtp_1
Xinput51 awaddr[23] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 awaddr[4] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_1
X_4584_ net370 _0316_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[17\] sky130_fd_sc_hd__dfxtp_1
Xinput73 wdata[11] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
X_3604_ cordic_inst.deg_handler_inst.theta_abs\[15\] _1771_ VGND VGND VPWR VPWR _1772_
+ sky130_fd_sc_hd__or2_1
Xinput84 wdata[21] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 wdata[31] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
X_3535_ net182 _1605_ _1745_ _1746_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a31o_1
X_3466_ net180 _1694_ _1695_ _1696_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a31o_1
X_2417_ net218 _0726_ _0730_ net221 net277 VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a221o_1
X_3397_ net267 _1635_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__xnor2_1
X_2348_ net284 _0669_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__a21oi_1
X_2279_ cordic_inst.deg_handler_inst.theta_abs\[18\] VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__inv_2
X_4018_ net92 _2009_ _2015_ net346 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o211a_1
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3320_ net220 _1557_ _1558_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__or3_1
X_3251_ _1488_ _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__nand2_1
X_3182_ _1459_ _1460_ cordic_inst.cordic_inst.x\[7\] net168 VGND VGND VPWR VPWR _0505_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2966_ cordic_inst.cordic_inst.x\[1\] _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__nand2_1
X_2897_ _1069_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nand2_1
X_4705_ net379 _0432_ _0127_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_4636_ net406 _0367_ net342 VGND VGND VPWR VPWR axi_controller.result_out\[13\] sky130_fd_sc_hd__dfrtp_1
X_4567_ net364 _0299_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_3518_ _1616_ _1619_ _1622_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__o21ai_1
X_4498_ net341 VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__inv_2
X_3449_ net180 _1682_ _1683_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2820_ net221 _1121_ _1122_ net218 net275 VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__a221o_1
X_2751_ net185 _1057_ _1060_ net168 cordic_inst.cordic_inst.y\[6\] VGND VGND VPWR
+ VPWR _0536_ sky130_fd_sc_hd__a32o_1
X_2682_ cordic_inst.cordic_inst.y\[26\] _0985_ _1012_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a21oi_1
X_4421_ net322 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__inv_2
X_4352_ net323 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
Xfanout408 net1 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_4
X_3303_ net222 _0706_ _0712_ _1541_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__and4b_1
X_4283_ cordic_inst.cordic_inst.sin_out\[31\] _2238_ net231 VGND VGND VPWR VPWR _2239_
+ sky130_fd_sc_hd__a21oi_1
X_3234_ net249 cordic_inst.cordic_inst.z\[30\] VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__nand2_1
X_3165_ _1309_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3096_ cordic_inst.cordic_inst.x\[27\] _1384_ _1387_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__o21ba_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3998_ _0611_ _2002_ _2004_ _0621_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a211oi_1
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2949_ _0602_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__and2_1
XFILLER_13_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4619_ net363 _0350_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3921_ axi_controller.read_addr_reg\[22\] net16 net196 VGND VGND VPWR VPWR _0288_
+ sky130_fd_sc_hd__mux2_1
X_3852_ net49 net48 net51 net50 VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__or4_1
X_2803_ _1104_ _1105_ net290 VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux2_1
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3783_ axi_controller.reg_input_data\[20\] axi_controller.reg_input_data\[19\] _1874_
+ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__o21ba_1
X_2734_ net184 _1041_ _1049_ net166 cordic_inst.cordic_inst.y\[12\] VGND VGND VPWR
+ VPWR _0542_ sky130_fd_sc_hd__a32o_1
X_2665_ _0819_ _0997_ _0812_ _0815_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__a211o_1
X_4404_ net320 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__inv_2
X_2596_ _0770_ _0773_ net250 VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a21o_1
Xfanout205 cordic_inst.sign_handler_inst.done_pulse VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4335_ net142 net191 net155 axi_controller.result_out\[8\] VGND VGND VPWR VPWR _0586_
+ sky130_fd_sc_hd__a22o_1
Xfanout227 _0613_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_4
Xfanout238 net239 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_2
Xfanout249 _0604_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_2
X_4266_ net256 _2221_ cordic_inst.cordic_inst.sin_out\[29\] VGND VGND VPWR VPWR _2224_
+ sky130_fd_sc_hd__a21o_1
X_4197_ cordic_inst.cordic_inst.cos_out\[20\] _2163_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__xnor2_1
X_3217_ cordic_inst.cordic_inst.y\[16\] cordic_inst.cordic_inst.sin_out\[16\] net213
+ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
X_3148_ _1367_ _1436_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ _1377_ _1381_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__nand2_1
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2450_ net245 _0699_ net170 VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a21oi_1
X_2381_ cordic_inst.cordic_inst.x\[0\] net222 _0711_ _0704_ net219 VGND VGND VPWR
+ VPWR _0716_ sky130_fd_sc_hd__a32o_1
X_4120_ cordic_inst.cordic_inst.cos_out\[10\] _2089_ net225 VGND VGND VPWR VPWR _2096_
+ sky130_fd_sc_hd__o21a_1
X_4051_ cordic_inst.cordic_inst.cos_out\[1\] cordic_inst.cordic_inst.cos_out\[0\]
+ net224 VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__o21a_1
X_3002_ _1189_ _1190_ net272 VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__o21a_1
Xinput5 araddr[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4953_ net402 _0582_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_1
X_3904_ axi_controller.read_addr_reg\[5\] net29 net198 VGND VGND VPWR VPWR _0271_
+ sky130_fd_sc_hd__mux2_1
X_4884_ net357 axi_controller.reg_input_data\[16\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3835_ _0610_ net68 VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__or2_1
X_3766_ axi_controller.reg_input_data\[22\] _1870_ axi_controller.reg_input_data\[23\]
+ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__o21a_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2717_ net184 _0972_ _1036_ net167 cordic_inst.cordic_inst.y\[16\] VGND VGND VPWR
+ VPWR _0546_ sky130_fd_sc_hd__a32o_1
X_3697_ cordic_inst.deg_handler_inst.theta_norm\[7\] _1824_ net252 VGND VGND VPWR
+ VPWR _1826_ sky130_fd_sc_hd__o21ai_1
X_2648_ cordic_inst.cordic_inst.y\[27\] _0981_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__nand2_1
X_2579_ cordic_inst.cordic_inst.y\[7\] _0872_ _0879_ _0913_ _0877_ VGND VGND VPWR
+ VPWR _0914_ sky130_fd_sc_hd__o221a_1
X_4318_ net129 net193 net157 axi_controller.result_out\[25\] VGND VGND VPWR VPWR _0569_
+ sky130_fd_sc_hd__a22o_1
X_4249_ axi_controller.result_out\[26\] _2209_ net201 VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3620_ cordic_inst.deg_handler_inst.theta_abs\[17\] _1773_ VGND VGND VPWR VPWR _1787_
+ sky130_fd_sc_hd__or2_2
X_3551_ cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.cos_out\[28\] net207
+ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
X_2502_ _0835_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nand2_1
X_3482_ _1639_ _1707_ _1708_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__o21a_1
X_2433_ net240 _0739_ net277 VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__a21oi_1
X_2364_ _0696_ _0698_ net285 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__mux2_1
X_4103_ cordic_inst.cordic_inst.sin_out\[8\] _2075_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__or2_1
X_2295_ _0601_ net244 VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__nor2_1
X_4034_ net97 _2019_ _2024_ net350 VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_35_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4936_ net385 _0565_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4867_ net376 _0077_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3818_ _1911_ _1912_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4798_ net386 _0525_ _0220_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[27\] sky130_fd_sc_hd__dfrtp_4
XFILLER_4_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3749_ cordic_inst.deg_handler_inst.theta_norm\[27\] _1858_ VGND VGND VPWR VPWR _0027_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2982_ net272 _1180_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4721_ net360 _0448_ _0143_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4652_ net385 _0383_ net325 VGND VGND VPWR VPWR axi_controller.result_out\[29\] sky130_fd_sc_hd__dfrtp_1
X_3603_ cordic_inst.deg_handler_inst.theta_abs\[14\] _1770_ VGND VGND VPWR VPWR _1771_
+ sky130_fd_sc_hd__or2_1
Xinput30 araddr[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput52 awaddr[24] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 awaddr[5] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
X_4583_ net380 _0315_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[16\] sky130_fd_sc_hd__dfxtp_1
Xinput41 awaddr[14] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput96 wdata[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput85 wdata[22] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_1
Xinput74 wdata[12] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
X_3534_ cordic_inst.cordic_inst.angle\[4\] net171 net160 cordic_inst.cordic_inst.z\[4\]
+ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__a22o_1
X_3465_ cordic_inst.cordic_inst.angle\[23\] net173 net161 cordic_inst.cordic_inst.z\[23\]
+ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__a22o_1
X_2416_ _0719_ _0727_ net235 VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__mux2_1
X_3396_ net280 _1576_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__nor2_1
X_2347_ net221 _0679_ net219 _0681_ net277 VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a221o_1
X_2278_ cordic_inst.cordic_inst.state\[1\] VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__inv_2
X_4017_ axi_controller.reg_input_data\[29\] _2008_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__or2_1
XFILLER_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4919_ net358 _0018_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3250_ cordic_inst.cordic_inst.z\[20\] _1487_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__or2_1
X_3181_ _1247_ _1282_ _1283_ net177 VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__a31o_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2965_ _1157_ _1267_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__xnor2_1
X_4704_ net386 _0431_ _0126_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_2896_ net244 _1151_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__nand2_1
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4635_ net401 _0366_ net338 VGND VGND VPWR VPWR axi_controller.result_out\[12\] sky130_fd_sc_hd__dfrtp_1
X_4566_ net370 _0298_ VGND VGND VPWR VPWR axi_controller.reg_done_flag sky130_fd_sc_hd__dfxtp_1
X_3517_ _1616_ _1619_ _1622_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__or3_1
X_4497_ net341 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_2
X_3448_ cordic_inst.cordic_inst.angle\[27\] net173 net161 cordic_inst.cordic_inst.z\[27\]
+ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__a22o_1
X_3379_ _1616_ _1617_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ _0877_ _0878_ _0913_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__a21o_1
XFILLER_8_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2681_ _0986_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__and2_1
X_4420_ net322 VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__inv_2
X_4351_ net321 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
X_3302_ net280 net288 VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__nand2_1
X_4282_ cordic_inst.cordic_inst.sin_out\[30\] _2224_ net256 VGND VGND VPWR VPWR _2238_
+ sky130_fd_sc_hd__o21a_1
X_3233_ cordic_inst.cordic_inst.y\[0\] cordic_inst.cordic_inst.sin_out\[0\] net208
+ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3164_ cordic_inst.cordic_inst.x\[12\] _1310_ _1443_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3095_ _1394_ _1397_ _1385_ _1389_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__and4bb_1
XFILLER_35_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3997_ _1961_ _1995_ _2003_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__a21oi_1
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2948_ _1131_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_20_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2879_ net262 _1149_ _1150_ _1152_ net243 net240 VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__mux4_1
X_4618_ net363 _0349_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4549_ net355 _0281_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3920_ axi_controller.read_addr_reg\[21\] net15 net196 VGND VGND VPWR VPWR _0287_
+ sky130_fd_sc_hd__mux2_1
X_3851_ net66 net38 net37 net40 VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__or4_1
X_3782_ _1880_ _1883_ axi_controller.reg_input_data\[21\] VGND VGND VPWR VPWR _1885_
+ sky130_fd_sc_hd__o21a_1
X_2802_ cordic_inst.cordic_inst.y\[18\] cordic_inst.cordic_inst.y\[19\] cordic_inst.cordic_inst.y\[20\]
+ cordic_inst.cordic_inst.y\[21\] net311 net300 VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__mux4_1
XFILLER_9_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2733_ _0930_ _1040_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__or2_1
XFILLER_8_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2664_ _0819_ _0997_ _0815_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a21o_1
X_4403_ net320 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__inv_2
X_2595_ _0928_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nor2_1
X_4334_ net143 net192 net155 axi_controller.result_out\[9\] VGND VGND VPWR VPWR _0585_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout228 net229 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_2
X_4265_ axi_controller.result_out\[28\] _2223_ net200 VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
Xfanout239 _0607_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_4
X_4196_ cordic_inst.cordic_inst.cos_out\[19\] _2155_ net227 VGND VGND VPWR VPWR _2163_
+ sky130_fd_sc_hd__o21a_1
X_3216_ cordic_inst.cordic_inst.y\[17\] cordic_inst.cordic_inst.sin_out\[17\] net212
+ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3147_ cordic_inst.cordic_inst.x\[16\] _1360_ _1361_ _1332_ VGND VGND VPWR VPWR _1436_
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3078_ _1379_ _1380_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__nor2_1
XFILLER_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2380_ cordic_inst.cordic_inst.x\[1\] net217 net216 _0710_ net276 VGND VGND VPWR
+ VPWR _0715_ sky130_fd_sc_hd__a221o_1
X_4050_ cordic_inst.cordic_inst.sin_out\[2\] _2034_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__xnor2_1
Xinput6 araddr[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_3001_ _1299_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__and2_1
XFILLER_36_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4952_ net407 _0581_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4883_ net357 axi_controller.reg_input_data\[15\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3903_ axi_controller.read_addr_reg\[4\] net28 net198 VGND VGND VPWR VPWR _0270_
+ sky130_fd_sc_hd__mux2_1
X_3834_ net111 axi_controller.state\[2\] net69 _0621_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__a31o_1
X_3765_ axi_controller.reg_input_data\[19\] _1869_ axi_controller.reg_input_data\[21\]
+ axi_controller.reg_input_data\[20\] VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3696_ cordic_inst.deg_handler_inst.theta_norm\[7\] _1825_ VGND VGND VPWR VPWR _0037_
+ sky130_fd_sc_hd__xnor2_1
X_2716_ _0968_ _0970_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__nand2_1
X_2647_ cordic_inst.cordic_inst.y\[27\] _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nor2_1
XFILLER_10_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2578_ _0906_ _0907_ _0912_ _0911_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__a31o_1
X_4317_ net130 net194 net157 axi_controller.result_out\[26\] VGND VGND VPWR VPWR _0568_
+ sky130_fd_sc_hd__a22o_1
X_4248_ net313 _2208_ _2206_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__a21o_1
XFILLER_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4179_ net226 _2147_ cordic_inst.cordic_inst.cos_out\[18\] VGND VGND VPWR VPWR _2148_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3550_ cordic_inst.cordic_inst.x\[29\] cordic_inst.cordic_inst.cos_out\[29\] net207
+ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
X_2501_ cordic_inst.cordic_inst.y\[20\] _0834_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__or2_1
XFILLER_6_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3481_ _1639_ _1707_ net175 VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__a21oi_1
X_2432_ net287 _0661_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2363_ _0641_ _0697_ net234 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__mux2_1
X_4102_ cordic_inst.cordic_inst.cos_out\[9\] _2079_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__xor2_1
X_2294_ net162 VGND VGND VPWR VPWR cordic_inst.cordic_inst.next_state\[1\] sky130_fd_sc_hd__inv_2
X_4033_ axi_controller.reg_input_data\[4\] _2018_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__or2_1
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4935_ net382 _0564_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_1
X_4866_ net376 _0076_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[30\] sky130_fd_sc_hd__dfxtp_1
X_3817_ axi_controller.reg_input_data\[28\] axi_controller.reg_input_data\[27\] _1908_
+ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__nor3_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4797_ net386 _0524_ _0219_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[26\] sky130_fd_sc_hd__dfrtp_2
X_3748_ net254 _1857_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__nand2_1
XFILLER_20_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3679_ cordic_inst.deg_handler_inst.theta_abs\[30\] net152 VGND VGND VPWR VPWR _0076_
+ sky130_fd_sc_hd__and2_1
Xoutput140 net140 VGND VGND VPWR VPWR rdata[6] sky130_fd_sc_hd__buf_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2981_ _1244_ _1247_ _1282_ _1243_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__a31o_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4720_ net360 _0447_ _0142_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4651_ net385 _0382_ net325 VGND VGND VPWR VPWR axi_controller.result_out\[28\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_26_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3602_ cordic_inst.deg_handler_inst.theta_abs\[13\] _1769_ VGND VGND VPWR VPWR _1770_
+ sky130_fd_sc_hd__or2_1
Xinput20 araddr[26] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 araddr[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput53 awaddr[25] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 awaddr[6] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
X_4582_ net369 _0314_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[15\] sky130_fd_sc_hd__dfxtp_1
Xinput42 awaddr[15] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_1
Xinput97 wdata[4] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
Xinput86 wdata[23] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
Xinput75 wdata[13] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
X_3533_ _1591_ _1602_ _1604_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_10_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3464_ _1491_ _1494_ _1693_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__or3_1
X_2415_ _0746_ _0749_ net277 VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__mux2_1
X_3395_ _1632_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__nor2_1
X_2346_ cordic_inst.cordic_inst.x\[11\] cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.x\[13\]
+ cordic_inst.cordic_inst.x\[14\] net309 net298 VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux4_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2277_ cordic_inst.deg_handler_inst.kuadran\[0\] VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__inv_2
X_4016_ net91 _2009_ _2014_ net348 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o211a_1
XFILLER_38_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4918_ net358 _0017_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_4849_ net359 _0057_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcordic_system_410 VGND VGND VPWR VPWR cordic_system_410/HI rresp[0] sky130_fd_sc_hd__conb_1
X_3180_ _1247_ _1282_ _1283_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2964_ net270 _1138_ _1147_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__and3_1
XFILLER_22_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4703_ net386 _0430_ _0125_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_2895_ net244 _1196_ _1197_ net215 VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a31o_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4634_ net401 _0365_ net338 VGND VGND VPWR VPWR axi_controller.result_out\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4565_ net355 _0297_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[31\] sky130_fd_sc_hd__dfxtp_1
X_3516_ cordic_inst.cordic_inst.angle\[10\] net171 net159 cordic_inst.cordic_inst.z\[10\]
+ _1733_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4496_ net337 VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__inv_2
X_3447_ _1660_ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__xnor2_1
X_3378_ cordic_inst.cordic_inst.z\[8\] _1615_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__nor2_1
X_2329_ net285 _0661_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_4_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2680_ _0979_ _0993_ _0989_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__o21a_1
X_4350_ net321 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
X_3301_ _1538_ _1539_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__nand2_1
XFILLER_4_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4281_ cordic_inst.cordic_inst.cos_out\[30\] _2227_ net223 cordic_inst.cordic_inst.cos_out\[31\]
+ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__o211a_1
X_3232_ cordic_inst.cordic_inst.y\[1\] cordic_inst.cordic_inst.sin_out\[1\] net214
+ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
X_3163_ net185 _1445_ _1448_ net168 cordic_inst.cordic_inst.x\[14\] VGND VGND VPWR
+ VPWR _0512_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_1_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3094_ _1379_ _1393_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__nor2_1
XFILLER_23_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3996_ _0624_ _1942_ _1998_ _2002_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__a31o_1
XFILLER_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947_ net251 _1178_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2878_ net241 _1150_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__nand2_1
X_4617_ net368 _0348_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_4548_ net355 _0280_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[14\] sky130_fd_sc_hd__dfxtp_1
X_4479_ net327 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_13_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3850_ net58 net65 net64 net67 VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__or4_1
X_3781_ axi_controller.reg_input_data\[21\] _1880_ _1883_ VGND VGND VPWR VPWR _1884_
+ sky130_fd_sc_hd__nor3_1
XFILLER_20_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2801_ cordic_inst.cordic_inst.y\[14\] cordic_inst.cordic_inst.y\[15\] cordic_inst.cordic_inst.y\[16\]
+ cordic_inst.cordic_inst.y\[17\] net310 net299 VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__mux4_1
XFILLER_13_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2732_ cordic_inst.cordic_inst.y\[13\] net166 _1048_ net184 VGND VGND VPWR VPWR _0543_
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2663_ _0815_ _0818_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__and2b_1
X_4402_ net320 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__inv_2
X_2594_ cordic_inst.cordic_inst.y\[12\] _0927_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__and2b_1
X_4333_ net113 net191 net155 axi_controller.result_out\[10\] VGND VGND VPWR VPWR _0584_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout218 net219 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_2
Xfanout229 net230 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
X_4264_ net313 _2219_ _2222_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__o21ai_1
Xfanout207 net209 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_4
X_3215_ cordic_inst.cordic_inst.y\[18\] cordic_inst.cordic_inst.sin_out\[18\] net212
+ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
X_4195_ cordic_inst.cordic_inst.sin_out\[20\] net261 _2159_ _2161_ VGND VGND VPWR
+ VPWR _2162_ sky130_fd_sc_hd__a31o_1
X_3146_ net185 _1432_ _1435_ net167 cordic_inst.cordic_inst.x\[18\] VGND VGND VPWR
+ VPWR _0516_ sky130_fd_sc_hd__a32o_1
XFILLER_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3077_ cordic_inst.cordic_inst.x\[24\] _1378_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__nor2_1
XFILLER_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3979_ axi_controller.write_addr_reg\[28\] net56 net189 VGND VGND VPWR VPWR _0327_
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 araddr[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_3000_ cordic_inst.cordic_inst.x\[14\] _1301_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__xor2_1
XFILLER_45_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4951_ net406 _0580_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_1
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4882_ net356 axi_controller.reg_input_data\[14\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3902_ axi_controller.read_addr_reg\[3\] net27 net197 VGND VGND VPWR VPWR _0269_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3833_ net111 net69 VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__nand2_1
X_3764_ axi_controller.reg_input_data\[17\] axi_controller.reg_input_data\[16\] _1868_
+ axi_controller.reg_input_data\[18\] VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_30_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3695_ net252 _1824_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__nand2_1
X_2715_ cordic_inst.cordic_inst.y\[17\] net166 _1035_ net184 VGND VGND VPWR VPWR _0547_
+ sky130_fd_sc_hd__a22o_1
X_2646_ _0804_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__xnor2_1
X_2577_ _0883_ _0885_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__nor2_1
X_4316_ net131 net194 net157 axi_controller.result_out\[27\] VGND VGND VPWR VPWR _0567_
+ sky130_fd_sc_hd__a22o_1
X_4247_ cordic_inst.cordic_inst.sin_out\[26\] _2207_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_40_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4178_ cordic_inst.cordic_inst.cos_out\[17\] cordic_inst.cordic_inst.cos_out\[16\]
+ _2132_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__or3_1
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3129_ _1337_ _1423_ _1335_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3480_ cordic_inst.cordic_inst.z\[18\] _1640_ _1706_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__a21o_1
X_2500_ cordic_inst.cordic_inst.y\[20\] _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__nand2_1
X_2431_ net286 _0662_ _0637_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__o21a_1
X_2362_ cordic_inst.cordic_inst.x\[24\] cordic_inst.cordic_inst.x\[25\] cordic_inst.cordic_inst.x\[26\]
+ cordic_inst.cordic_inst.x\[27\] net305 net295 VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux4_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2293_ net181 net174 VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__nor2_2
X_4101_ cordic_inst.cordic_inst.cos_out\[8\] cordic_inst.cordic_inst.cos_out\[7\]
+ _2068_ net225 VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__o31a_1
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4032_ net96 _2019_ _2023_ net350 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__o211a_1
XFILLER_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4934_ net385 _0563_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4865_ net389 _0074_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[29\] sky130_fd_sc_hd__dfxtp_1
X_3816_ axi_controller.reg_input_data\[29\] _1910_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__xnor2_1
X_4796_ net386 _0523_ _0218_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[25\] sky130_fd_sc_hd__dfrtp_2
X_3747_ cordic_inst.deg_handler_inst.theta_norm\[26\] cordic_inst.deg_handler_inst.theta_norm\[25\]
+ _1854_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__or3_1
X_3678_ cordic_inst.deg_handler_inst.theta_abs\[29\] net153 VGND VGND VPWR VPWR _0074_
+ sky130_fd_sc_hd__and2_1
Xoutput130 net130 VGND VGND VPWR VPWR rdata[26] sky130_fd_sc_hd__buf_2
Xoutput141 net141 VGND VGND VPWR VPWR rdata[7] sky130_fd_sc_hd__buf_2
X_2629_ _0939_ _0963_ _0962_ _0948_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout390 net391 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2980_ _1243_ _1244_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__nand2b_1
X_4650_ net384 _0381_ net325 VGND VGND VPWR VPWR axi_controller.result_out\[27\] sky130_fd_sc_hd__dfrtp_1
Xinput21 araddr[27] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
X_3601_ cordic_inst.deg_handler_inst.theta_abs\[12\] _1768_ VGND VGND VPWR VPWR _1769_
+ sky130_fd_sc_hd__or2_1
Xinput10 araddr[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput43 awaddr[16] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
Xinput54 awaddr[26] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
X_4581_ net363 _0313_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[14\] sky130_fd_sc_hd__dfxtp_1
Xinput32 araddr[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput98 wdata[5] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
Xinput65 awaddr[7] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
Xinput76 wdata[14] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_1
Xinput87 wdata[24] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
X_3532_ cordic_inst.cordic_inst.angle\[5\] net171 net160 cordic_inst.cordic_inst.z\[5\]
+ _1744_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__a221o_1
X_3463_ _1491_ _1693_ _1494_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__o21ai_1
X_2414_ net285 _0747_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__o21ai_2
X_3394_ cordic_inst.cordic_inst.z\[16\] _1631_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__and2b_1
X_2345_ net286 net291 VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__and2b_1
XFILLER_29_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2276_ net318 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
X_4015_ axi_controller.reg_input_data\[28\] _2008_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__or2_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4917_ net357 _0016_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_4848_ net359 _0056_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[12\] sky130_fd_sc_hd__dfxtp_1
X_4779_ net397 _0506_ _0201_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2963_ cordic_inst.cordic_inst.x\[2\] _1265_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__nand2_1
X_4702_ net386 _0429_ _0124_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2894_ net238 _1088_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__or2_1
X_4633_ net401 _0364_ net338 VGND VGND VPWR VPWR axi_controller.result_out\[10\] sky130_fd_sc_hd__dfrtp_1
X_4564_ net351 _0296_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[30\] sky130_fd_sc_hd__dfxtp_1
X_3515_ net175 _1732_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__nor2_1
X_4495_ net338 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__inv_2
X_3446_ net249 cordic_inst.cordic_inst.z\[26\] _1680_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__a21boi_1
X_3377_ cordic_inst.cordic_inst.z\[8\] _1615_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__and2_1
X_2328_ net234 _0649_ _0635_ net238 VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__a211o_1
XFILLER_45_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2259_ cordic_inst.cordic_inst.y\[18\] VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__inv_2
XFILLER_38_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3300_ cordic_inst.cordic_inst.z\[11\] _1537_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__nand2_1
X_4280_ cordic_inst.deg_handler_inst.kuadran\[0\] _2232_ cordic_inst.cordic_inst.cos_out\[31\]
+ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__o21ba_1
X_3231_ cordic_inst.cordic_inst.y\[2\] cordic_inst.cordic_inst.sin_out\[2\] net214
+ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
X_3162_ _1303_ _1444_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3093_ _1382_ _1385_ _1389_ _1395_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__and4b_1
X_3995_ net107 _0624_ _1943_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__o21ai_1
X_2946_ _1247_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__nand2_1
X_2877_ _1170_ _1179_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4616_ net368 _0347_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[1\] sky130_fd_sc_hd__dfxtp_1
X_4547_ net351 _0279_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[13\] sky130_fd_sc_hd__dfxtp_1
X_4478_ net327 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__inv_2
X_3429_ cordic_inst.cordic_inst.z\[29\] cordic_inst.cordic_inst.z\[28\] net249 VGND
+ VGND VPWR VPWR _1668_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3780_ axi_controller.reg_input_data\[20\] axi_controller.reg_input_data\[19\] VGND
+ VGND VPWR VPWR _1883_ sky130_fd_sc_hd__and2_1
X_2800_ net275 _1089_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a21o_1
XFILLER_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2731_ _0935_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4401_ net320 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__inv_2
X_2662_ _0983_ _0992_ _0994_ _0995_ _0821_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a41o_1
X_2593_ _0927_ cordic_inst.cordic_inst.y\[12\] VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__and2b_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4332_ net114 net191 net156 axi_controller.result_out\[11\] VGND VGND VPWR VPWR _0583_
+ sky130_fd_sc_hd__a22o_1
Xfanout208 net209 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_4
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout219 net220 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
X_4263_ net231 _2220_ _2221_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__or3b_1
X_3214_ cordic_inst.cordic_inst.y\[19\] cordic_inst.cordic_inst.sin_out\[19\] net214
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
X_4194_ net316 _2160_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__nand2_1
X_3145_ _1358_ _1431_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__nand2_1
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3076_ cordic_inst.cordic_inst.x\[24\] _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__and2_1
XFILLER_36_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3978_ axi_controller.write_addr_reg\[27\] net55 net189 VGND VGND VPWR VPWR _0326_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2929_ net215 _1227_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__or2_1
XFILLER_19_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 araddr[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4950_ net406 _0579_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3901_ axi_controller.read_addr_reg\[2\] net24 net195 VGND VGND VPWR VPWR _0268_
+ sky130_fd_sc_hd__mux2_1
X_4881_ net356 axi_controller.reg_input_data\[13\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3832_ _0620_ _1919_ _1918_ cordic_inst.state\[0\] VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3763_ _1864_ _1865_ _1866_ _1867_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__or4_1
X_3694_ cordic_inst.deg_handler_inst.theta_norm\[6\] _1822_ VGND VGND VPWR VPWR _1824_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2714_ _0868_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__xor2_1
X_2645_ net170 _0798_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__nor2_1
X_4315_ net132 net194 net157 axi_controller.result_out\[28\] VGND VGND VPWR VPWR _0566_
+ sky130_fd_sc_hd__a22o_1
X_2576_ cordic_inst.cordic_inst.y\[4\] _0884_ _0886_ _0885_ VGND VGND VPWR VPWR _0911_
+ sky130_fd_sc_hd__a31o_1
X_4246_ cordic_inst.cordic_inst.sin_out\[25\] _2199_ net256 VGND VGND VPWR VPWR _2207_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4177_ cordic_inst.cordic_inst.sin_out\[18\] net260 _2143_ _2145_ VGND VGND VPWR
+ VPWR _2146_ sky130_fd_sc_hd__a31o_1
XFILLER_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3128_ _1339_ _1422_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__or2_1
XFILLER_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3059_ cordic_inst.cordic_inst.x\[16\] _1360_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_38_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2430_ _0677_ _0763_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nor2_1
X_2361_ _0694_ _0695_ net292 VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux2_1
X_4100_ axi_controller.result_out\[8\] net202 _2078_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__o21ba_1
X_2292_ _0614_ cordic_inst.cordic_inst.state\[0\] VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__and2_1
X_4031_ axi_controller.reg_input_data\[3\] _2018_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__or2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4933_ net380 axi_controller.done _0257_ VGND VGND VPWR VPWR cordic_inst.done_d sky130_fd_sc_hd__dfrtp_1
X_4864_ net376 _0073_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[28\] sky130_fd_sc_hd__dfxtp_1
X_3815_ _1877_ _1900_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__and2_1
X_4795_ net386 _0522_ _0217_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[24\] sky130_fd_sc_hd__dfrtp_2
X_3746_ cordic_inst.deg_handler_inst.theta_norm\[26\] _1856_ VGND VGND VPWR VPWR _0026_
+ sky130_fd_sc_hd__xnor2_1
X_3677_ cordic_inst.deg_handler_inst.theta_abs\[28\] net152 VGND VGND VPWR VPWR _0073_
+ sky130_fd_sc_hd__and2_1
Xoutput131 net131 VGND VGND VPWR VPWR rdata[27] sky130_fd_sc_hd__buf_2
Xoutput142 net142 VGND VGND VPWR VPWR rdata[8] sky130_fd_sc_hd__buf_2
X_2628_ _0941_ _0945_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__or2_1
Xoutput120 net120 VGND VGND VPWR VPWR rdata[17] sky130_fd_sc_hd__buf_2
X_2559_ _0735_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__xor2_1
X_4229_ net257 _2191_ cordic_inst.cordic_inst.sin_out\[24\] VGND VGND VPWR VPWR _2192_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout391 net408 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_2
Xfanout380 net382 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4580_ net363 _0312_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[13\] sky130_fd_sc_hd__dfxtp_1
Xinput11 araddr[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_3600_ cordic_inst.deg_handler_inst.theta_abs\[11\] _1767_ VGND VGND VPWR VPWR _1768_
+ sky130_fd_sc_hd__or2_1
Xinput22 araddr[28] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput44 awaddr[17] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
Xinput55 awaddr[27] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xinput33 araddr[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
X_3531_ net175 _1606_ _1743_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__nor3_1
Xinput66 awaddr[8] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput77 wdata[15] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
Xinput88 wdata[25] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
Xinput99 wdata[6] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
X_3462_ _1493_ _1692_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__nor2_1
X_3393_ _1631_ cordic_inst.cordic_inst.z\[16\] VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__and2b_1
X_2413_ net234 _0641_ _0635_ net238 VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a211o_1
X_2344_ cordic_inst.cordic_inst.x\[7\] cordic_inst.cordic_inst.x\[8\] cordic_inst.cordic_inst.x\[9\]
+ cordic_inst.cordic_inst.x\[10\] net309 net298 VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux4_1
X_2275_ net315 VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__inv_2
XFILLER_38_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4014_ net90 _2009_ _2013_ net348 VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o211a_1
XFILLER_38_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4916_ net358 _0015_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4847_ net359 _0055_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4778_ net396 _0505_ _0200_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3729_ cordic_inst.deg_handler_inst.theta_norm\[19\] _1844_ net253 VGND VGND VPWR
+ VPWR _1846_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2962_ _1164_ _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4701_ net386 _0428_ _0123_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_4632_ net401 _0363_ net338 VGND VGND VPWR VPWR axi_controller.result_out\[9\] sky130_fd_sc_hd__dfrtp_1
X_2893_ net285 _1099_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__or2_1
X_4563_ net351 _0295_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[29\] sky130_fd_sc_hd__dfxtp_1
X_3514_ _1546_ _1623_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__xor2_1
X_4494_ net338 VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__inv_2
X_3445_ _1663_ _1679_ _1661_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__o21ai_1
X_3376_ net266 _1614_ _1613_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__mux2_1
X_2327_ net234 _0649_ _0635_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__a21oi_1
X_2258_ cordic_inst.cordic_inst.y\[28\] VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__inv_2
XFILLER_26_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3230_ cordic_inst.cordic_inst.y\[3\] cordic_inst.cordic_inst.sin_out\[3\] net214
+ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
X_3161_ cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.next_state\[1\] _1446_
+ _1447_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o22a_1
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3092_ _1393_ _1394_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__nor2_1
X_3994_ _0610_ net145 _0619_ net350 _1928_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a41o_1
X_2945_ cordic_inst.cordic_inst.x\[6\] _1246_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__nand2b_1
X_2876_ _1103_ _1116_ _1131_ _1177_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_20_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4615_ net368 _0346_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[0\] sky130_fd_sc_hd__dfxtp_1
X_4546_ net362 _0278_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[12\] sky130_fd_sc_hd__dfxtp_1
X_4477_ net331 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__inv_2
X_3428_ _1477_ _1666_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__nor2_1
X_3359_ cordic_inst.cordic_inst.z\[1\] _1595_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_28_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2730_ _0928_ _1041_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__and2b_1
X_2661_ _0983_ _0992_ _0994_ _0995_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__and4_1
X_4400_ net320 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
X_2592_ _0772_ _0921_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4331_ net115 net192 net156 axi_controller.result_out\[12\] VGND VGND VPWR VPWR _0582_
+ sky130_fd_sc_hd__a22o_1
Xfanout209 _1472_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__buf_2
X_4262_ net256 _2214_ cordic_inst.cordic_inst.sin_out\[28\] VGND VGND VPWR VPWR _2221_
+ sky130_fd_sc_hd__a21o_1
X_3213_ cordic_inst.cordic_inst.y\[20\] cordic_inst.cordic_inst.sin_out\[20\] net214
+ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_4193_ net261 _2159_ cordic_inst.cordic_inst.sin_out\[20\] VGND VGND VPWR VPWR _2160_
+ sky130_fd_sc_hd__a21o_1
XFILLER_28_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3144_ _1433_ _1434_ cordic_inst.cordic_inst.x\[19\] net167 VGND VGND VPWR VPWR _0517_
+ sky130_fd_sc_hd__a2bb2o_1
X_3075_ _1211_ _1221_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3977_ axi_controller.write_addr_reg\[26\] net54 net189 VGND VGND VPWR VPWR _0325_
+ sky130_fd_sc_hd__mux2_1
X_2928_ cordic_inst.cordic_inst.x\[30\] _1229_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__xor2_1
X_2859_ net263 _1073_ _1078_ _1112_ net232 net237 VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__mux4_2
X_4529_ net353 _0261_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 araddr[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4880_ net356 axi_controller.reg_input_data\[12\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3900_ axi_controller.read_addr_reg\[1\] net13 net197 VGND VGND VPWR VPWR _0267_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3831_ cordic_inst.state\[1\] _1919_ cordic_inst.state\[2\] VGND VGND VPWR VPWR _0007_
+ sky130_fd_sc_hd__a21o_1
X_3762_ axi_controller.reg_input_data\[7\] axi_controller.reg_input_data\[6\] axi_controller.reg_input_data\[5\]
+ axi_controller.reg_input_data\[4\] VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__or4_1
XFILLER_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3693_ cordic_inst.deg_handler_inst.theta_norm\[6\] _1823_ VGND VGND VPWR VPWR _0036_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2713_ _0860_ _0972_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__nand2_1
X_2644_ _0974_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nor2_1
X_2575_ cordic_inst.cordic_inst.y\[4\] _0886_ _0908_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a21o_1
X_4314_ net133 net194 net157 axi_controller.result_out\[29\] VGND VGND VPWR VPWR _0565_
+ sky130_fd_sc_hd__a22o_1
X_4245_ _0605_ cordic_inst.deg_handler_inst.kuadran\[0\] _2203_ _2205_ VGND VGND VPWR
+ VPWR _2206_ sky130_fd_sc_hd__o31a_1
X_4176_ net315 _2144_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__nand2_1
X_3127_ _1369_ _1421_ _1346_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__a21o_1
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3058_ cordic_inst.cordic_inst.x\[16\] _1360_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_38_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2360_ cordic_inst.cordic_inst.x\[20\] cordic_inst.cordic_inst.x\[21\] cordic_inst.cordic_inst.x\[22\]
+ cordic_inst.cordic_inst.x\[23\] net312 net301 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux4_1
XFILLER_2_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2291_ _0614_ cordic_inst.cordic_inst.state\[0\] VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4030_ net93 _2019_ _2022_ net350 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o211a_1
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4932_ net368 _0562_ VGND VGND VPWR VPWR axi_controller.start_pulse_reg sky130_fd_sc_hd__dfxtp_1
X_4863_ net375 _0072_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[27\] sky130_fd_sc_hd__dfxtp_1
X_3814_ axi_controller.reg_input_data\[28\] _1909_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4794_ net392 _0521_ _0216_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[23\] sky130_fd_sc_hd__dfrtp_4
X_3745_ cordic_inst.deg_handler_inst.theta_norm\[25\] _1854_ net254 VGND VGND VPWR
+ VPWR _1856_ sky130_fd_sc_hd__o21ai_1
Xoutput110 net110 VGND VGND VPWR VPWR bresp[1] sky130_fd_sc_hd__buf_2
X_3676_ cordic_inst.deg_handler_inst.theta_abs\[27\] net152 VGND VGND VPWR VPWR _0072_
+ sky130_fd_sc_hd__and2_1
Xoutput132 net132 VGND VGND VPWR VPWR rdata[28] sky130_fd_sc_hd__buf_2
Xoutput143 net143 VGND VGND VPWR VPWR rdata[9] sky130_fd_sc_hd__buf_2
X_2627_ _0953_ _0957_ _0952_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__o21a_1
Xoutput121 net121 VGND VGND VPWR VPWR rdata[18] sky130_fd_sc_hd__buf_2
XFILLER_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2558_ net247 _0699_ _0717_ net272 VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__o211a_1
X_2489_ cordic_inst.cordic_inst.y\[22\] _0822_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__or2_1
X_4228_ cordic_inst.cordic_inst.sin_out\[23\] cordic_inst.cordic_inst.sin_out\[22\]
+ _2176_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__or3_1
XFILLER_28_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4159_ net315 _2129_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__nand2_1
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout381 net382 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_2
Xfanout392 net393 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_2
Xfanout370 net371 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_2
Xinput12 araddr[19] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput45 awaddr[18] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 aresetn VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 araddr[29] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
X_3530_ _1570_ _1575_ _1605_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__and3b_1
Xinput56 awaddr[28] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
Xinput67 awaddr[9] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xinput78 wdata[16] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
Xinput89 wdata[26] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
X_3461_ _1486_ _1691_ _1497_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__o21a_1
X_3392_ _1507_ net266 _1630_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__mux2_1
X_2412_ _0695_ _0697_ net290 VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__mux2_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2343_ net286 net291 VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__nor2_1
X_2274_ net110 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__inv_2
X_4013_ axi_controller.reg_input_data\[27\] _2008_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__or2_1
X_4915_ net359 _0014_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_4846_ net359 _0054_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ net391 _0504_ _0199_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[6\] sky130_fd_sc_hd__dfrtp_4
X_3728_ cordic_inst.deg_handler_inst.theta_norm\[19\] _1845_ VGND VGND VPWR VPWR _0018_
+ sky130_fd_sc_hd__xnor2_1
X_3659_ cordic_inst.deg_handler_inst.theta_abs\[18\] net152 net149 _1807_ VGND VGND
+ VPWR VPWR _0062_ sky130_fd_sc_hd__a22o_1
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2961_ _1148_ _1157_ net270 VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__o21a_1
XFILLER_34_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4700_ net384 _0427_ _0122_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_4631_ net398 _0362_ net336 VGND VGND VPWR VPWR axi_controller.result_out\[8\] sky130_fd_sc_hd__dfrtp_1
X_2892_ _1170_ _1179_ _1188_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__or4_2
XFILLER_7_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4562_ net362 _0294_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[28\] sky130_fd_sc_hd__dfxtp_1
X_4493_ net335 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__inv_2
X_3513_ cordic_inst.cordic_inst.angle\[11\] net171 net159 cordic_inst.cordic_inst.z\[11\]
+ _1731_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a221o_1
X_3444_ _1658_ _1659_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__nor2_1
X_3375_ net266 _0712_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__nand2_1
X_2326_ _0646_ _0660_ net236 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux2_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4829_ net393 _0556_ _0251_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3160_ _1299_ _1302_ _1445_ net177 VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__a31o_1
X_3091_ cordic_inst.cordic_inst.x\[25\] _1392_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3993_ net350 _2001_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and2_1
X_2944_ _1246_ cordic_inst.cordic_inst.x\[6\] VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__nand2b_2
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2875_ _1170_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_20_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4614_ net381 _0005_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.kuadran\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4545_ net354 _0277_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[11\] sky130_fd_sc_hd__dfxtp_1
X_4476_ net331 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__inv_2
X_3427_ _1658_ _1659_ _1662_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3358_ _1583_ _1584_ cordic_inst.cordic_inst.z\[0\] VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2309_ net242 _0643_ net170 VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__a21o_1
XFILLER_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3289_ _1520_ _1527_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2660_ _0982_ _0985_ cordic_inst.cordic_inst.y\[26\] VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__nand3b_1
X_2591_ _0920_ _0925_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__or2_1
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4330_ net116 net192 net156 axi_controller.result_out\[13\] VGND VGND VPWR VPWR _0581_
+ sky130_fd_sc_hd__a22o_1
X_4261_ cordic_inst.cordic_inst.sin_out\[28\] net256 _2214_ VGND VGND VPWR VPWR _2220_
+ sky130_fd_sc_hd__and3_1
X_3212_ cordic_inst.cordic_inst.y\[21\] cordic_inst.cordic_inst.sin_out\[21\] net214
+ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux2_1
X_4192_ cordic_inst.cordic_inst.sin_out\[19\] _2151_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__or2_1
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3143_ _1355_ _1357_ _1432_ net177 VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__a31o_1
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3074_ _1332_ _1368_ _1376_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__a21bo_1
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3976_ axi_controller.write_addr_reg\[25\] net53 net189 VGND VGND VPWR VPWR _0324_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2927_ _1229_ cordic_inst.cordic_inst.x\[30\] VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and2b_1
X_2858_ _1105_ _1111_ net290 VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__mux2_1
X_2789_ net241 _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__nand2_1
X_4528_ net353 _0260_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[10\] sky130_fd_sc_hd__dfxtp_1
X_4459_ net329 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__inv_2
XFILLER_46_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3830_ cordic_inst.done_d axi_controller.done VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__nand2b_1
X_3761_ axi_controller.reg_input_data\[3\] axi_controller.reg_input_data\[2\] axi_controller.reg_input_data\[1\]
+ axi_controller.reg_input_data\[0\] VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__or4_1
X_2712_ net186 _1030_ _1033_ net167 cordic_inst.cordic_inst.y\[18\] VGND VGND VPWR
+ VPWR _0548_ sky130_fd_sc_hd__a32o_1
XFILLER_9_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3692_ net252 _1822_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_30_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2643_ _0976_ _0977_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__or2_1
X_2574_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__inv_2
X_4313_ net135 net194 net157 axi_controller.result_out\[30\] VGND VGND VPWR VPWR _0564_
+ sky130_fd_sc_hd__a22o_1
X_4244_ net313 _2204_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__nor2_1
X_4175_ net260 _2143_ cordic_inst.cordic_inst.sin_out\[18\] VGND VGND VPWR VPWR _2144_
+ sky130_fd_sc_hd__a21o_1
X_3126_ _1375_ _1420_ _1343_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__a21o_1
X_3057_ _1201_ _1217_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_38_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3959_ axi_controller.write_addr_reg\[8\] net66 net187 VGND VGND VPWR VPWR _0307_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2290_ _0614_ cordic_inst.cordic_inst.state\[0\] VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__nor2_1
X_4931_ net372 _0032_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4862_ net375 _0071_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3813_ _1908_ _1906_ axi_controller.reg_input_data\[27\] VGND VGND VPWR VPWR _1909_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4793_ net392 _0520_ _0215_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_9_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3744_ cordic_inst.deg_handler_inst.theta_norm\[25\] _1855_ VGND VGND VPWR VPWR _0025_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3675_ cordic_inst.deg_handler_inst.theta_abs\[26\] net152 VGND VGND VPWR VPWR _0071_
+ sky130_fd_sc_hd__and2_1
X_2626_ _0915_ _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__or2_1
Xoutput122 net122 VGND VGND VPWR VPWR rdata[19] sky130_fd_sc_hd__buf_2
Xoutput133 net133 VGND VGND VPWR VPWR rdata[29] sky130_fd_sc_hd__buf_2
Xoutput111 net111 VGND VGND VPWR VPWR bvalid sky130_fd_sc_hd__buf_2
Xoutput144 net144 VGND VGND VPWR VPWR rresp[1] sky130_fd_sc_hd__buf_2
X_2557_ cordic_inst.cordic_inst.y\[2\] _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__and2_1
X_2488_ cordic_inst.cordic_inst.y\[22\] _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__nand2_1
X_4227_ cordic_inst.cordic_inst.cos_out\[24\] net223 _2188_ net316 VGND VGND VPWR
+ VPWR _2190_ sky130_fd_sc_hd__a31o_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4158_ net260 _2128_ cordic_inst.cordic_inst.sin_out\[16\] VGND VGND VPWR VPWR _2129_
+ sky130_fd_sc_hd__a21o_1
X_4089_ net225 _2068_ cordic_inst.cordic_inst.cos_out\[7\] VGND VGND VPWR VPWR _2069_
+ sky130_fd_sc_hd__a21oi_1
X_3109_ _1236_ _1401_ _1237_ _1234_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__a211o_1
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_2
Xfanout371 net388 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_2
Xfanout382 net383 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_2
Xfanout393 net408 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_2
XFILLER_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 araddr[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_30_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput46 awaddr[19] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 arvalid VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput24 araddr[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput57 awaddr[29] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 awvalid VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput79 wdata[17] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
X_3460_ _1650_ _1654_ _1490_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__a21o_1
X_2411_ net283 _0744_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a21oi_1
X_3391_ net241 _1578_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__nand2_1
X_2342_ net265 _0655_ _0658_ _0675_ net244 _0607_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux4_1
X_4012_ net89 _2009_ _2012_ net346 VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o211a_1
X_2273_ axi_controller.state\[0\] VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__inv_2
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4914_ net359 _0013_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_4845_ net366 _0084_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4776_ net390 _0503_ _0198_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3727_ net253 _1844_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__nand2_1
X_3658_ cordic_inst.deg_handler_inst.theta_abs\[18\] _1787_ VGND VGND VPWR VPWR _1807_
+ sky130_fd_sc_hd__xnor2_1
X_3589_ net180 net161 net303 VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux2_1
X_2609_ _0677_ _0943_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__xor2_1
XFILLER_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout190 _1929_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_2
XFILLER_19_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2960_ cordic_inst.cordic_inst.x\[3\] _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _1190_ _1192_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__or3_1
X_4630_ net398 _0361_ net336 VGND VGND VPWR VPWR axi_controller.result_out\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4561_ net354 _0293_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[27\] sky130_fd_sc_hd__dfxtp_1
X_4492_ net334 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__inv_2
X_3512_ _1540_ _1729_ _1730_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__o21ba_1
X_3443_ cordic_inst.cordic_inst.angle\[28\] net174 net162 cordic_inst.cordic_inst.z\[28\]
+ _1678_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a221o_1
X_3374_ _1498_ _1510_ _1577_ _1612_ net232 VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__o32a_1
X_2325_ cordic_inst.cordic_inst.x\[19\] cordic_inst.cordic_inst.x\[20\] cordic_inst.cordic_inst.x\[21\]
+ cordic_inst.cordic_inst.x\[22\] net311 net300 VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux4_1
XFILLER_38_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4828_ net392 _0555_ _0250_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[25\] sky130_fd_sc_hd__dfrtp_4
X_4759_ net394 _0486_ _0181_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_31_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3090_ cordic_inst.cordic_inst.x\[25\] _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__and2_1
X_3992_ net93 net313 _1999_ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__mux2_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2943_ _1116_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__xor2_1
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2874_ _1173_ _1176_ net275 VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4613_ net351 _0345_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[31\] sky130_fd_sc_hd__dfxtp_1
X_4544_ net355 _0276_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[10\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap154 _0743_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
X_4475_ net332 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__inv_2
X_3426_ _1663_ _1664_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__nor2_1
X_3357_ cordic_inst.cordic_inst.z\[1\] _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__and2_1
X_2308_ net239 _0642_ _0637_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a21bo_1
X_3288_ _1525_ _1526_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ cordic_inst.cordic_inst.y\[14\] _0923_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4260_ cordic_inst.cordic_inst.cos_out\[28\] _2218_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__xnor2_1
X_4191_ _2154_ _2158_ axi_controller.result_out\[19\] net205 VGND VGND VPWR VPWR _0373_
+ sky130_fd_sc_hd__o2bb2a_1
X_3211_ cordic_inst.cordic_inst.y\[22\] cordic_inst.cordic_inst.sin_out\[22\] net208
+ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux2_1
X_3142_ _1357_ _1432_ _1355_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__a21oi_1
X_3073_ _1349_ _1375_ _1372_ _1370_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__o211a_1
XFILLER_35_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3975_ axi_controller.write_addr_reg\[24\] net52 net190 VGND VGND VPWR VPWR _0323_
+ sky130_fd_sc_hd__mux2_1
X_2926_ _1077_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2857_ net218 _1108_ _1158_ net283 VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__a22o_1
XFILLER_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2788_ net233 _1087_ _1071_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a21o_1
X_4527_ net352 _0259_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4458_ net329 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__inv_2
X_3409_ _1646_ _1647_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__nor2_1
X_4389_ net324 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
XFILLER_46_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3760_ axi_controller.reg_input_data\[15\] axi_controller.reg_input_data\[14\] axi_controller.reg_input_data\[13\]
+ axi_controller.reg_input_data\[12\] VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__or4_1
X_2711_ _0858_ _1029_ _0854_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_30_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3691_ cordic_inst.deg_handler_inst.theta_norm\[5\] cordic_inst.deg_handler_inst.theta_norm\[4\]
+ _1819_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_10_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2642_ cordic_inst.cordic_inst.y\[24\] _0975_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__nor2_1
X_2573_ _0906_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and2_1
X_4312_ net136 net194 net157 axi_controller.result_out\[31\] VGND VGND VPWR VPWR _0563_
+ sky130_fd_sc_hd__a22o_1
X_4243_ cordic_inst.deg_handler_inst.kuadran\[0\] _2203_ _0605_ VGND VGND VPWR VPWR
+ _2204_ sky130_fd_sc_hd__o21a_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4174_ cordic_inst.cordic_inst.sin_out\[17\] cordic_inst.cordic_inst.sin_out\[16\]
+ _2128_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__or3_1
X_3125_ _1359_ _1362_ _1367_ _1332_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__or4b_1
X_3056_ _1355_ _1358_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__or2_1
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3958_ axi_controller.write_addr_reg\[7\] net65 net187 VGND VGND VPWR VPWR _0306_
+ sky130_fd_sc_hd__mux2_1
X_3889_ axi_controller.reg_input_data\[11\] _1964_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__or2_1
X_2909_ _1070_ _1181_ net274 VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4930_ net375 _0031_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4861_ net374 _0070_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[25\] sky130_fd_sc_hd__dfxtp_1
X_3812_ _1907_ _1908_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_15_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4792_ net392 _0519_ _0214_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[21\] sky130_fd_sc_hd__dfrtp_2
X_3743_ net255 _1854_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__nand2_1
XFILLER_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3674_ cordic_inst.deg_handler_inst.theta_abs\[25\] net153 VGND VGND VPWR VPWR _0070_
+ sky130_fd_sc_hd__and2_1
X_2625_ _0936_ _0948_ _0955_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__or4_1
Xoutput112 net112 VGND VGND VPWR VPWR rdata[0] sky130_fd_sc_hd__buf_2
Xoutput123 net123 VGND VGND VPWR VPWR rdata[1] sky130_fd_sc_hd__buf_2
Xoutput134 net134 VGND VGND VPWR VPWR rdata[2] sky130_fd_sc_hd__buf_2
Xoutput145 net145 VGND VGND VPWR VPWR rvalid sky130_fd_sc_hd__buf_2
X_2556_ _0738_ _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__xnor2_1
X_2487_ _0794_ _0799_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__xnor2_1
X_4226_ net224 _2188_ cordic_inst.cordic_inst.cos_out\[24\] VGND VGND VPWR VPWR _2189_
+ sky130_fd_sc_hd__a21oi_1
X_4157_ cordic_inst.cordic_inst.sin_out\[15\] _2123_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__or2_1
X_3108_ _1234_ _1237_ _1401_ _1236_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__o211ai_1
X_4088_ cordic_inst.cordic_inst.cos_out\[6\] cordic_inst.cordic_inst.cos_out\[5\]
+ cordic_inst.cordic_inst.cos_out\[4\] _2048_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__or4_2
X_3039_ cordic_inst.cordic_inst.x\[20\] _1340_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__or2_1
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout350 net34 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_2
Xfanout361 net388 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_2
Xfanout372 net373 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_2
Xfanout383 net387 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_2
Xfanout394 net408 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 awaddr[0] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 araddr[30] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 araddr[20] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput58 awaddr[2] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput69 bready VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
Xinput47 awaddr[1] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
X_2410_ net218 _0700_ _0704_ net221 VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a22o_1
X_3390_ _1532_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__nand2_1
X_2341_ net239 _0658_ _0637_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a21bo_1
X_2272_ net296 VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__inv_2
X_4011_ axi_controller.reg_input_data\[26\] _2008_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__or2_1
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4913_ net359 _0012_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4844_ net366 _0083_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[8\] sky130_fd_sc_hd__dfxtp_1
X_4775_ net390 _0502_ _0197_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[4\] sky130_fd_sc_hd__dfrtp_4
X_3726_ cordic_inst.deg_handler_inst.theta_norm\[18\] _1842_ VGND VGND VPWR VPWR _1844_
+ sky130_fd_sc_hd__or2_1
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3657_ _1774_ _1787_ net149 net151 cordic_inst.deg_handler_inst.theta_abs\[17\] VGND
+ VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a32o_1
X_3588_ net296 net161 _1509_ net179 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a22o_1
X_2608_ net154 _0758_ _0764_ net250 VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__a31o_1
XFILLER_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2539_ cordic_inst.cordic_inst.y\[7\] _0872_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__nor2_1
XFILLER_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4209_ net224 _2173_ cordic_inst.cordic_inst.cos_out\[22\] VGND VGND VPWR VPWR _2174_
+ sky130_fd_sc_hd__a21o_1
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout180 net181 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_2
Xfanout191 net192 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_2
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2890_ net262 _1075_ _1114_ _1106_ net238 net243 VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__mux4_2
XFILLER_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4560_ net355 _0292_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4491_ net334 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__inv_2
X_3511_ _1540_ _1729_ net175 VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__a21o_1
X_3442_ _1477_ _1666_ _1677_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__a21oi_1
X_3373_ net280 net302 VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__or2_1
X_2324_ _0655_ _0658_ net285 VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux2_1
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4827_ net392 _0554_ _0249_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[24\] sky130_fd_sc_hd__dfrtp_4
X_4758_ net403 _0485_ _0180_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_3709_ cordic_inst.deg_handler_inst.theta_norm\[12\] _1833_ VGND VGND VPWR VPWR _0011_
+ sky130_fd_sc_hd__xnor2_1
X_4689_ net405 _0416_ _0111_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3991_ net350 _2000_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2_1
X_2942_ _1131_ _1178_ net251 VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a21o_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2873_ net286 _1174_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_20_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4612_ net352 _0344_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[30\] sky130_fd_sc_hd__dfxtp_1
X_4543_ net351 _0275_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[9\] sky130_fd_sc_hd__dfxtp_1
X_4474_ net332 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__inv_2
X_3425_ cordic_inst.cordic_inst.z\[27\] cordic_inst.cordic_inst.z\[26\] net249 VGND
+ VGND VPWR VPWR _1664_ sky130_fd_sc_hd__o21a_1
X_3356_ _1585_ _1587_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__xnor2_1
X_3287_ cordic_inst.cordic_inst.z\[15\] _1524_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__nand2_1
X_2307_ net234 _0641_ _0635_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__a21o_1
XFILLER_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3210_ cordic_inst.cordic_inst.y\[23\] cordic_inst.cordic_inst.sin_out\[23\] net208
+ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux2_1
X_4190_ _2156_ _2157_ net205 VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__o21a_1
X_3141_ _1358_ _1431_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__or2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3072_ _1359_ _1365_ _1373_ _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__o31a_1
XFILLER_36_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3974_ axi_controller.write_addr_reg\[23\] net51 net189 VGND VGND VPWR VPWR _0322_
+ sky130_fd_sc_hd__mux2_1
X_2925_ net269 _1227_ _1226_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__a21oi_1
X_2856_ net216 _1142_ _1144_ _0713_ net275 VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a221o_1
X_2787_ net274 _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__nor2_1
X_4526_ net352 _0258_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[8\] sky130_fd_sc_hd__dfxtp_1
X_4457_ net322 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__inv_2
X_3408_ cordic_inst.cordic_inst.z\[17\] _1644_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__and2_1
X_4388_ net324 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
X_3339_ _1498_ _1577_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__nor2_1
XFILLER_39_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2710_ _1031_ _1032_ cordic_inst.cordic_inst.y\[19\] net167 VGND VGND VPWR VPWR _0549_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3690_ cordic_inst.deg_handler_inst.theta_norm\[5\] _1821_ VGND VGND VPWR VPWR _0035_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2641_ cordic_inst.cordic_inst.y\[24\] _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__and2_1
X_2572_ cordic_inst.cordic_inst.y\[4\] _0886_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_10_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4311_ net194 _1976_ _1987_ _2252_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__and4b_4
X_4242_ cordic_inst.cordic_inst.cos_out\[25\] _2196_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__nor2_1
X_4173_ _2139_ _2142_ axi_controller.result_out\[17\] net204 VGND VGND VPWR VPWR _0371_
+ sky130_fd_sc_hd__o2bb2a_1
X_3124_ net181 _1382_ _1419_ net164 cordic_inst.cordic_inst.x\[24\] VGND VGND VPWR
+ VPWR _0522_ sky130_fd_sc_hd__a32o_1
XFILLER_28_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3055_ cordic_inst.cordic_inst.x\[18\] _1356_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3957_ axi_controller.write_addr_reg\[6\] net64 net187 VGND VGND VPWR VPWR _0305_
+ sky130_fd_sc_hd__mux2_1
X_2908_ net242 _1183_ net215 VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__a21o_1
X_3888_ net72 _1965_ _1968_ net346 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__o211a_1
X_2839_ cordic_inst.cordic_inst.y\[4\] cordic_inst.cordic_inst.y\[5\] net308 VGND
+ VGND VPWR VPWR _1142_ sky130_fd_sc_hd__mux2_1
XFILLER_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4509_ net332 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__inv_2
XFILLER_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4860_ net372 _0069_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ axi_controller.reg_input_data\[26\] axi_controller.reg_input_data\[25\] _1903_
+ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_15_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4791_ net394 _0518_ _0213_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[20\] sky130_fd_sc_hd__dfrtp_4
X_3742_ cordic_inst.deg_handler_inst.theta_norm\[24\] _1852_ VGND VGND VPWR VPWR _1854_
+ sky130_fd_sc_hd__or2_1
X_3673_ cordic_inst.deg_handler_inst.theta_abs\[24\] net152 VGND VGND VPWR VPWR _0069_
+ sky130_fd_sc_hd__and2_1
X_2624_ _0957_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nand2_1
Xoutput124 net124 VGND VGND VPWR VPWR rdata[20] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR rdata[10] sky130_fd_sc_hd__buf_2
Xoutput135 net135 VGND VGND VPWR VPWR rdata[30] sky130_fd_sc_hd__buf_2
Xoutput146 net146 VGND VGND VPWR VPWR wready sky130_fd_sc_hd__buf_2
X_2555_ _0718_ _0735_ net272 VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__o21ai_1
X_2486_ _0817_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__or2_1
X_4225_ cordic_inst.cordic_inst.cos_out\[23\] cordic_inst.cordic_inst.cos_out\[22\]
+ _2173_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__or3_1
X_4156_ axi_controller.result_out\[15\] net204 _2127_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__o21ba_1
X_3107_ cordic_inst.cordic_inst.x\[30\] net163 _1408_ net179 VGND VGND VPWR VPWR _0528_
+ sky130_fd_sc_hd__a22o_1
X_4087_ net258 _2065_ cordic_inst.cordic_inst.sin_out\[7\] VGND VGND VPWR VPWR _2067_
+ sky130_fd_sc_hd__a21oi_1
X_3038_ cordic_inst.cordic_inst.x\[20\] _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__nand2_1
XFILLER_11_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout340 net344 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__buf_4
Xfanout373 net374 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
Xfanout351 net354 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_2
Xfanout362 net365 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_2
Xfanout384 net387 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_2
Xfanout395 net408 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput37 awaddr[10] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput15 araddr[21] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 araddr[31] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput59 awaddr[30] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
Xinput48 awaddr[20] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
XFILLER_6_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2340_ _0673_ _0674_ net292 VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__mux2_1
X_2271_ net289 VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__inv_2
X_4010_ net88 _2009_ _2011_ net347 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__o211a_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4912_ net359 _0011_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4843_ net366 _0082_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[7\] sky130_fd_sc_hd__dfxtp_1
X_4774_ net389 _0501_ _0196_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3725_ cordic_inst.deg_handler_inst.theta_norm\[18\] _1843_ VGND VGND VPWR VPWR _0017_
+ sky130_fd_sc_hd__xnor2_1
X_3656_ _1773_ net147 _1806_ net151 cordic_inst.deg_handler_inst.theta_abs\[16\] VGND
+ VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a32o_1
X_3587_ net179 _1576_ _1581_ net161 net289 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a32o_1
X_2607_ _0940_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2538_ cordic_inst.cordic_inst.y\[7\] _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__and2_1
X_2469_ net273 _0797_ _0803_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a21o_1
X_4208_ cordic_inst.cordic_inst.cos_out\[21\] _2166_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__or2_1
X_4139_ cordic_inst.cordic_inst.cos_out\[13\] net227 _2111_ net315 VGND VGND VPWR
+ VPWR _2113_ sky130_fd_sc_hd__a31o_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout192 net193 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_4
Xfanout181 net182 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xfanout170 _0630_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
XFILLER_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3510_ _1545_ _1623_ _1544_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4490_ net330 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
X_3441_ net176 _1667_ VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__or2_1
X_3372_ _1554_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__or2_1
X_2323_ net265 _0632_ _0640_ _0656_ _0609_ net234 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux4_2
XFILLER_38_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4826_ net394 _0553_ _0248_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[23\] sky130_fd_sc_hd__dfrtp_4
X_4757_ net404 _0484_ _0179_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3708_ net253 _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__nand2_1
X_4688_ net405 _0415_ _0110_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_3639_ cordic_inst.deg_handler_inst.theta_abs\[8\] _1764_ VGND VGND VPWR VPWR _1798_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3990_ net71 net319 _1999_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__mux2_1
X_2941_ cordic_inst.cordic_inst.x\[7\] _1242_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__nand2_1
XFILLER_30_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4611_ net352 _0343_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2872_ net233 _1079_ _1071_ net238 VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__a211o_1
XFILLER_31_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4542_ net351 _0274_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[8\] sky130_fd_sc_hd__dfxtp_1
X_4473_ net344 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__inv_2
X_3424_ cordic_inst.cordic_inst.z\[25\] cordic_inst.cordic_inst.z\[24\] net248 VGND
+ VGND VPWR VPWR _1663_ sky130_fd_sc_hd__o21a_1
X_3355_ cordic_inst.cordic_inst.z\[2\] _1593_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__nand2_1
X_3286_ cordic_inst.cordic_inst.z\[15\] _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__or2_1
X_2306_ cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.x\[29\] cordic_inst.cordic_inst.x\[30\]
+ net265 net305 net296 VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4809_ net396 _0536_ _0231_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[6\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ _1373_ _1430_ _1365_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__a21o_1
X_3071_ _1354_ _1357_ _1353_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__a21o_1
X_3973_ axi_controller.write_addr_reg\[22\] net50 net189 VGND VGND VPWR VPWR _0321_
+ sky130_fd_sc_hd__mux2_1
X_2924_ net274 _1191_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__nor2_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2855_ _1104_ _1107_ net235 VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__mux2_1
X_2786_ net238 _1088_ _1070_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__a21boi_1
X_4525_ net368 _0004_ VGND VGND VPWR VPWR axi_controller.state\[3\] sky130_fd_sc_hd__dfxtp_1
X_4456_ net323 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__inv_2
X_3407_ _1645_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__inv_2
X_4387_ net324 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
X_3338_ _0711_ _1576_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__nor2_1
X_3269_ net222 _0707_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__nand2_1
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2640_ _0795_ _0801_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2571_ _0902_ _0904_ _0889_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4310_ net82 net103 _1930_ _1994_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__and4_1
X_4241_ axi_controller.result_out\[25\] _2202_ net201 VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux2_1
XFILLER_4_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4172_ net314 _2141_ net204 VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__o21a_1
X_3123_ _1377_ _1381_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__or2_1
X_3054_ cordic_inst.cordic_inst.x\[18\] _1356_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__nand2_1
XFILLER_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3956_ axi_controller.write_addr_reg\[5\] net63 net188 VGND VGND VPWR VPWR _0304_
+ sky130_fd_sc_hd__mux2_1
X_2907_ net246 _1115_ _1068_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a21o_1
X_3887_ axi_controller.reg_input_data\[10\] _1964_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__or2_1
X_2838_ _1139_ _1140_ net291 VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__mux2_1
X_2769_ net263 net295 VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__and2_1
XFILLER_2_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4508_ net332 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__inv_2
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4439_ net343 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__inv_2
XFILLER_46_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3810_ axi_controller.reg_input_data\[27\] _1905_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_15_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4790_ net403 _0517_ _0212_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[19\] sky130_fd_sc_hd__dfrtp_2
X_3741_ cordic_inst.deg_handler_inst.theta_norm\[24\] _1853_ VGND VGND VPWR VPWR _0024_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3672_ cordic_inst.deg_handler_inst.theta_abs\[23\] cordic_inst.deg_handler_inst.theta_abs\[31\]
+ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__and2_1
X_2623_ _0598_ _0956_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__nand2_1
Xoutput125 net125 VGND VGND VPWR VPWR rdata[21] sky130_fd_sc_hd__buf_2
X_2554_ cordic_inst.cordic_inst.y\[3\] _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__and2_1
Xoutput114 net114 VGND VGND VPWR VPWR rdata[11] sky130_fd_sc_hd__buf_2
Xoutput136 net136 VGND VGND VPWR VPWR rdata[31] sky130_fd_sc_hd__buf_2
X_2485_ _0595_ _0816_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__and2_1
X_4224_ axi_controller.result_out\[24\] net201 VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__nor2_1
X_4155_ _2121_ _2122_ _2126_ net204 VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__o211a_1
X_3106_ _1231_ _1402_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__xor2_1
X_4086_ cordic_inst.cordic_inst.sin_out\[7\] net258 _2065_ VGND VGND VPWR VPWR _2066_
+ sky130_fd_sc_hd__and3_1
X_3037_ _1208_ _1218_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__xor2_1
XFILLER_36_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3939_ axi_controller.read_addr_reg\[29\] axi_controller.read_addr_reg\[30\] VGND
+ VGND VPWR VPWR _1982_ sky130_fd_sc_hd__nand2_1
XFILLER_3_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout330 net345 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__buf_2
Xfanout341 net342 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__buf_4
Xfanout374 net378 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_2
Xfanout352 net354 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_2
Xfanout363 net364 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
Xfanout385 net387 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_2
Xfanout396 net397 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 araddr[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
Xinput16 araddr[22] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput49 awaddr[21] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 awaddr[11] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
X_2270_ net282 VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__inv_2
XFILLER_38_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4911_ net360 _0010_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4842_ net366 _0081_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4773_ net389 _0500_ _0195_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3724_ net253 _1842_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__nand2_1
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3655_ cordic_inst.deg_handler_inst.theta_abs\[16\] _1772_ VGND VGND VPWR VPWR _1806_
+ sky130_fd_sc_hd__nand2_1
X_2606_ _0938_ cordic_inst.cordic_inst.y\[11\] VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__and2b_1
X_3586_ _1756_ _1757_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and2_1
X_2537_ _0684_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__xor2_1
X_2468_ net273 _0796_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21o_1
X_4207_ axi_controller.result_out\[21\] _2172_ net205 VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
X_2399_ net284 _0728_ _0732_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__a211o_1
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4138_ net227 _2111_ cordic_inst.cordic_inst.cos_out\[13\] VGND VGND VPWR VPWR _2112_
+ sky130_fd_sc_hd__a21oi_1
X_4069_ net202 _2051_ _2044_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout182 _0626_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_4
Xfanout171 net172 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xfanout160 _0629_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
Xfanout193 _1927_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3440_ net181 _1675_ _1676_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a21o_1
X_3371_ _1561_ _1608_ _1556_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__o21ba_1
X_2322_ _0640_ _0656_ _0609_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4825_ net394 _0552_ _0247_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[22\] sky130_fd_sc_hd__dfrtp_2
X_4756_ net407 _0483_ _0178_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_3707_ cordic_inst.deg_handler_inst.theta_norm\[11\] cordic_inst.deg_handler_inst.theta_norm\[10\]
+ _1829_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__or3_1
X_4687_ net400 _0414_ _0109_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3638_ _1764_ net147 _1797_ net150 cordic_inst.deg_handler_inst.theta_abs\[7\] VGND
+ VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a32o_1
X_3569_ cordic_inst.cordic_inst.x\[10\] cordic_inst.cordic_inst.cos_out\[10\] net211
+ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2940_ cordic_inst.cordic_inst.x\[7\] _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__nor2_1
X_2871_ _1133_ _1135_ net291 VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__mux2_1
X_4610_ net357 _0342_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4541_ net364 _0273_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4472_ net344 VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__inv_2
X_3423_ _1660_ _1661_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__nand2_1
X_3354_ _1582_ _1588_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__xor2_1
X_3285_ net267 _1481_ _1523_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__mux2_1
X_2305_ cordic_inst.cordic_inst.x\[28\] cordic_inst.cordic_inst.x\[29\] net304 VGND
+ VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux2_1
XFILLER_39_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4808_ net396 _0535_ _0230_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[5\] sky130_fd_sc_hd__dfrtp_2
X_4739_ net390 _0466_ _0161_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_8_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3070_ cordic_inst.cordic_inst.x\[16\] _1360_ _1364_ cordic_inst.cordic_inst.x\[17\]
+ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__a22oi_1
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3972_ axi_controller.write_addr_reg\[21\] net49 net190 VGND VGND VPWR VPWR _0320_
+ sky130_fd_sc_hd__mux2_1
X_2923_ _1082_ _1225_ net269 VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__o21a_1
X_2854_ _1153_ _1155_ _1156_ _1151_ net243 VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__o32a_1
X_2785_ _1084_ _1087_ net291 VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__mux2_1
X_4524_ net368 _0003_ VGND VGND VPWR VPWR axi_controller.state\[2\] sky130_fd_sc_hd__dfxtp_1
X_4455_ net322 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__inv_2
X_3406_ cordic_inst.cordic_inst.z\[17\] _1644_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__or2_1
X_4386_ net324 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
X_3337_ net296 net303 net289 VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__a21o_1
X_3268_ net248 _0705_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__or2_1
X_3199_ _0603_ net174 VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__nor2_1
XFILLER_27_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2570_ _0902_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4240_ axi_controller.mode _2197_ _2198_ _2200_ _2201_ VGND VGND VPWR VPWR _2202_
+ sky130_fd_sc_hd__o32ai_1
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4171_ cordic_inst.cordic_inst.cos_out\[17\] _2140_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__xnor2_1
X_3122_ cordic_inst.cordic_inst.x\[25\] net163 _1418_ net181 VGND VGND VPWR VPWR _0523_
+ sky130_fd_sc_hd__a22o_1
X_3053_ _1204_ _1350_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__xor2_1
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3955_ axi_controller.write_addr_reg\[4\] net62 net188 VGND VGND VPWR VPWR _0303_
+ sky130_fd_sc_hd__mux2_1
X_2906_ _1206_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__nand2_1
X_3886_ net102 _1965_ _1967_ net347 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o211a_1
X_2837_ cordic_inst.cordic_inst.y\[12\] cordic_inst.cordic_inst.y\[13\] cordic_inst.cordic_inst.y\[14\]
+ cordic_inst.cordic_inst.y\[15\] net310 net299 VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__mux4_2
XFILLER_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2768_ net263 net293 VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and2_1
X_2699_ cordic_inst.cordic_inst.y\[23\] net165 _1025_ net186 VGND VGND VPWR VPWR _0553_
+ sky130_fd_sc_hd__a22o_1
X_4507_ net333 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__inv_2
X_4438_ net343 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
X_4369_ net337 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3740_ net254 _1852_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__nand2_1
X_3671_ net149 _1814_ _1815_ net152 cordic_inst.deg_handler_inst.theta_abs\[22\] VGND
+ VGND VPWR VPWR _0067_ sky130_fd_sc_hd__a32o_1
X_2622_ _0598_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__or2_1
X_2553_ _0742_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__xnor2_1
Xoutput115 net115 VGND VGND VPWR VPWR rdata[12] sky130_fd_sc_hd__buf_2
Xoutput126 net126 VGND VGND VPWR VPWR rdata[22] sky130_fd_sc_hd__buf_2
Xoutput137 net137 VGND VGND VPWR VPWR rdata[3] sky130_fd_sc_hd__buf_2
X_2484_ cordic_inst.cordic_inst.y\[29\] _0814_ _0817_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a21oi_1
X_4223_ _2183_ _2186_ axi_controller.result_out\[23\] net201 VGND VGND VPWR VPWR _0377_
+ sky130_fd_sc_hd__o2bb2a_1
X_4154_ _2124_ _2125_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__or2_1
X_4085_ cordic_inst.cordic_inst.sin_out\[6\] cordic_inst.cordic_inst.sin_out\[5\]
+ cordic_inst.cordic_inst.sin_out\[4\] _2045_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__or4_1
X_3105_ net179 _1406_ _1407_ net163 net265 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a32o_1
XFILLER_28_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3036_ _1337_ _1338_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__nand2_1
XFILLER_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3938_ axi_controller.read_addr_reg\[17\] _1980_ axi_controller.read_addr_reg\[2\]
+ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__or3b_1
X_3869_ axi_controller.write_addr_reg\[12\] axi_controller.write_addr_reg\[15\] axi_controller.write_addr_reg\[14\]
+ axi_controller.write_addr_reg\[17\] VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__or4_1
Xfanout320 axi_controller.rst VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_4
Xfanout331 net333 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__buf_4
Xfanout375 net377 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
Xfanout353 net354 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_1
Xfanout342 net343 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_2
Xfanout364 net365 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_2
Xfanout397 net408 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout386 net387 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 araddr[23] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 araddr[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 awaddr[12] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4910_ net360 _0009_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4841_ net366 _0080_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[5\] sky130_fd_sc_hd__dfxtp_1
X_4772_ net390 _0499_ _0194_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[1\] sky130_fd_sc_hd__dfrtp_2
X_3723_ cordic_inst.deg_handler_inst.theta_norm\[17\] cordic_inst.deg_handler_inst.theta_norm\[16\]
+ _1839_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__or3_1
X_3654_ _1772_ net147 _1805_ net151 cordic_inst.deg_handler_inst.theta_abs\[15\] VGND
+ VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a32o_1
X_2605_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__inv_2
X_3585_ net158 _1580_ net282 VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__a21o_1
X_2536_ _0693_ _0743_ _0757_ net250 VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__a31o_1
X_2467_ net273 _0795_ _0801_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__a21bo_1
X_4206_ net316 _2170_ _2171_ _2167_ _2168_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__a32o_1
X_2398_ cordic_inst.cordic_inst.x\[1\] net222 _0711_ _0730_ net219 VGND VGND VPWR
+ VPWR _0733_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_39_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4137_ cordic_inst.cordic_inst.cos_out\[12\] cordic_inst.cordic_inst.cos_out\[11\]
+ cordic_inst.cordic_inst.cos_out\[10\] _2089_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__or4_2
X_4068_ net228 _2046_ _2047_ _2049_ _2050_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__o32a_1
X_3019_ cordic_inst.cordic_inst.x\[10\] _1320_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__or2_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout161 net162 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net186 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_4
Xfanout172 _0628_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_4
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_2
Xfanout194 _1927_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_34_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3370_ _1561_ _1608_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__nor2_1
X_2321_ cordic_inst.cordic_inst.x\[26\] cordic_inst.cordic_inst.x\[27\] net304 VGND
+ VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4824_ net395 _0551_ _0246_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[21\] sky130_fd_sc_hd__dfrtp_2
X_4755_ net407 _0482_ _0177_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3706_ cordic_inst.deg_handler_inst.theta_norm\[11\] _1831_ VGND VGND VPWR VPWR _0010_
+ sky130_fd_sc_hd__xnor2_1
X_4686_ net400 _0413_ _0108_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3637_ cordic_inst.deg_handler_inst.theta_abs\[7\] _1763_ VGND VGND VPWR VPWR _1797_
+ sky130_fd_sc_hd__nand2_1
X_3568_ cordic_inst.cordic_inst.x\[11\] cordic_inst.cordic_inst.cos_out\[11\] net211
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2519_ _0852_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__nand2_1
X_3499_ cordic_inst.cordic_inst.angle\[15\] net172 net159 cordic_inst.cordic_inst.z\[15\]
+ _1721_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__a221o_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2870_ net286 _1171_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4540_ net364 _0272_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_4471_ net340 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__inv_2
X_3422_ net268 cordic_inst.cordic_inst.z\[26\] VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__xnor2_1
X_3353_ cordic_inst.cordic_inst.z\[3\] _1590_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__xnor2_1
X_3284_ _0707_ _1521_ net280 VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__a21o_1
X_2304_ _0606_ _0638_ net170 VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a21o_1
XFILLER_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4807_ net396 _0534_ _0229_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[4\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2999_ cordic_inst.cordic_inst.x\[14\] _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__nand2_1
X_4738_ net389 _0465_ _0160_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[31\] sky130_fd_sc_hd__dfrtp_1
X_4669_ net351 _0398_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[23\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_8_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3971_ axi_controller.write_addr_reg\[20\] net48 net189 VGND VGND VPWR VPWR _0319_
+ sky130_fd_sc_hd__mux2_1
X_2922_ net269 _1214_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a21o_1
X_2853_ cordic_inst.cordic_inst.y\[1\] net221 _0711_ _1121_ net218 VGND VGND VPWR
+ VPWR _1156_ sky130_fd_sc_hd__a32o_1
X_2784_ cordic_inst.cordic_inst.y\[27\] cordic_inst.cordic_inst.y\[28\] cordic_inst.cordic_inst.y\[29\]
+ cordic_inst.cordic_inst.y\[30\] net304 net295 VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__mux4_1
XFILLER_8_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4523_ net370 _0002_ VGND VGND VPWR VPWR axi_controller.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_4454_ net323 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__inv_2
X_3405_ net248 _1643_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__xnor2_1
X_4385_ net324 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
X_3336_ cordic_inst.cordic_inst.z\[4\] _1574_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__nand2_1
X_3267_ cordic_inst.cordic_inst.z\[13\] _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__and2_1
XFILLER_27_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3198_ net180 _1148_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__nand2_1
XFILLER_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4170_ cordic_inst.cordic_inst.cos_out\[16\] _2132_ net226 VGND VGND VPWR VPWR _2140_
+ sky130_fd_sc_hd__o21a_1
X_3121_ _1395_ _1417_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__xnor2_1
X_3052_ _1353_ _1354_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_18_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3954_ axi_controller.write_addr_reg\[3\] net61 net190 VGND VGND VPWR VPWR _0302_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3885_ axi_controller.reg_input_data\[9\] _1964_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__or2_1
X_2905_ net276 _1176_ _1069_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__o21a_1
X_2836_ cordic_inst.cordic_inst.y\[8\] cordic_inst.cordic_inst.y\[9\] cordic_inst.cordic_inst.y\[10\]
+ cordic_inst.cordic_inst.y\[11\] net308 net297 VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__mux4_2
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2767_ net263 net282 VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__nand2_2
X_2698_ _0830_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__xnor2_1
X_4506_ net333 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__inv_2
X_4437_ net341 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__inv_2
X_4368_ net338 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
X_4299_ axi_controller.reg_input_data\[21\] _2242_ VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__or2_1
X_3319_ net237 net302 VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__and2_1
XFILLER_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3670_ _1783_ _1808_ _0617_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__o21ai_1
X_2621_ _0760_ _0949_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__xnor2_1
X_2552_ _0718_ _0735_ _0738_ net272 VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__o31a_1
Xoutput116 net116 VGND VGND VPWR VPWR rdata[13] sky130_fd_sc_hd__buf_2
Xoutput127 net127 VGND VGND VPWR VPWR rdata[23] sky130_fd_sc_hd__buf_2
Xoutput138 net138 VGND VGND VPWR VPWR rdata[4] sky130_fd_sc_hd__buf_2
X_4222_ net316 _2185_ net201 VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__o21a_1
X_2483_ cordic_inst.cordic_inst.y\[29\] _0814_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__nand2_1
X_4153_ cordic_inst.cordic_inst.sin_out\[15\] net260 _2123_ net229 VGND VGND VPWR
+ VPWR _2125_ sky130_fd_sc_hd__a31o_1
X_4084_ axi_controller.result_out\[7\] net202 VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__nor2_1
X_3104_ _1230_ _1403_ _1405_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__or3_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3035_ cordic_inst.cordic_inst.x\[22\] _1336_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__or2_1
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3937_ axi_controller.read_addr_reg\[16\] axi_controller.read_addr_reg\[19\] axi_controller.read_addr_reg\[18\]
+ axi_controller.read_addr_reg\[21\] VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__or4_1
X_3868_ axi_controller.write_addr_reg\[8\] axi_controller.write_addr_reg\[11\] axi_controller.write_addr_reg\[10\]
+ axi_controller.write_addr_reg\[13\] VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__or4_1
X_3799_ axi_controller.reg_input_data\[23\] _1892_ axi_controller.reg_input_data\[24\]
+ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__a21oi_1
X_2819_ cordic_inst.cordic_inst.y\[9\] cordic_inst.cordic_inst.y\[10\] cordic_inst.cordic_inst.y\[11\]
+ cordic_inst.cordic_inst.y\[12\] net308 net297 VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux4_2
Xfanout321 net328 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_4
Xfanout310 net311 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_4
Xfanout332 net333 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_2
Xfanout354 net361 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_2
Xfanout365 net388 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_2
Xfanout343 net344 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
Xfanout376 net377 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout398 net399 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_2
Xfanout387 net388 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 araddr[24] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 araddr[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4840_ net367 _0079_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4771_ net390 _0498_ _0193_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[0\] sky130_fd_sc_hd__dfrtp_1
X_3722_ cordic_inst.deg_handler_inst.theta_norm\[17\] _1841_ VGND VGND VPWR VPWR _0016_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3653_ cordic_inst.deg_handler_inst.theta_abs\[15\] _1771_ VGND VGND VPWR VPWR _1805_
+ sky130_fd_sc_hd__nand2_1
X_2604_ cordic_inst.cordic_inst.y\[11\] _0938_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nand2b_1
X_3584_ _1755_ _1756_ net274 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
X_2535_ _0743_ _0757_ net250 VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21oi_1
X_2466_ net271 _0652_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a21oi_1
X_4205_ cordic_inst.cordic_inst.sin_out\[21\] net261 _2169_ VGND VGND VPWR VPWR _2171_
+ sky130_fd_sc_hd__nand3_1
X_2397_ cordic_inst.cordic_inst.x\[2\] net217 _0709_ _0731_ net275 VGND VGND VPWR
+ VPWR _0732_ sky130_fd_sc_hd__a221o_1
X_4136_ _2108_ _2109_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4067_ cordic_inst.cordic_inst.cos_out\[4\] net226 _2048_ net314 VGND VGND VPWR VPWR
+ _2050_ sky130_fd_sc_hd__a31o_1
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3018_ cordic_inst.cordic_inst.x\[10\] _1320_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__nand2_1
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout162 net164 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_2
Xfanout151 net153 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
Xfanout173 _0628_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
Xfanout195 net199 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net186 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_2
XFILLER_43_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2320_ _0653_ _0654_ net292 VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_18_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4823_ net395 _0550_ _0245_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[20\] sky130_fd_sc_hd__dfrtp_4
X_4754_ net406 _0481_ _0176_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3705_ cordic_inst.deg_handler_inst.theta_norm\[10\] _1829_ net252 VGND VGND VPWR
+ VPWR _1831_ sky130_fd_sc_hd__o21ai_1
X_4685_ net401 _0412_ _0107_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3636_ _1763_ net147 _1796_ net150 cordic_inst.deg_handler_inst.theta_abs\[6\] VGND
+ VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a32o_1
X_3567_ cordic_inst.cordic_inst.x\[12\] cordic_inst.cordic_inst.cos_out\[12\] net210
+ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_2518_ _0596_ _0851_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__nand2_1
X_3498_ _1527_ _1719_ _1720_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__a21oi_1
X_2449_ _0631_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nand2_1
XFILLER_29_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4119_ cordic_inst.cordic_inst.sin_out\[11\] net258 _2093_ net228 VGND VGND VPWR
+ VPWR _2095_ sky130_fd_sc_hd__a31o_1
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4470_ net340 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__inv_2
X_3421_ net268 cordic_inst.cordic_inst.z\[27\] VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__xnor2_1
X_3352_ cordic_inst.cordic_inst.z\[3\] _1590_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__and2_1
X_2303_ net286 _0636_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__o21ai_1
X_3283_ _1521_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__inv_2
XFILLER_38_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4806_ net391 _0533_ _0228_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2998_ _1193_ _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4737_ net376 _0464_ _0159_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[30\] sky130_fd_sc_hd__dfrtp_1
X_4668_ net357 _0397_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[22\] sky130_fd_sc_hd__dfxtp_1
X_3619_ net153 _1786_ cordic_inst.deg_handler_inst.theta_abs\[0\] VGND VGND VPWR VPWR
+ _0053_ sky130_fd_sc_hd__o21a_1
X_4599_ net369 _0331_ VGND VGND VPWR VPWR axi_controller.rst sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_8_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3970_ axi_controller.write_addr_reg\[19\] net46 net190 VGND VGND VPWR VPWR _0318_
+ sky130_fd_sc_hd__mux2_1
X_2921_ net269 _1213_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__a21o_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2852_ cordic_inst.cordic_inst.y\[2\] net217 net216 _1154_ net275 VGND VGND VPWR
+ VPWR _1155_ sky130_fd_sc_hd__a221o_1
X_2783_ cordic_inst.cordic_inst.y\[29\] cordic_inst.cordic_inst.y\[30\] net304 VGND
+ VGND VPWR VPWR _1086_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4522_ net370 _0001_ VGND VGND VPWR VPWR axi_controller.state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4453_ net324 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__inv_2
X_3404_ net288 net302 _1498_ _1502_ net280 VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__a2111o_1
X_4384_ net324 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
X_3335_ _1481_ net266 _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__mux2_1
X_3266_ net267 _1503_ _1504_ _1501_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3197_ net181 _1272_ _1469_ net165 cordic_inst.cordic_inst.x\[1\] VGND VGND VPWR
+ VPWR _0499_ sky130_fd_sc_hd__a32o_1
XFILLER_27_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3120_ _1377_ _1381_ _1379_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__a21oi_1
X_3051_ cordic_inst.cordic_inst.x\[19\] _1352_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__nand2_1
XFILLER_36_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ axi_controller.write_addr_reg\[2\] net58 net187 VGND VGND VPWR VPWR _0301_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3884_ net101 _1965_ _1966_ net346 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__o211a_1
X_2904_ _1069_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__nand2_1
X_2835_ net242 _1137_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__or2_1
X_2766_ net262 net276 VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nand2_1
X_2697_ _0825_ _1023_ _0823_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__a21bo_1
X_4505_ net333 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__inv_2
X_4436_ net341 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__inv_2
X_4367_ net334 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
X_3318_ net280 net237 _0712_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__a21oi_1
X_4298_ net83 _2243_ _2248_ net346 VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o211a_1
X_3249_ cordic_inst.cordic_inst.z\[20\] _1487_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__nand2_1
XFILLER_27_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2620_ _0952_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nand2_1
X_2551_ _0750_ _0880_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__xnor2_1
Xoutput128 net128 VGND VGND VPWR VPWR rdata[24] sky130_fd_sc_hd__buf_2
Xoutput139 net139 VGND VGND VPWR VPWR rdata[5] sky130_fd_sc_hd__buf_2
Xoutput117 net117 VGND VGND VPWR VPWR rdata[14] sky130_fd_sc_hd__buf_2
X_2482_ _0595_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__nor2_1
X_4221_ cordic_inst.cordic_inst.cos_out\[23\] _2184_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__xnor2_1
X_4152_ net260 _2123_ cordic_inst.cordic_inst.sin_out\[15\] VGND VGND VPWR VPWR _2124_
+ sky130_fd_sc_hd__a21oi_1
X_4083_ axi_controller.result_out\[6\] _2063_ net202 VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux2_1
X_3103_ _1230_ _1403_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__o21ai_1
X_3034_ cordic_inst.cordic_inst.x\[22\] _1336_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__nand2_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3936_ _1976_ _1978_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__nand2_1
X_3867_ axi_controller.write_addr_reg\[1\] axi_controller.write_addr_reg\[0\] _1949_
+ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__or3_1
X_3798_ _1896_ _1897_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__xnor2_1
X_2818_ cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.y\[6\] cordic_inst.cordic_inst.y\[7\]
+ cordic_inst.cordic_inst.y\[8\] net308 net297 VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__mux4_1
X_2749_ net185 _1058_ _1059_ net168 cordic_inst.cordic_inst.y\[7\] VGND VGND VPWR
+ VPWR _0537_ sky130_fd_sc_hd__a32o_1
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4419_ net323 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__inv_2
Xfanout322 net323 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__buf_4
Xfanout311 net312 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_4
Xfanout300 cordic_inst.cordic_inst.i\[1\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_2
Xfanout355 net361 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_2
Xfanout366 net367 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_2
Xfanout333 net345 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__buf_4
Xfanout344 net345 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_2
Xfanout399 net402 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_2
Xfanout388 net1 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_2
Xfanout377 net378 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_2
XFILLER_27_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput19 araddr[25] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4770_ net381 _0497_ _0192_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_3721_ cordic_inst.deg_handler_inst.theta_norm\[16\] _1839_ net253 VGND VGND VPWR
+ VPWR _1841_ sky130_fd_sc_hd__o21ai_1
X_3652_ _1771_ net147 _1804_ net151 cordic_inst.deg_handler_inst.theta_abs\[14\] VGND
+ VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a32o_1
X_3583_ net174 _1755_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__nor2_1
X_2603_ _0769_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__xnor2_1
X_2534_ _0850_ _0854_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__or3b_1
X_2465_ _0789_ _0791_ _0793_ _0794_ net271 VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__o41a_1
X_4204_ net261 _2169_ cordic_inst.cordic_inst.sin_out\[21\] VGND VGND VPWR VPWR _2170_
+ sky130_fd_sc_hd__a21o_1
X_2396_ cordic_inst.cordic_inst.x\[3\] cordic_inst.cordic_inst.x\[4\] net307 VGND
+ VGND VPWR VPWR _0731_ sky130_fd_sc_hd__mux2_1
X_4135_ cordic_inst.cordic_inst.sin_out\[13\] net260 _2107_ net229 VGND VGND VPWR
+ VPWR _2109_ sky130_fd_sc_hd__a31o_1
XFILLER_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4066_ net226 _2048_ cordic_inst.cordic_inst.cos_out\[4\] VGND VGND VPWR VPWR _2049_
+ sky130_fd_sc_hd__a21oi_1
X_3017_ _1187_ _1319_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__xor2_1
XFILLER_37_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4968_ net108 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
X_4899_ net358 _0052_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_3919_ axi_controller.read_addr_reg\[20\] net14 net196 VGND VGND VPWR VPWR _0286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xcordic_system_409 VGND VGND VPWR VPWR cordic_system_409/HI bresp[0] sky130_fd_sc_hd__conb_1
Xfanout152 net153 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
Xfanout174 _0628_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xfanout163 net164 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_2
Xfanout185 net186 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net199 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_2
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4822_ net395 _0549_ _0244_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[19\] sky130_fd_sc_hd__dfrtp_4
X_4753_ net405 _0480_ _0175_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3704_ cordic_inst.deg_handler_inst.theta_norm\[10\] _1830_ VGND VGND VPWR VPWR _0009_
+ sky130_fd_sc_hd__xnor2_1
X_4684_ net396 _0411_ _0106_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3635_ cordic_inst.deg_handler_inst.theta_abs\[6\] _1762_ VGND VGND VPWR VPWR _1796_
+ sky130_fd_sc_hd__nand2_1
XFILLER_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3566_ cordic_inst.cordic_inst.x\[13\] cordic_inst.cordic_inst.cos_out\[13\] net212
+ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
X_3497_ _1527_ _1719_ net179 VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__o21ai_1
X_2517_ _0596_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__or2_1
X_2448_ net245 _0725_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__nand2_1
X_2379_ net222 _0711_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__nand2_1
XFILLER_29_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4118_ net258 _2093_ cordic_inst.cordic_inst.sin_out\[11\] VGND VGND VPWR VPWR _2094_
+ sky130_fd_sc_hd__a21oi_1
X_4049_ cordic_inst.cordic_inst.sin_out\[1\] cordic_inst.cordic_inst.sin_out\[0\]
+ net261 VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3420_ net267 cordic_inst.cordic_inst.z\[25\] VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__xor2_1
X_3351_ _1579_ _1589_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__xor2_1
X_2302_ net264 net286 VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nand2_2
X_3282_ net237 net303 VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4805_ net391 _0532_ _0227_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2997_ _1189_ _1190_ _1192_ net272 VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__o31a_1
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4736_ net389 _0463_ _0158_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[29\] sky130_fd_sc_hd__dfrtp_1
X_4667_ net357 _0396_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[21\] sky130_fd_sc_hd__dfxtp_2
X_3618_ _1785_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__inv_2
X_4598_ net385 _0330_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3549_ cordic_inst.cordic_inst.x\[30\] cordic_inst.cordic_inst.cos_out\[30\] net207
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2920_ net269 _1212_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__a21o_1
XFILLER_16_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2851_ cordic_inst.cordic_inst.y\[3\] cordic_inst.cordic_inst.y\[4\] net311 VGND
+ VGND VPWR VPWR _1154_ sky130_fd_sc_hd__mux2_1
X_2782_ cordic_inst.cordic_inst.y\[27\] cordic_inst.cordic_inst.y\[28\] net304 VGND
+ VGND VPWR VPWR _1085_ sky130_fd_sc_hd__mux2_1
XFILLER_31_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4521_ net380 _0000_ _0087_ VGND VGND VPWR VPWR cordic_inst.state\[2\] sky130_fd_sc_hd__dfrtp_1
X_4452_ net325 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__inv_2
X_3403_ _1639_ _1641_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__nand2_1
X_4383_ net326 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
X_3334_ net280 _1499_ _1571_ _1572_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__a31o_1
X_3265_ net248 net206 VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__or2_1
X_3196_ _1271_ _1270_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__nand2b_1
XFILLER_27_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4719_ net360 _0446_ _0141_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3050_ cordic_inst.cordic_inst.x\[19\] _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__nor2_1
XFILLER_35_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3952_ axi_controller.write_addr_reg\[1\] net47 net187 VGND VGND VPWR VPWR _0300_
+ sky130_fd_sc_hd__mux2_1
X_3883_ axi_controller.reg_input_data\[8\] _1964_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__or2_1
X_2903_ net246 _1130_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__nand2_1
X_2834_ _1079_ _1133_ _1135_ _1132_ net239 net233 VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__mux4_2
X_2765_ net263 net274 VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__and2_1
X_4504_ net345 VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__inv_2
X_2696_ _0842_ _1022_ _0841_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__a21bo_1
X_4435_ net338 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__inv_2
X_4366_ net336 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
X_3317_ _1554_ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__or2_1
X_4297_ axi_controller.reg_input_data\[20\] _2242_ VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__or2_1
X_3248_ net268 _0708_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__xnor2_1
X_3179_ cordic_inst.cordic_inst.x\[8\] net158 _1458_ net178 VGND VGND VPWR VPWR _0506_
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2550_ _0599_ _0882_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__nor2_1
Xoutput129 net129 VGND VGND VPWR VPWR rdata[25] sky130_fd_sc_hd__buf_2
X_2481_ _0644_ _0805_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__xnor2_1
Xoutput118 net118 VGND VGND VPWR VPWR rdata[15] sky130_fd_sc_hd__buf_2
X_4220_ cordic_inst.cordic_inst.cos_out\[22\] _2173_ net224 VGND VGND VPWR VPWR _2184_
+ sky130_fd_sc_hd__o21a_1
XFILLER_5_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4151_ cordic_inst.cordic_inst.sin_out\[14\] cordic_inst.cordic_inst.sin_out\[13\]
+ _2107_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__or3_1
X_4082_ net228 _2059_ _2061_ _2062_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__a22o_1
X_3102_ _1002_ _1404_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__xor2_1
X_3033_ _1210_ _1219_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_34_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3935_ axi_controller.read_addr_reg\[3\] axi_controller.read_addr_reg\[4\] axi_controller.read_addr_reg\[5\]
+ _1977_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__and4bb_1
XFILLER_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3866_ axi_controller.write_addr_reg\[2\] axi_controller.write_addr_reg\[7\] axi_controller.write_addr_reg\[6\]
+ axi_controller.write_addr_reg\[9\] VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__or4_1
X_3797_ axi_controller.reg_input_data\[24\] _1893_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__xnor2_1
X_2817_ cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.y\[6\] net308 VGND
+ VGND VPWR VPWR _1120_ sky130_fd_sc_hd__mux2_1
X_2748_ _0873_ _0914_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nand2b_1
X_4418_ net322 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__inv_2
X_2679_ _0976_ _0979_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__or2_1
Xfanout323 net328 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_4
Xfanout301 cordic_inst.cordic_inst.i\[1\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_2
Xfanout312 cordic_inst.cordic_inst.i\[0\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__buf_2
Xfanout334 net335 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_4
Xfanout356 net361 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlymetal6s2s_1
X_4349_ net321 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
Xfanout345 axi_controller.rst VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_2
Xfanout378 net388 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_2
Xfanout389 net390 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_2
Xfanout367 net371 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_2
XFILLER_27_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3720_ cordic_inst.deg_handler_inst.theta_norm\[16\] _1840_ VGND VGND VPWR VPWR _0015_
+ sky130_fd_sc_hd__xnor2_1
X_3651_ cordic_inst.deg_handler_inst.theta_abs\[14\] _1770_ VGND VGND VPWR VPWR _1804_
+ sky130_fd_sc_hd__nand2_1
X_3582_ net282 net180 _1580_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__and3_1
X_2602_ net154 _0758_ _0765_ net250 VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__a31o_1
X_2533_ _0858_ _0861_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__and2b_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2464_ _0789_ _0791_ _0793_ net271 VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__o31ai_1
X_4203_ cordic_inst.cordic_inst.sin_out\[20\] cordic_inst.cordic_inst.sin_out\[19\]
+ _2151_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__or3_1
X_2395_ cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.x\[6\] cordic_inst.cordic_inst.x\[7\]
+ cordic_inst.cordic_inst.x\[8\] net308 net297 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__mux4_1
X_4134_ net260 _2107_ cordic_inst.cordic_inst.sin_out\[13\] VGND VGND VPWR VPWR _2108_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_28_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4065_ cordic_inst.cordic_inst.cos_out\[3\] cordic_inst.cordic_inst.cos_out\[2\]
+ cordic_inst.cordic_inst.cos_out\[1\] cordic_inst.cordic_inst.cos_out\[0\] VGND VGND
+ VPWR VPWR _2048_ sky130_fd_sc_hd__or4_4
X_3016_ _1180_ _1185_ net272 VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4898_ net373 _0051_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3918_ axi_controller.read_addr_reg\[19\] net12 net197 VGND VGND VPWR VPWR _0285_
+ sky130_fd_sc_hd__mux2_1
X_3849_ net63 net62 net61 VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__nand3b_1
XFILLER_22_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout153 _1781_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xfanout164 _0629_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout186 _0626_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_2
Xfanout197 net199 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4821_ net403 _0548_ _0243_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[18\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_44_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4752_ net406 _0479_ _0174_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_4683_ net399 _0410_ _0105_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3703_ net252 _1829_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__nand2_1
X_3634_ _1762_ net147 _1795_ net150 cordic_inst.deg_handler_inst.theta_abs\[5\] VGND
+ VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a32o_1
X_3565_ cordic_inst.cordic_inst.x\[14\] cordic_inst.cordic_inst.cos_out\[14\] net212
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
X_3496_ _1518_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__nor2_1
X_2516_ _0667_ _0845_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__xor2_1
X_2447_ _0771_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nor2_1
X_2378_ net232 net222 VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_3_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4117_ cordic_inst.cordic_inst.sin_out\[10\] _2086_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__or2_1
X_4048_ axi_controller.result_out\[1\] _2033_ net202 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3350_ net267 _1582_ _1588_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__a21boi_1
X_2301_ net233 _0634_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a21oi_1
X_3281_ _1518_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__or2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4804_ net391 _0531_ _0226_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[1\] sky130_fd_sc_hd__dfrtp_2
X_4735_ net376 _0462_ _0157_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[28\] sky130_fd_sc_hd__dfrtp_1
X_2996_ _1297_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__and2b_1
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4666_ net351 _0395_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[20\] sky130_fd_sc_hd__dfxtp_2
X_3617_ cordic_inst.deg_handler_inst.theta_abs\[23\] _1784_ _1779_ VGND VGND VPWR
+ VPWR _1785_ sky130_fd_sc_hd__a21o_1
X_4597_ net382 _0329_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[30\] sky130_fd_sc_hd__dfxtp_1
X_3548_ net265 cordic_inst.cordic_inst.cos_out\[31\] net207 VGND VGND VPWR VPWR _0433_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3479_ _1632_ _1647_ _1705_ _1641_ _1645_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__o311a_1
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2850_ net283 _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__and2_1
XFILLER_31_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2781_ cordic_inst.cordic_inst.y\[23\] cordic_inst.cordic_inst.y\[24\] cordic_inst.cordic_inst.y\[25\]
+ cordic_inst.cordic_inst.y\[26\] net307 net301 VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__mux4_1
X_4520_ net380 _0007_ _0086_ VGND VGND VPWR VPWR cordic_inst.state\[1\] sky130_fd_sc_hd__dfrtp_1
X_4451_ net326 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__inv_2
X_3402_ cordic_inst.cordic_inst.z\[18\] _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__xor2_1
X_4382_ net326 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
X_3333_ net241 net294 net302 net288 VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3264_ net280 net206 _1501_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__a21oi_1
X_3195_ cordic_inst.cordic_inst.x\[2\] net158 _1468_ net176 VGND VGND VPWR VPWR _0500_
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2979_ _1254_ _1258_ _1278_ _1252_ _1249_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__a311o_2
X_4718_ net360 _0445_ _0140_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4649_ net384 _0380_ net326 VGND VGND VPWR VPWR axi_controller.result_out\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3951_ axi_controller.write_addr_reg\[0\] net36 net187 VGND VGND VPWR VPWR _0299_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2902_ net244 _1163_ _1202_ _1203_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a211o_1
X_3882_ net104 _1963_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__nand2_2
X_2833_ _1079_ _1135_ net233 VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__mux2_1
X_2764_ _0600_ _1067_ _1066_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux2_1
X_4503_ net340 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__inv_2
X_2695_ _0835_ _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__nand2_1
X_4434_ net337 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__inv_2
X_4365_ net336 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
X_3316_ cordic_inst.cordic_inst.z\[7\] _1553_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__nor2_1
X_4296_ net81 _2243_ _2247_ net347 VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_16_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3247_ _1484_ _1485_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__or2_1
X_3178_ _1290_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput108 net108 VGND VGND VPWR VPWR arready sky130_fd_sc_hd__buf_2
X_2480_ cordic_inst.cordic_inst.y\[29\] _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__nor2_1
Xoutput119 net119 VGND VGND VPWR VPWR rdata[16] sky130_fd_sc_hd__buf_2
X_4150_ cordic_inst.cordic_inst.cos_out\[15\] net226 _2120_ net315 VGND VGND VPWR
+ VPWR _2122_ sky130_fd_sc_hd__a31o_1
X_3101_ _1077_ _1226_ _1227_ net269 VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__o31a_1
X_4081_ cordic_inst.cordic_inst.sin_out\[6\] _2060_ net228 VGND VGND VPWR VPWR _2062_
+ sky130_fd_sc_hd__a21oi_1
X_3032_ cordic_inst.cordic_inst.x\[23\] _1334_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3934_ axi_controller.read_addr_reg\[1\] axi_controller.read_addr_reg\[0\] axi_controller.read_addr_reg\[7\]
+ axi_controller.read_addr_reg\[6\] VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__nor4_1
X_3865_ _1944_ _1945_ _1946_ _1947_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__or4_1
XFILLER_32_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2816_ _1117_ _1118_ net290 VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__mux2_1
X_3796_ axi_controller.reg_input_data\[23\] _1890_ _1874_ VGND VGND VPWR VPWR _1896_
+ sky130_fd_sc_hd__o21ba_1
X_2747_ _0873_ _0874_ _0878_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__o211ai_1
X_2678_ net182 _0997_ _1009_ net163 cordic_inst.cordic_inst.y\[28\] VGND VGND VPWR
+ VPWR _0558_ sky130_fd_sc_hd__a32o_1
X_4417_ net322 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
Xfanout313 axi_controller.mode VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_4
Xfanout302 net303 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_2
Xfanout357 net361 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_2
Xfanout346 net348 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__buf_2
Xfanout335 net339 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_2
Xfanout324 net325 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_4
X_4348_ net318 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
Xfanout379 net383 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_2
Xfanout368 net370 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_2
X_4279_ net200 _2235_ _2230_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_1_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3650_ _1770_ net147 _1803_ net151 cordic_inst.deg_handler_inst.theta_abs\[13\] VGND
+ VGND VPWR VPWR _0057_ sky130_fd_sc_hd__a32o_1
X_2601_ _0926_ _0930_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__nand3b_1
X_3581_ cordic_inst.cordic_inst.start cordic_inst.state\[2\] _0620_ _0618_ VGND VGND
+ VPWR VPWR _0400_ sky130_fd_sc_hd__o211a_1
X_2532_ _0844_ _0864_ _0865_ _0832_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__o221a_1
X_2463_ net279 _0766_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nor2_1
X_4202_ cordic_inst.cordic_inst.cos_out\[21\] net227 _2166_ net316 VGND VGND VPWR
+ VPWR _2168_ sky130_fd_sc_hd__a31oi_1
X_2394_ cordic_inst.cordic_inst.x\[5\] cordic_inst.cordic_inst.x\[6\] net307 VGND
+ VGND VPWR VPWR _0729_ sky130_fd_sc_hd__mux2_1
X_4133_ cordic_inst.cordic_inst.sin_out\[12\] _2099_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__or2_1
X_4064_ net259 _2045_ cordic_inst.cordic_inst.sin_out\[4\] VGND VGND VPWR VPWR _2047_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_39_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3015_ _1316_ _1317_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__nand2b_1
X_4897_ net372 _0050_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_3917_ axi_controller.read_addr_reg\[18\] net11 net196 VGND VGND VPWR VPWR _0284_
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3848_ net349 _1931_ _1930_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a21o_1
X_3779_ axi_controller.reg_input_data\[20\] _1882_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout165 net169 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_4
Xfanout187 _1929_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_4
Xfanout176 net178 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_4
Xfanout198 net199 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4820_ net404 _0547_ _0242_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[17\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_44_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ net400 _0478_ _0173_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4682_ net399 _0409_ _0104_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3702_ cordic_inst.deg_handler_inst.theta_norm\[9\] _1827_ VGND VGND VPWR VPWR _1829_
+ sky130_fd_sc_hd__or2_1
X_3633_ cordic_inst.deg_handler_inst.theta_abs\[5\] _1761_ VGND VGND VPWR VPWR _1795_
+ sky130_fd_sc_hd__nand2_1
X_3564_ cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.cos_out\[15\] net212
+ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
X_3495_ _1520_ _1717_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__nor2_1
X_2515_ _0849_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__inv_2
X_2446_ _0672_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__nand2_1
X_4116_ net203 _2092_ _2085_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__a21oi_1
X_2377_ net294 net302 VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4047_ _2030_ _2032_ net230 VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__mux2_1
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4949_ net407 _0578_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3280_ cordic_inst.cordic_inst.z\[14\] _1517_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__nor2_1
X_2300_ net264 net291 VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4803_ net389 _0530_ _0225_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.y\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4734_ net376 _0461_ _0156_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[27\] sky130_fd_sc_hd__dfrtp_1
X_2995_ cordic_inst.cordic_inst.x\[15\] _1296_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__nand2_1
X_4665_ net352 _0394_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[19\] sky130_fd_sc_hd__dfxtp_2
X_3616_ _1782_ _1783_ _0617_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__o21ai_1
X_4596_ net381 _0328_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[29\] sky130_fd_sc_hd__dfxtp_1
X_3547_ cordic_inst.cordic_inst.angle\[0\] net171 net159 cordic_inst.cordic_inst.z\[0\]
+ _1754_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3478_ _1629_ _1634_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__and2_1
X_2429_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2780_ cordic_inst.cordic_inst.y\[25\] cordic_inst.cordic_inst.y\[26\] net304 VGND
+ VGND VPWR VPWR _1083_ sky130_fd_sc_hd__mux2_1
X_4450_ net325 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__inv_2
X_3401_ net249 _1508_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__xnor2_1
X_4381_ net331 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
X_3332_ net302 _0705_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__nor2_1
X_3263_ net288 net294 net302 VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__nor3_1
X_3194_ _1274_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__and2_1
XFILLER_38_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2978_ _1254_ _1258_ _1278_ _1252_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__a31o_1
X_4717_ net359 _0444_ _0139_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4648_ net393 _0379_ net326 VGND VGND VPWR VPWR axi_controller.result_out\[25\] sky130_fd_sc_hd__dfrtp_1
X_4579_ net369 _0311_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3950_ axi_controller.done _1992_ net349 _0085_ _1918_ VGND VGND VPWR VPWR _0298_
+ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_18_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2901_ net244 _1163_ net215 VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__a21o_1
XFILLER_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3881_ net104 _1963_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__and2_1
X_2832_ cordic_inst.cordic_inst.y\[24\] cordic_inst.cordic_inst.y\[25\] cordic_inst.cordic_inst.y\[26\]
+ cordic_inst.cordic_inst.y\[27\] net304 net295 VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__mux4_1
XFILLER_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2763_ _0600_ net173 VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nor2_1
X_4502_ net340 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__inv_2
XFILLER_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2694_ _0864_ _0973_ _0837_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a21o_1
X_4433_ net337 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__inv_2
X_4364_ net334 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
X_4295_ axi_controller.reg_input_data\[19\] _2242_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__or2_1
X_3315_ cordic_inst.cordic_inst.z\[7\] _1553_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__and2_1
X_3246_ _1481_ _1483_ cordic_inst.cordic_inst.z\[21\] VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__a21oi_1
X_3177_ _1284_ _1289_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__nand2_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput109 net109 VGND VGND VPWR VPWR awready sky130_fd_sc_hd__buf_2
XFILLER_5_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3100_ _1236_ _1238_ _1401_ _1234_ _1231_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__a311oi_1
X_4080_ cordic_inst.cordic_inst.sin_out\[6\] _2060_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__or2_1
X_3031_ _1220_ _1333_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3933_ _1974_ _1975_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__nor2_1
X_3864_ axi_controller.write_addr_reg\[24\] axi_controller.write_addr_reg\[27\] axi_controller.write_addr_reg\[26\]
+ axi_controller.write_addr_reg\[28\] VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__or4b_1
X_2815_ cordic_inst.cordic_inst.y\[17\] cordic_inst.cordic_inst.y\[18\] cordic_inst.cordic_inst.y\[19\]
+ cordic_inst.cordic_inst.y\[20\] net311 net300 VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__mux4_1
X_3795_ _1891_ _1895_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__xnor2_1
X_2746_ _0876_ _0879_ _0913_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__or3b_1
X_2677_ _0821_ _0996_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__nand2_1
X_4416_ net321 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__inv_2
Xfanout314 axi_controller.mode VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_4
Xfanout303 cordic_inst.cordic_inst.i\[0\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_2
Xfanout347 net348 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__buf_2
Xfanout336 net339 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_4
X_4347_ net318 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
Xfanout325 net328 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net370 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_1
Xfanout358 net361 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_2
X_4278_ net313 _2231_ _2232_ _2233_ _2234_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__o32a_1
X_3229_ cordic_inst.cordic_inst.y\[4\] cordic_inst.cordic_inst.sin_out\[4\] net211
+ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux2_1
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3580_ cordic_inst.cordic_inst.done cordic_inst.cordic_inst.state\[0\] cordic_inst.cordic_inst.state\[1\]
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o21a_1
X_2600_ _0933_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__nor2_1
X_2531_ _0823_ _0828_ _0829_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a21o_1
X_4201_ net227 _2166_ cordic_inst.cordic_inst.cos_out\[21\] VGND VGND VPWR VPWR _2167_
+ sky130_fd_sc_hd__a21o_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2462_ net242 _0676_ net170 VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__a21o_1
X_2393_ _0726_ _0727_ net290 VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__mux2_1
X_4132_ _2102_ _2106_ axi_controller.result_out\[12\] net203 VGND VGND VPWR VPWR _0366_
+ sky130_fd_sc_hd__o2bb2a_1
X_4063_ cordic_inst.cordic_inst.sin_out\[4\] net259 _2045_ VGND VGND VPWR VPWR _2046_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3014_ cordic_inst.cordic_inst.x\[11\] _1315_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__nand2_1
X_4965_ net380 _0594_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_1
X_3916_ axi_controller.read_addr_reg\[17\] net10 net197 VGND VGND VPWR VPWR _0283_
+ sky130_fd_sc_hd__mux2_1
X_4896_ net372 _0049_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_3847_ axi_controller.state\[0\] net68 net107 _1920_ axi_controller.state\[2\] VGND
+ VGND VPWR VPWR _1931_ sky130_fd_sc_hd__a32o_1
X_3778_ _1874_ _1880_ axi_controller.reg_input_data\[19\] VGND VGND VPWR VPWR _1882_
+ sky130_fd_sc_hd__mux2_1
X_2729_ net184 _1043_ _1046_ net166 cordic_inst.cordic_inst.y\[14\] VGND VGND VPWR
+ VPWR _0544_ sky130_fd_sc_hd__a32o_1
Xfanout155 net156 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_2
Xfanout188 _1929_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
Xfanout177 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_4
Xfanout166 net167 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
Xfanout199 _1926_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ net400 _0477_ _0172_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.sin_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_4681_ net399 _0408_ _0103_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3701_ cordic_inst.deg_handler_inst.theta_norm\[9\] _1828_ VGND VGND VPWR VPWR _0039_
+ sky130_fd_sc_hd__xnor2_1
X_3632_ _1761_ net148 _1794_ net150 cordic_inst.deg_handler_inst.theta_abs\[4\] VGND
+ VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a32o_1
X_3563_ cordic_inst.cordic_inst.x\[16\] cordic_inst.cordic_inst.cos_out\[16\] net212
+ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3494_ _1515_ _1627_ _1530_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__a21o_1
X_2514_ cordic_inst.cordic_inst.y\[19\] _0847_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__xor2_1
X_2445_ _0776_ _0777_ _0779_ _0773_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__o211a_1
X_4115_ net228 _2087_ _2088_ _2090_ _2091_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__o32a_1
X_2376_ net295 net305 VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nor2_2
X_4046_ cordic_inst.cordic_inst.cos_out\[1\] _2031_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4948_ net407 _0577_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_1
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4879_ net356 axi_controller.reg_input_data\[11\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2994_ cordic_inst.cordic_inst.x\[15\] _1296_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__nor2_1
X_4802_ net383 _0529_ _0224_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4733_ net375 _0460_ _0155_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[26\] sky130_fd_sc_hd__dfrtp_1
X_4664_ net352 _0393_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[18\] sky130_fd_sc_hd__dfxtp_1
X_4595_ net381 _0327_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[28\] sky130_fd_sc_hd__dfxtp_1
X_3615_ cordic_inst.deg_handler_inst.theta_abs\[20\] cordic_inst.deg_handler_inst.theta_abs\[21\]
+ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__nand2_1
X_3546_ _1597_ _1753_ net182 VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__o21a_1
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3477_ _1703_ _1704_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__nand2_1
X_2428_ _0760_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__or2_1
X_2359_ cordic_inst.cordic_inst.x\[16\] cordic_inst.cordic_inst.x\[17\] cordic_inst.cordic_inst.x\[18\]
+ cordic_inst.cordic_inst.x\[19\] net310 net299 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_27_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4029_ axi_controller.reg_input_data\[2\] _2018_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3400_ _1637_ _1638_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__and2_1
X_4380_ net331 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
X_3331_ _1568_ _1569_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__nor2_1
X_3262_ _1499_ _1500_ net281 VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__a21oi_1
X_3193_ _1269_ _1272_ _1273_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__nand3_1
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2977_ _1252_ _1253_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__or2_1
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4716_ net367 _0443_ _0138_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4647_ net393 _0378_ net326 VGND VGND VPWR VPWR axi_controller.result_out\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4578_ net363 _0310_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3529_ cordic_inst.cordic_inst.angle\[6\] net171 net160 cordic_inst.cordic_inst.z\[6\]
+ _1742_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a221o_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2900_ net276 _1168_ _1069_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__o21ai_2
X_3880_ _0622_ _1962_ _1943_ _1922_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__and4bb_4
X_2831_ _1132_ _1133_ net291 VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__mux2_1
X_2762_ net183 _0718_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__nand2_1
XFILLER_8_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ net341 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__inv_2
X_4432_ net337 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__inv_2
X_2693_ cordic_inst.cordic_inst.y\[24\] net169 _1019_ _1020_ VGND VGND VPWR VPWR _0554_
+ sky130_fd_sc_hd__a22o_1
X_4363_ net334 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
X_4294_ net80 _2243_ _2246_ net347 VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__o211a_1
X_3314_ net266 _1481_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__mux2_1
X_3245_ cordic_inst.cordic_inst.z\[21\] _1481_ _1483_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__and3_1
X_3176_ cordic_inst.cordic_inst.x\[9\] net158 _1455_ _1456_ VGND VGND VPWR VPWR _0507_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_37_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3030_ _1068_ _1090_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__or2_1
XFILLER_17_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3932_ axi_controller.read_addr_reg\[9\] axi_controller.read_addr_reg\[8\] axi_controller.read_addr_reg\[11\]
+ axi_controller.read_addr_reg\[10\] VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__or4_1
X_3863_ axi_controller.write_addr_reg\[29\] axi_controller.write_addr_reg\[30\] axi_controller.write_addr_reg\[31\]
+ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__nand3_1
X_2814_ cordic_inst.cordic_inst.y\[13\] cordic_inst.cordic_inst.y\[14\] cordic_inst.cordic_inst.y\[15\]
+ cordic_inst.cordic_inst.y\[16\] net310 net299 VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__mux4_1
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3794_ axi_controller.reg_input_data\[23\] _1880_ _1894_ VGND VGND VPWR VPWR _1895_
+ sky130_fd_sc_hd__a21oi_1
X_2745_ net185 _1037_ _1056_ net166 cordic_inst.cordic_inst.y\[8\] VGND VGND VPWR
+ VPWR _0538_ sky130_fd_sc_hd__a32o_1
X_2676_ cordic_inst.cordic_inst.y\[29\] net163 _1008_ net182 VGND VGND VPWR VPWR _0559_
+ sky130_fd_sc_hd__a22o_1
X_4415_ net321 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
Xfanout304 net305 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_4
X_4346_ net255 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
Xfanout348 net34 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_2
Xfanout337 net338 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_4
Xfanout326 net327 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__buf_4
Xfanout315 net316 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_2
Xfanout359 net360 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_2
X_4277_ cordic_inst.cordic_inst.sin_out\[30\] net256 _2224_ net231 VGND VGND VPWR
+ VPWR _2234_ sky130_fd_sc_hd__a31o_1
X_3228_ cordic_inst.cordic_inst.y\[5\] cordic_inst.cordic_inst.sin_out\[5\] net211
+ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
XFILLER_27_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3159_ _1302_ _1445_ _1299_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ _0835_ _0841_ _0842_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__a21bo_1
X_2461_ _0637_ _0761_ net279 VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__a21oi_1
X_4200_ cordic_inst.cordic_inst.cos_out\[20\] cordic_inst.cordic_inst.cos_out\[19\]
+ _2155_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__or3_1
X_2392_ cordic_inst.cordic_inst.x\[13\] cordic_inst.cordic_inst.x\[14\] cordic_inst.cordic_inst.x\[15\]
+ cordic_inst.cordic_inst.x\[16\] net310 net300 VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__mux4_2
X_4131_ _2104_ _2105_ net203 VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__o21a_1
X_4062_ cordic_inst.cordic_inst.sin_out\[3\] cordic_inst.cordic_inst.sin_out\[2\]
+ cordic_inst.cordic_inst.sin_out\[1\] cordic_inst.cordic_inst.sin_out\[0\] VGND VGND
+ VPWR VPWR _2045_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_39_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3013_ cordic_inst.cordic_inst.x\[11\] _1315_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nor2_1
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4964_ net399 _0593_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_1
X_3915_ axi_controller.read_addr_reg\[16\] net9 net197 VGND VGND VPWR VPWR _0282_
+ sky130_fd_sc_hd__mux2_1
X_4895_ net373 _0048_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3846_ net349 net107 axi_controller.state\[3\] VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__and3_1
X_3777_ axi_controller.reg_input_data\[19\] _1881_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__xor2_1
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2728_ _0925_ _1042_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__nand2_1
X_2659_ _0984_ _0986_ _0989_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__nand4_1
X_4329_ net117 net192 net156 axi_controller.result_out\[14\] VGND VGND VPWR VPWR _0580_
+ sky130_fd_sc_hd__a22o_1
Xfanout156 _2256_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_2
Xfanout189 net190 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_4
Xfanout178 _0627_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_2
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XFILLER_43_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3700_ net252 _1827_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__nand2_1
X_4680_ net396 _0407_ _0102_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.cos_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3631_ cordic_inst.deg_handler_inst.theta_abs\[4\] _1760_ VGND VGND VPWR VPWR _1794_
+ sky130_fd_sc_hd__nand2_1
X_3562_ cordic_inst.cordic_inst.x\[17\] cordic_inst.cordic_inst.cos_out\[17\] net212
+ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
X_2513_ cordic_inst.cordic_inst.y\[19\] _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nor2_1
X_3493_ cordic_inst.cordic_inst.angle\[16\] net172 net159 cordic_inst.cordic_inst.z\[16\]
+ _1716_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a221o_1
X_2444_ _0601_ _0636_ _0691_ _0686_ net240 net244 VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__mux4_2
X_2375_ cordic_inst.cordic_inst.x\[2\] cordic_inst.cordic_inst.x\[3\] net312 VGND
+ VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux2_1
X_4114_ cordic_inst.cordic_inst.cos_out\[10\] net225 _2089_ net314 VGND VGND VPWR
+ VPWR _2091_ sky130_fd_sc_hd__a31o_1
X_4045_ cordic_inst.cordic_inst.cos_out\[0\] net223 VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__nand2_1
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4947_ net407 _0576_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_1
X_4878_ net356 axi_controller.reg_input_data\[10\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3829_ cordic_inst.sign_handler_inst.done_d cordic_inst.cordic_inst.done VGND VGND
+ VPWR VPWR cordic_inst.sign_handler_inst.done_pulse sky130_fd_sc_hd__and2b_1
XFILLER_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2993_ _1198_ _1216_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__xnor2_1
X_4801_ net383 _0528_ _0223_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[30\] sky130_fd_sc_hd__dfrtp_4
X_4732_ net375 _0459_ _0154_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4663_ net352 _0392_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[17\] sky130_fd_sc_hd__dfxtp_1
X_3614_ cordic_inst.deg_handler_inst.theta_abs\[18\] cordic_inst.deg_handler_inst.theta_abs\[19\]
+ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__nor2_1
X_4594_ net385 _0326_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[27\] sky130_fd_sc_hd__dfxtp_1
X_3545_ cordic_inst.cordic_inst.z\[0\] _1583_ _1584_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__and3_1
X_3476_ cordic_inst.cordic_inst.angle\[20\] net173 net161 cordic_inst.cordic_inst.z\[20\]
+ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__a22oi_1
X_2427_ net264 _0721_ _0724_ _0728_ net244 _0607_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__mux4_1
X_2358_ net247 _0692_ _0689_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o21ai_2
XFILLER_28_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2289_ axi_controller.read_addr_reg\[31\] VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__inv_2
XFILLER_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4028_ net82 _2019_ _2021_ net349 VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__o211a_1
XFILLER_25_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3330_ cordic_inst.cordic_inst.z\[5\] _1567_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__nor2_1
X_3261_ net294 net303 VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__nand2_1
X_3192_ net183 _1277_ _1466_ net165 cordic_inst.cordic_inst.x\[3\] VGND VGND VPWR
+ VPWR _0501_ sky130_fd_sc_hd__a32o_1
XFILLER_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2976_ _1258_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__nand2_1
X_4715_ net367 _0442_ _0137_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4646_ net392 _0377_ net331 VGND VGND VPWR VPWR axi_controller.result_out\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4577_ net363 _0309_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3528_ _1563_ _1607_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__a21oi_1
X_3459_ cordic_inst.cordic_inst.angle\[24\] net173 net161 cordic_inst.cordic_inst.z\[24\]
+ _1690_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__a221o_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2830_ cordic_inst.cordic_inst.y\[20\] cordic_inst.cordic_inst.y\[21\] cordic_inst.cordic_inst.y\[22\]
+ cordic_inst.cordic_inst.y\[23\] net307 net301 VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__mux4_1
X_2761_ net183 _0898_ _1065_ net165 cordic_inst.cordic_inst.y\[1\] VGND VGND VPWR
+ VPWR _0531_ sky130_fd_sc_hd__a32o_1
X_4500_ net342 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__inv_2
X_2692_ net177 _0979_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__nor2_1
XFILLER_8_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4431_ net337 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__inv_2
XANTENNA_1 _2028_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4362_ net335 VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
X_4293_ axi_controller.reg_input_data\[18\] _2242_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__or2_1
X_3313_ net281 _0707_ _1521_ _1510_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__a31o_1
X_3244_ _1482_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__inv_2
XFILLER_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3175_ _1295_ _1439_ net178 VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__a21o_1
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2959_ _1169_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__xor2_1
XFILLER_22_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4629_ net398 _0360_ net336 VGND VGND VPWR VPWR axi_controller.result_out\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3931_ axi_controller.read_addr_reg\[13\] axi_controller.read_addr_reg\[12\] axi_controller.read_addr_reg\[15\]
+ axi_controller.read_addr_reg\[14\] VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3862_ axi_controller.write_addr_reg\[16\] axi_controller.write_addr_reg\[19\] axi_controller.write_addr_reg\[18\]
+ axi_controller.write_addr_reg\[21\] VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__or4_1
X_2813_ net243 _1115_ _1110_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__o21ai_2
X_3793_ axi_controller.reg_input_data\[23\] _1892_ _1893_ VGND VGND VPWR VPWR _1894_
+ sky130_fd_sc_hd__o21a_1
X_2744_ _0915_ _0959_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nand2_1
X_2675_ _0998_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__xnor2_1
X_4414_ net321 VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__inv_2
X_4345_ cordic_inst.deg_handler_inst.theta_abs\[31\] VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
Xfanout305 net306 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_2
Xfanout316 axi_controller.mode VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_4
Xfanout327 net328 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__buf_2
Xfanout338 net339 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_4
X_4276_ net256 _2224_ cordic_inst.cordic_inst.sin_out\[30\] VGND VGND VPWR VPWR _2233_
+ sky130_fd_sc_hd__a21oi_1
Xfanout349 net34 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__buf_2
X_3227_ cordic_inst.cordic_inst.y\[6\] cordic_inst.cordic_inst.sin_out\[6\] net211
+ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux2_1
X_3158_ _1303_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nand2_1
X_3089_ _1222_ _1391_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2460_ net246 _0759_ net170 VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21o_1
X_2391_ cordic_inst.cordic_inst.x\[9\] cordic_inst.cordic_inst.x\[10\] cordic_inst.cordic_inst.x\[11\]
+ cordic_inst.cordic_inst.x\[12\] net309 net298 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__mux4_1
X_4130_ cordic_inst.cordic_inst.cos_out\[12\] net225 _2103_ net314 VGND VGND VPWR
+ VPWR _2105_ sky130_fd_sc_hd__a31o_1
X_4061_ axi_controller.result_out\[4\] net202 VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__nor2_1
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3012_ _1098_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4963_ net398 _0592_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3914_ axi_controller.read_addr_reg\[15\] net8 net196 VGND VGND VPWR VPWR _0281_
+ sky130_fd_sc_hd__mux2_1
X_4894_ net373 _0047_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_3845_ net349 _0622_ axi_controller.state\[3\] net188 VGND VGND VPWR VPWR _0004_
+ sky130_fd_sc_hd__a31o_1
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3776_ _1874_ _1880_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__nand2_1
X_2727_ cordic_inst.cordic_inst.y\[15\] net166 _1045_ net184 VGND VGND VPWR VPWR _0545_
+ sky130_fd_sc_hd__a22o_1
X_2658_ cordic_inst.cordic_inst.y\[25\] _0988_ _0976_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a21o_1
X_2589_ cordic_inst.cordic_inst.y\[14\] _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__nand2_1
X_4328_ net118 net192 net156 axi_controller.result_out\[15\] VGND VGND VPWR VPWR _0579_
+ sky130_fd_sc_hd__a22o_1
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
Xfanout179 net182 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_2
X_4259_ cordic_inst.deg_handler_inst.kuadran\[0\] _2211_ VGND VGND VPWR VPWR _2218_
+ sky130_fd_sc_hd__nor2_1
Xfanout157 _2256_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_4
XFILLER_28_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3630_ _1760_ net148 _1793_ net150 cordic_inst.deg_handler_inst.theta_abs\[3\] VGND
+ VGND VPWR VPWR _0078_ sky130_fd_sc_hd__a32o_1
X_3561_ cordic_inst.cordic_inst.x\[18\] cordic_inst.cordic_inst.cos_out\[18\] net212
+ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
X_2512_ _0666_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__xnor2_1
X_3492_ _1629_ _1634_ _1715_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__o21a_1
X_2443_ _0776_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nor2_1
X_2374_ net283 net290 net301 VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__nor3b_1
X_4113_ net226 _2089_ cordic_inst.cordic_inst.cos_out\[10\] VGND VGND VPWR VPWR _2090_
+ sky130_fd_sc_hd__a21oi_1
X_4044_ cordic_inst.cordic_inst.sin_out\[1\] _2029_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4946_ net403 _0575_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_1
X_4877_ net356 axi_controller.reg_input_data\[9\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3828_ _0618_ _1918_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__nor2_1
X_3759_ axi_controller.reg_input_data\[11\] axi_controller.reg_input_data\[10\] axi_controller.reg_input_data\[9\]
+ axi_controller.reg_input_data\[8\] VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__or4_1
XFILLER_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4800_ net383 _0527_ _0222_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[29\] sky130_fd_sc_hd__dfrtp_4
X_2992_ _1293_ _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__nand2b_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4731_ net372 _0458_ _0153_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[24\] sky130_fd_sc_hd__dfrtp_1
X_4662_ net352 _0391_ VGND VGND VPWR VPWR axi_controller.reg_input_data\[16\] sky130_fd_sc_hd__dfxtp_1
X_3613_ cordic_inst.deg_handler_inst.theta_abs\[31\] _1780_ VGND VGND VPWR VPWR _1781_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4593_ net381 _0325_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[26\] sky130_fd_sc_hd__dfxtp_1
X_3544_ cordic_inst.cordic_inst.angle\[1\] net172 net160 cordic_inst.cordic_inst.z\[1\]
+ _1752_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__a221o_1
X_3475_ _1490_ _1650_ _1654_ _1702_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__a31o_1
X_2426_ net238 _0724_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nand2_1
X_2357_ net264 _0634_ _0657_ _0654_ net234 net240 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__mux4_2
X_2288_ axi_controller.state\[3\] VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__inv_2
X_4027_ axi_controller.reg_input_data\[1\] _2018_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__or2_1
XFILLER_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4929_ net375 _0029_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_8_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3260_ net288 net294 VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__nand2_1
X_3191_ _1266_ _1274_ _1276_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__nand3_1
XFILLER_35_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2975_ _1263_ _1277_ _1260_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a21o_1
X_4714_ net366 _0441_ _0136_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4645_ net394 _0376_ net331 VGND VGND VPWR VPWR axi_controller.result_out\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4576_ net364 _0308_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[9\] sky130_fd_sc_hd__dfxtp_1
X_3527_ net175 _1608_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__or2_1
X_3458_ _1689_ net180 _1658_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__and3b_1
X_3389_ _1625_ _1626_ _1529_ _1533_ _1535_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__a2111o_1
X_2409_ _0694_ _0701_ net235 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__mux2_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2760_ _0896_ _0897_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nand2_1
XFILLER_8_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2691_ _0974_ _0978_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__nand2_1
XANTENNA_2 net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4430_ net336 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__inv_2
X_4361_ net329 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
X_4292_ net79 _2243_ _2245_ net346 VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o211a_1
X_3312_ _1550_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__inv_2
X_3243_ net268 _0714_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__nor2_1
X_3174_ _1295_ _1439_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__nor2_1
XFILLER_39_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ _1148_ _1157_ _1164_ net270 VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__o31a_1
X_4628_ net398 _0359_ net336 VGND VGND VPWR VPWR axi_controller.result_out\[5\] sky130_fd_sc_hd__dfrtp_1
X_2889_ net262 _1127_ _1129_ _1119_ net242 net239 VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__mux4_2
X_4559_ net355 _0291_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3930_ axi_controller.read_addr_reg\[31\] net26 net195 VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3861_ axi_controller.write_addr_reg\[20\] axi_controller.write_addr_reg\[23\] axi_controller.write_addr_reg\[22\]
+ axi_controller.write_addr_reg\[25\] VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__or4_1
X_3792_ axi_controller.reg_input_data\[23\] _1892_ _1880_ VGND VGND VPWR VPWR _1893_
+ sky130_fd_sc_hd__a21oi_1
X_2812_ net262 _1074_ _1113_ _1111_ net234 net238 VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__mux4_1
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2743_ net184 _1054_ _1055_ net166 cordic_inst.cordic_inst.y\[9\] VGND VGND VPWR
+ VPWR _0539_ sky130_fd_sc_hd__a32o_1
X_2674_ _0817_ _0997_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__and2b_1
X_4413_ net321 VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__inv_2
X_4344_ _2257_ net112 net194 VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux2_1
Xfanout339 net344 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_2
Xfanout306 cordic_inst.cordic_inst.i\[0\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout317 net319 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_4
Xfanout328 axi_controller.rst VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_4
X_4275_ net223 _2227_ cordic_inst.cordic_inst.cos_out\[30\] VGND VGND VPWR VPWR _2232_
+ sky130_fd_sc_hd__a21oi_1
X_3226_ cordic_inst.cordic_inst.y\[7\] cordic_inst.cordic_inst.sin_out\[7\] net210
+ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
X_3157_ _1326_ _1443_ _1307_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__o21a_1
X_3088_ net215 _1212_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__or2_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2390_ _0721_ _0724_ net285 VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__mux2_1
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4060_ axi_controller.result_out\[3\] _2043_ net202 VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3011_ _1180_ _1185_ _1187_ net272 VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o31a_1
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4962_ net398 _0591_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_1
X_4893_ net373 _0046_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_3913_ axi_controller.read_addr_reg\[14\] net7 net196 VGND VGND VPWR VPWR _0280_
+ sky130_fd_sc_hd__mux2_1
X_3844_ axi_controller.state\[0\] net349 net68 _0622_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__and4_1
X_3775_ axi_controller.reg_input_data\[31\] _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__nand2_2
X_2726_ _0920_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__xnor2_1
X_2657_ _0979_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__nand2_1
X_2588_ _0779_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__xor2_2
Xfanout147 net149 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
X_4327_ net119 net192 net156 axi_controller.result_out\[16\] VGND VGND VPWR VPWR _0578_
+ sky130_fd_sc_hd__a22o_1
X_4258_ axi_controller.result_out\[27\] net200 _2216_ _2217_ VGND VGND VPWR VPWR _0381_
+ sky130_fd_sc_hd__o22a_1
Xfanout169 _0629_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_2
Xfanout158 cordic_inst.cordic_inst.next_state\[1\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_4
X_3209_ cordic_inst.cordic_inst.y\[24\] cordic_inst.cordic_inst.sin_out\[24\] net208
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_1
X_4189_ cordic_inst.cordic_inst.cos_out\[19\] net227 _2155_ net314 VGND VGND VPWR
+ VPWR _2157_ sky130_fd_sc_hd__a31o_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3560_ cordic_inst.cordic_inst.x\[19\] cordic_inst.cordic_inst.cos_out\[19\] net212
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
XFILLER_6_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2511_ _0667_ _0787_ net273 VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o21a_1
XFILLER_6_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3491_ net175 _1705_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__nor2_1
X_2442_ net286 _0754_ _0637_ net274 VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__o211a_1
X_2373_ net282 net293 net295 net305 VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nor4b_1
X_4112_ cordic_inst.cordic_inst.cos_out\[9\] cordic_inst.cordic_inst.cos_out\[8\]
+ cordic_inst.cordic_inst.cos_out\[7\] _2068_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__or4_2
X_4043_ cordic_inst.cordic_inst.sin_out\[0\] net261 VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4945_ net403 _0574_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4876_ net356 axi_controller.reg_input_data\[8\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3827_ axi_controller.reg_done_flag axi_controller.start_pulse_reg VGND VGND VPWR
+ VPWR _1918_ sky130_fd_sc_hd__nand2b_1
X_3758_ cordic_inst.deg_handler_inst.theta_norm\[30\] cordic_inst.deg_handler_inst.theta_norm\[29\]
+ _1861_ net254 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and4bb_1
X_2709_ _0850_ _0852_ _1030_ net177 VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__a31o_1
X_3689_ cordic_inst.deg_handler_inst.theta_norm\[4\] _1819_ net252 VGND VGND VPWR
+ VPWR _1821_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2991_ _1292_ cordic_inst.cordic_inst.x\[9\] VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__nand2b_1
X_4730_ net376 _0457_ _0152_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[23\] sky130_fd_sc_hd__dfrtp_1
X_4661_ net389 cordic_inst.cordic_inst.done net322 VGND VGND VPWR VPWR cordic_inst.sign_handler_inst.done_d
+ sky130_fd_sc_hd__dfrtp_1
X_3612_ cordic_inst.deg_handler_inst.theta_abs\[22\] _1776_ _1779_ cordic_inst.deg_handler_inst.theta_abs\[23\]
+ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__a211oi_1
X_4592_ net381 _0324_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[25\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_24_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3543_ _1597_ _1598_ _1751_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__a21oi_1
X_3474_ net180 _1691_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__nand2_1
X_2425_ net264 _0696_ _0698_ _0702_ net244 net240 VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__mux4_2
X_2356_ net235 _0657_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__o21ai_1
X_2287_ axi_controller.write_addr_reg\[4\] VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__inv_2
X_4026_ net71 _2019_ _2020_ net349 VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_27_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4928_ net375 _0028_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4859_ net372 _0068_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3190_ cordic_inst.cordic_inst.x\[4\] net158 _1465_ net177 VGND VGND VPWR VPWR _0502_
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2974_ _1266_ _1274_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a21o_1
X_4713_ net367 _0440_ _0135_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4644_ net394 _0375_ net333 VGND VGND VPWR VPWR axi_controller.result_out\[21\] sky130_fd_sc_hd__dfrtp_1
X_4575_ net363 _0307_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3526_ cordic_inst.cordic_inst.angle\[7\] net171 net160 cordic_inst.cordic_inst.z\[7\]
+ _1740_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__a221o_1
X_3457_ _1480_ _1655_ _1657_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__and3_1
X_2408_ _0718_ _0735_ _0738_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nor4b_2
X_3388_ _1625_ _1626_ _1535_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__a21o_1
X_2339_ cordic_inst.cordic_inst.x\[14\] cordic_inst.cordic_inst.x\[15\] cordic_inst.cordic_inst.x\[16\]
+ cordic_inst.cordic_inst.x\[17\] net310 net299 VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4009_ axi_controller.reg_input_data\[25\] _2008_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__or2_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2690_ net186 _1017_ _1018_ net169 cordic_inst.cordic_inst.y\[25\] VGND VGND VPWR
+ VPWR _0555_ sky130_fd_sc_hd__a32o_1
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4360_ net329 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
X_3311_ cordic_inst.cordic_inst.z\[9\] _1549_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__or2_1
X_4291_ axi_controller.reg_input_data\[17\] _2242_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__or2_1
X_3242_ net268 _0714_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__nand2_2
XFILLER_39_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3173_ net185 _1441_ _1454_ net168 cordic_inst.cordic_inst.x\[10\] VGND VGND VPWR
+ VPWR _0508_ sky130_fd_sc_hd__a32o_1
XFILLER_23_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2957_ _1257_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__or2_1
XFILLER_41_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2888_ net241 _1129_ _1070_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__a21boi_1
X_4627_ net399 _0358_ net336 VGND VGND VPWR VPWR axi_controller.result_out\[4\] sky130_fd_sc_hd__dfrtp_1
X_4558_ net354 _0290_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[24\] sky130_fd_sc_hd__dfxtp_1
X_4489_ net330 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__inv_2
X_3509_ cordic_inst.cordic_inst.angle\[12\] net172 net159 cordic_inst.cordic_inst.z\[12\]
+ _1728_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a221o_1
XFILLER_17_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3860_ axi_controller.state\[0\] axi_controller.state\[3\] VGND VGND VPWR VPWR _1943_
+ sky130_fd_sc_hd__or2_1
X_3791_ axi_controller.reg_input_data\[22\] axi_controller.reg_input_data\[21\] _1883_
+ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__or3_1
X_2811_ _1111_ _1113_ net291 VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__mux2_1
X_2742_ _0957_ _1037_ _0955_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__a21o_1
X_4412_ net321 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__inv_2
X_2673_ net181 _1000_ _1006_ net164 cordic_inst.cordic_inst.y\[30\] VGND VGND VPWR
+ VPWR _0560_ sky130_fd_sc_hd__a32o_1
X_4343_ axi_controller.reg_done_flag _1990_ _2254_ axi_controller.result_out\[0\]
+ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__a22o_1
Xfanout329 net345 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_4
Xfanout307 net312 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_4
Xfanout318 net319 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_2
X_4274_ cordic_inst.cordic_inst.cos_out\[30\] net223 _2227_ VGND VGND VPWR VPWR _2231_
+ sky130_fd_sc_hd__and3_1
X_3225_ cordic_inst.cordic_inst.y\[8\] cordic_inst.cordic_inst.sin_out\[8\] net210
+ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
X_3156_ _1311_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__nor2_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3087_ _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__inv_2
XFILLER_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3989_ axi_controller.state\[0\] _1998_ _1996_ _1995_ VGND VGND VPWR VPWR _1999_
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3010_ _1304_ _1309_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4961_ net398 _0590_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4892_ net373 _0045_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_3912_ axi_controller.read_addr_reg\[13\] net6 net195 VGND VGND VPWR VPWR _0279_
+ sky130_fd_sc_hd__mux2_1
X_3843_ net199 _1928_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__or2_1
XFILLER_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3774_ _1876_ _1878_ axi_controller.reg_input_data\[24\] VGND VGND VPWR VPWR _1879_
+ sky130_fd_sc_hd__or3b_1
XFILLER_9_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2725_ cordic_inst.cordic_inst.y\[14\] _0923_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__a21bo_1
X_2656_ _0984_ _0986_ _0989_ _0990_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__and4_1
X_2587_ _0771_ _0772_ _0778_ net271 VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__o31ai_2
X_4326_ net120 net192 net156 axi_controller.result_out\[17\] VGND VGND VPWR VPWR _0577_
+ sky130_fd_sc_hd__a22o_1
Xfanout159 _0629_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
X_4257_ _2211_ _2212_ net200 VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__o21ai_1
X_4188_ net227 _2155_ cordic_inst.cordic_inst.cos_out\[19\] VGND VGND VPWR VPWR _2156_
+ sky130_fd_sc_hd__a21oi_1
X_3208_ cordic_inst.cordic_inst.y\[25\] cordic_inst.cordic_inst.sin_out\[25\] net209
+ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux2_1
X_3139_ _1332_ _1361_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__nand2_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3490_ net179 _1712_ _1713_ _1714_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__a31o_1
X_2510_ net271 _0787_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__nand2_1
X_2441_ net277 _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nor2_1
X_2372_ net294 net303 VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nand2b_2
X_4111_ net259 _2086_ cordic_inst.cordic_inst.sin_out\[10\] VGND VGND VPWR VPWR _2088_
+ sky130_fd_sc_hd__a21oi_1
X_4042_ axi_controller.result_out\[0\] _2028_ net200 VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4944_ net395 _0573_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4875_ net365 axi_controller.reg_input_data\[7\] VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_norm\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3826_ net274 _0614_ _1917_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.next_state\[0\]
+ sky130_fd_sc_hd__o21a_1
X_3757_ cordic_inst.deg_handler_inst.theta_norm\[30\] _1863_ VGND VGND VPWR VPWR _0031_
+ sky130_fd_sc_hd__xor2_1
X_2708_ _0852_ _1030_ _0850_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a21oi_1
X_3688_ cordic_inst.deg_handler_inst.theta_norm\[4\] _1820_ VGND VGND VPWR VPWR _0034_
+ sky130_fd_sc_hd__xnor2_1
X_2639_ _0844_ _0869_ _0968_ _0970_ _0867_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__o41a_1
X_4309_ net194 _1990_ _2254_ _2255_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_2_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2990_ cordic_inst.cordic_inst.x\[9\] _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__and2b_1
XFILLER_9_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4660_ net377 _0390_ _0092_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.i\[4\] sky130_fd_sc_hd__dfrtp_1
X_3611_ _1777_ _1778_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__or2_1
X_4591_ net385 _0323_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3542_ net175 _1599_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__or2_1
X_3473_ net180 _1699_ _1700_ _1701_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a31o_1
X_2424_ net239 _0698_ _0637_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__a21bo_1
X_2355_ net290 _0654_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__or2_1
X_2286_ net107 VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__inv_2
X_4025_ axi_controller.reg_input_data\[0\] _2018_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__or2_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4927_ net372 _0027_ VGND VGND VPWR VPWR cordic_inst.deg_handler_inst.theta_abs\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_4858_ net372 _0067_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.angle\[22\] sky130_fd_sc_hd__dfxtp_1
X_3809_ _1905_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__inv_2
XFILLER_21_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4789_ net404 _0516_ _0211_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.x\[18\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_7_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2973_ _1263_ _1275_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__nand2_1
XFILLER_34_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4712_ net367 _0439_ _0134_ VGND VGND VPWR VPWR cordic_inst.cordic_inst.z\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4643_ net394 _0374_ net333 VGND VGND VPWR VPWR axi_controller.result_out\[20\] sky130_fd_sc_hd__dfrtp_1
X_4574_ net364 _0306_ VGND VGND VPWR VPWR axi_controller.write_addr_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3525_ _1556_ _1609_ _1739_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__a21oi_1
X_3456_ cordic_inst.cordic_inst.angle\[25\] net173 net161 cordic_inst.cordic_inst.z\[25\]
+ _1688_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__a221o_1
X_2407_ _0740_ _0741_ net277 _0664_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__a2bb2o_1
X_3387_ _1554_ _1610_ _1618_ _1622_ _1547_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__o2111ai_2
X_2338_ cordic_inst.cordic_inst.x\[10\] cordic_inst.cordic_inst.x\[11\] cordic_inst.cordic_inst.x\[12\]
+ cordic_inst.cordic_inst.x\[13\] net309 net298 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux4_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2269_ net274 VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__inv_2
X_4008_ net87 _2009_ _2010_ net346 VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o211a_1
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3310_ net266 _1481_ _1548_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__mux2_1
X_4290_ net78 _2243_ _2244_ net347 VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__o211a_1
X_3241_ _1478_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__nand2_1
X_3172_ _1293_ _1440_ _1323_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2956_ cordic_inst.cordic_inst.x\[4\] _1256_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__nor2_1
X_2887_ net262 _1080_ _1174_ _1171_ net238 net242 VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__mux4_2
X_4626_ net398 _0357_ net339 VGND VGND VPWR VPWR axi_controller.result_out\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4557_ net362 _0289_ VGND VGND VPWR VPWR axi_controller.read_addr_reg\[23\] sky130_fd_sc_hd__dfxtp_1
X_4488_ net330 VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__inv_2
X_3508_ _1727_ net179 _1627_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__and3b_1
X_3439_ cordic_inst.cordic_inst.angle\[29\] net174 net162 cordic_inst.cordic_inst.z\[29\]
+ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__a22o_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3790_ _1874_ _1890_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__nor2_1
X_2810_ _1078_ _1112_ net232 VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__mux2_1
XFILLER_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2741_ _0955_ _0957_ _1037_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nand3_1
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4411_ net328 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__inv_2
X_2672_ _0812_ _0999_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__nand2_1
X_4342_ net123 net191 net155 axi_controller.result_out\[1\] VGND VGND VPWR VPWR _0593_
+ sky130_fd_sc_hd__a22o_1
Xfanout319 axi_controller.rst VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__buf_2
Xfanout308 net311 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_4
X_4273_ axi_controller.result_out\[30\] net200 VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__nor2_1
X_3224_ cordic_inst.cordic_inst.y\[9\] cordic_inst.cordic_inst.sin_out\[9\] net210
+ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
.ends

