module cordic_system (aclk,
    aresetn,
    arready,
    arvalid,
    awready,
    awvalid,
    bready,
    bvalid,
    rready,
    rvalid,
    wready,
    wvalid,
    araddr,
    awaddr,
    bresp,
    rdata,
    rresp,
    wdata,
    wstrb);
 input aclk;
 input aresetn;
 output arready;
 input arvalid;
 output awready;
 input awvalid;
 input bready;
 output bvalid;
 input rready;
 output rvalid;
 output wready;
 input wvalid;
 input [31:0] araddr;
 input [31:0] awaddr;
 output [1:0] bresp;
 output [31:0] rdata;
 output [1:0] rresp;
 input [31:0] wdata;
 input [3:0] wstrb;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire \axi_controller.done ;
 wire \axi_controller.mode ;
 wire \axi_controller.read_addr_reg[0] ;
 wire \axi_controller.read_addr_reg[10] ;
 wire \axi_controller.read_addr_reg[11] ;
 wire \axi_controller.read_addr_reg[12] ;
 wire \axi_controller.read_addr_reg[13] ;
 wire \axi_controller.read_addr_reg[14] ;
 wire \axi_controller.read_addr_reg[15] ;
 wire \axi_controller.read_addr_reg[16] ;
 wire \axi_controller.read_addr_reg[17] ;
 wire \axi_controller.read_addr_reg[18] ;
 wire \axi_controller.read_addr_reg[19] ;
 wire \axi_controller.read_addr_reg[1] ;
 wire \axi_controller.read_addr_reg[20] ;
 wire \axi_controller.read_addr_reg[21] ;
 wire \axi_controller.read_addr_reg[22] ;
 wire \axi_controller.read_addr_reg[23] ;
 wire \axi_controller.read_addr_reg[24] ;
 wire \axi_controller.read_addr_reg[25] ;
 wire \axi_controller.read_addr_reg[26] ;
 wire \axi_controller.read_addr_reg[27] ;
 wire \axi_controller.read_addr_reg[28] ;
 wire \axi_controller.read_addr_reg[29] ;
 wire \axi_controller.read_addr_reg[2] ;
 wire \axi_controller.read_addr_reg[30] ;
 wire \axi_controller.read_addr_reg[31] ;
 wire \axi_controller.read_addr_reg[3] ;
 wire \axi_controller.read_addr_reg[4] ;
 wire \axi_controller.read_addr_reg[5] ;
 wire \axi_controller.read_addr_reg[6] ;
 wire \axi_controller.read_addr_reg[7] ;
 wire \axi_controller.read_addr_reg[8] ;
 wire \axi_controller.read_addr_reg[9] ;
 wire \axi_controller.reg_done_flag ;
 wire \axi_controller.reg_input_data[0] ;
 wire \axi_controller.reg_input_data[10] ;
 wire \axi_controller.reg_input_data[11] ;
 wire \axi_controller.reg_input_data[12] ;
 wire \axi_controller.reg_input_data[13] ;
 wire \axi_controller.reg_input_data[14] ;
 wire \axi_controller.reg_input_data[15] ;
 wire \axi_controller.reg_input_data[16] ;
 wire \axi_controller.reg_input_data[17] ;
 wire \axi_controller.reg_input_data[18] ;
 wire \axi_controller.reg_input_data[19] ;
 wire \axi_controller.reg_input_data[1] ;
 wire \axi_controller.reg_input_data[20] ;
 wire \axi_controller.reg_input_data[21] ;
 wire \axi_controller.reg_input_data[22] ;
 wire \axi_controller.reg_input_data[23] ;
 wire \axi_controller.reg_input_data[24] ;
 wire \axi_controller.reg_input_data[25] ;
 wire \axi_controller.reg_input_data[26] ;
 wire \axi_controller.reg_input_data[27] ;
 wire \axi_controller.reg_input_data[28] ;
 wire \axi_controller.reg_input_data[29] ;
 wire \axi_controller.reg_input_data[2] ;
 wire \axi_controller.reg_input_data[30] ;
 wire \axi_controller.reg_input_data[31] ;
 wire \axi_controller.reg_input_data[3] ;
 wire \axi_controller.reg_input_data[4] ;
 wire \axi_controller.reg_input_data[5] ;
 wire \axi_controller.reg_input_data[6] ;
 wire \axi_controller.reg_input_data[7] ;
 wire \axi_controller.reg_input_data[8] ;
 wire \axi_controller.reg_input_data[9] ;
 wire \axi_controller.result_out[0] ;
 wire \axi_controller.result_out[10] ;
 wire \axi_controller.result_out[11] ;
 wire \axi_controller.result_out[12] ;
 wire \axi_controller.result_out[13] ;
 wire \axi_controller.result_out[14] ;
 wire \axi_controller.result_out[15] ;
 wire \axi_controller.result_out[16] ;
 wire \axi_controller.result_out[17] ;
 wire \axi_controller.result_out[18] ;
 wire \axi_controller.result_out[19] ;
 wire \axi_controller.result_out[1] ;
 wire \axi_controller.result_out[20] ;
 wire \axi_controller.result_out[21] ;
 wire \axi_controller.result_out[22] ;
 wire \axi_controller.result_out[23] ;
 wire \axi_controller.result_out[24] ;
 wire \axi_controller.result_out[25] ;
 wire \axi_controller.result_out[26] ;
 wire \axi_controller.result_out[27] ;
 wire \axi_controller.result_out[28] ;
 wire \axi_controller.result_out[29] ;
 wire \axi_controller.result_out[2] ;
 wire \axi_controller.result_out[30] ;
 wire \axi_controller.result_out[31] ;
 wire \axi_controller.result_out[3] ;
 wire \axi_controller.result_out[4] ;
 wire \axi_controller.result_out[5] ;
 wire \axi_controller.result_out[6] ;
 wire \axi_controller.result_out[7] ;
 wire \axi_controller.result_out[8] ;
 wire \axi_controller.result_out[9] ;
 wire \axi_controller.rst ;
 wire \axi_controller.start_pulse_reg ;
 wire \axi_controller.state[0] ;
 wire \axi_controller.state[1] ;
 wire \axi_controller.state[2] ;
 wire \axi_controller.state[3] ;
 wire \axi_controller.write_addr_reg[0] ;
 wire \axi_controller.write_addr_reg[10] ;
 wire \axi_controller.write_addr_reg[11] ;
 wire \axi_controller.write_addr_reg[12] ;
 wire \axi_controller.write_addr_reg[13] ;
 wire \axi_controller.write_addr_reg[14] ;
 wire \axi_controller.write_addr_reg[15] ;
 wire \axi_controller.write_addr_reg[16] ;
 wire \axi_controller.write_addr_reg[17] ;
 wire \axi_controller.write_addr_reg[18] ;
 wire \axi_controller.write_addr_reg[19] ;
 wire \axi_controller.write_addr_reg[1] ;
 wire \axi_controller.write_addr_reg[20] ;
 wire \axi_controller.write_addr_reg[21] ;
 wire \axi_controller.write_addr_reg[22] ;
 wire \axi_controller.write_addr_reg[23] ;
 wire \axi_controller.write_addr_reg[24] ;
 wire \axi_controller.write_addr_reg[25] ;
 wire \axi_controller.write_addr_reg[26] ;
 wire \axi_controller.write_addr_reg[27] ;
 wire \axi_controller.write_addr_reg[28] ;
 wire \axi_controller.write_addr_reg[29] ;
 wire \axi_controller.write_addr_reg[2] ;
 wire \axi_controller.write_addr_reg[30] ;
 wire \axi_controller.write_addr_reg[31] ;
 wire \axi_controller.write_addr_reg[3] ;
 wire \axi_controller.write_addr_reg[4] ;
 wire \axi_controller.write_addr_reg[5] ;
 wire \axi_controller.write_addr_reg[6] ;
 wire \axi_controller.write_addr_reg[7] ;
 wire \axi_controller.write_addr_reg[8] ;
 wire \axi_controller.write_addr_reg[9] ;
 wire net410;
 wire \cordic_inst.cordic_inst.angle[0] ;
 wire \cordic_inst.cordic_inst.angle[10] ;
 wire \cordic_inst.cordic_inst.angle[11] ;
 wire \cordic_inst.cordic_inst.angle[12] ;
 wire \cordic_inst.cordic_inst.angle[13] ;
 wire \cordic_inst.cordic_inst.angle[14] ;
 wire \cordic_inst.cordic_inst.angle[15] ;
 wire \cordic_inst.cordic_inst.angle[16] ;
 wire \cordic_inst.cordic_inst.angle[17] ;
 wire \cordic_inst.cordic_inst.angle[18] ;
 wire \cordic_inst.cordic_inst.angle[19] ;
 wire \cordic_inst.cordic_inst.angle[1] ;
 wire \cordic_inst.cordic_inst.angle[20] ;
 wire \cordic_inst.cordic_inst.angle[21] ;
 wire \cordic_inst.cordic_inst.angle[22] ;
 wire \cordic_inst.cordic_inst.angle[23] ;
 wire \cordic_inst.cordic_inst.angle[24] ;
 wire \cordic_inst.cordic_inst.angle[25] ;
 wire \cordic_inst.cordic_inst.angle[26] ;
 wire \cordic_inst.cordic_inst.angle[27] ;
 wire \cordic_inst.cordic_inst.angle[28] ;
 wire \cordic_inst.cordic_inst.angle[29] ;
 wire \cordic_inst.cordic_inst.angle[2] ;
 wire \cordic_inst.cordic_inst.angle[30] ;
 wire \cordic_inst.cordic_inst.angle[31] ;
 wire \cordic_inst.cordic_inst.angle[3] ;
 wire \cordic_inst.cordic_inst.angle[4] ;
 wire \cordic_inst.cordic_inst.angle[5] ;
 wire \cordic_inst.cordic_inst.angle[6] ;
 wire \cordic_inst.cordic_inst.angle[7] ;
 wire \cordic_inst.cordic_inst.angle[8] ;
 wire \cordic_inst.cordic_inst.angle[9] ;
 wire \cordic_inst.cordic_inst.cos_out[0] ;
 wire \cordic_inst.cordic_inst.cos_out[10] ;
 wire \cordic_inst.cordic_inst.cos_out[11] ;
 wire \cordic_inst.cordic_inst.cos_out[12] ;
 wire \cordic_inst.cordic_inst.cos_out[13] ;
 wire \cordic_inst.cordic_inst.cos_out[14] ;
 wire \cordic_inst.cordic_inst.cos_out[15] ;
 wire \cordic_inst.cordic_inst.cos_out[16] ;
 wire \cordic_inst.cordic_inst.cos_out[17] ;
 wire \cordic_inst.cordic_inst.cos_out[18] ;
 wire \cordic_inst.cordic_inst.cos_out[19] ;
 wire \cordic_inst.cordic_inst.cos_out[1] ;
 wire \cordic_inst.cordic_inst.cos_out[20] ;
 wire \cordic_inst.cordic_inst.cos_out[21] ;
 wire \cordic_inst.cordic_inst.cos_out[22] ;
 wire \cordic_inst.cordic_inst.cos_out[23] ;
 wire \cordic_inst.cordic_inst.cos_out[24] ;
 wire \cordic_inst.cordic_inst.cos_out[25] ;
 wire \cordic_inst.cordic_inst.cos_out[26] ;
 wire \cordic_inst.cordic_inst.cos_out[27] ;
 wire \cordic_inst.cordic_inst.cos_out[28] ;
 wire \cordic_inst.cordic_inst.cos_out[29] ;
 wire \cordic_inst.cordic_inst.cos_out[2] ;
 wire \cordic_inst.cordic_inst.cos_out[30] ;
 wire \cordic_inst.cordic_inst.cos_out[31] ;
 wire \cordic_inst.cordic_inst.cos_out[3] ;
 wire \cordic_inst.cordic_inst.cos_out[4] ;
 wire \cordic_inst.cordic_inst.cos_out[5] ;
 wire \cordic_inst.cordic_inst.cos_out[6] ;
 wire \cordic_inst.cordic_inst.cos_out[7] ;
 wire \cordic_inst.cordic_inst.cos_out[8] ;
 wire \cordic_inst.cordic_inst.cos_out[9] ;
 wire \cordic_inst.cordic_inst.done ;
 wire \cordic_inst.cordic_inst.i[0] ;
 wire \cordic_inst.cordic_inst.i[1] ;
 wire \cordic_inst.cordic_inst.i[2] ;
 wire \cordic_inst.cordic_inst.i[3] ;
 wire \cordic_inst.cordic_inst.i[4] ;
 wire \cordic_inst.cordic_inst.next_state[0] ;
 wire \cordic_inst.cordic_inst.next_state[1] ;
 wire \cordic_inst.cordic_inst.sin_out[0] ;
 wire \cordic_inst.cordic_inst.sin_out[10] ;
 wire \cordic_inst.cordic_inst.sin_out[11] ;
 wire \cordic_inst.cordic_inst.sin_out[12] ;
 wire \cordic_inst.cordic_inst.sin_out[13] ;
 wire \cordic_inst.cordic_inst.sin_out[14] ;
 wire \cordic_inst.cordic_inst.sin_out[15] ;
 wire \cordic_inst.cordic_inst.sin_out[16] ;
 wire \cordic_inst.cordic_inst.sin_out[17] ;
 wire \cordic_inst.cordic_inst.sin_out[18] ;
 wire \cordic_inst.cordic_inst.sin_out[19] ;
 wire \cordic_inst.cordic_inst.sin_out[1] ;
 wire \cordic_inst.cordic_inst.sin_out[20] ;
 wire \cordic_inst.cordic_inst.sin_out[21] ;
 wire \cordic_inst.cordic_inst.sin_out[22] ;
 wire \cordic_inst.cordic_inst.sin_out[23] ;
 wire \cordic_inst.cordic_inst.sin_out[24] ;
 wire \cordic_inst.cordic_inst.sin_out[25] ;
 wire \cordic_inst.cordic_inst.sin_out[26] ;
 wire \cordic_inst.cordic_inst.sin_out[27] ;
 wire \cordic_inst.cordic_inst.sin_out[28] ;
 wire \cordic_inst.cordic_inst.sin_out[29] ;
 wire \cordic_inst.cordic_inst.sin_out[2] ;
 wire \cordic_inst.cordic_inst.sin_out[30] ;
 wire \cordic_inst.cordic_inst.sin_out[31] ;
 wire \cordic_inst.cordic_inst.sin_out[3] ;
 wire \cordic_inst.cordic_inst.sin_out[4] ;
 wire \cordic_inst.cordic_inst.sin_out[5] ;
 wire \cordic_inst.cordic_inst.sin_out[6] ;
 wire \cordic_inst.cordic_inst.sin_out[7] ;
 wire \cordic_inst.cordic_inst.sin_out[8] ;
 wire \cordic_inst.cordic_inst.sin_out[9] ;
 wire \cordic_inst.cordic_inst.start ;
 wire \cordic_inst.cordic_inst.state[0] ;
 wire \cordic_inst.cordic_inst.state[1] ;
 wire \cordic_inst.cordic_inst.x[0] ;
 wire \cordic_inst.cordic_inst.x[10] ;
 wire \cordic_inst.cordic_inst.x[11] ;
 wire \cordic_inst.cordic_inst.x[12] ;
 wire \cordic_inst.cordic_inst.x[13] ;
 wire \cordic_inst.cordic_inst.x[14] ;
 wire \cordic_inst.cordic_inst.x[15] ;
 wire \cordic_inst.cordic_inst.x[16] ;
 wire \cordic_inst.cordic_inst.x[17] ;
 wire \cordic_inst.cordic_inst.x[18] ;
 wire \cordic_inst.cordic_inst.x[19] ;
 wire \cordic_inst.cordic_inst.x[1] ;
 wire \cordic_inst.cordic_inst.x[20] ;
 wire \cordic_inst.cordic_inst.x[21] ;
 wire \cordic_inst.cordic_inst.x[22] ;
 wire \cordic_inst.cordic_inst.x[23] ;
 wire \cordic_inst.cordic_inst.x[24] ;
 wire \cordic_inst.cordic_inst.x[25] ;
 wire \cordic_inst.cordic_inst.x[26] ;
 wire \cordic_inst.cordic_inst.x[27] ;
 wire \cordic_inst.cordic_inst.x[28] ;
 wire \cordic_inst.cordic_inst.x[29] ;
 wire \cordic_inst.cordic_inst.x[2] ;
 wire \cordic_inst.cordic_inst.x[30] ;
 wire \cordic_inst.cordic_inst.x[31] ;
 wire \cordic_inst.cordic_inst.x[3] ;
 wire \cordic_inst.cordic_inst.x[4] ;
 wire \cordic_inst.cordic_inst.x[5] ;
 wire \cordic_inst.cordic_inst.x[6] ;
 wire \cordic_inst.cordic_inst.x[7] ;
 wire \cordic_inst.cordic_inst.x[8] ;
 wire \cordic_inst.cordic_inst.x[9] ;
 wire \cordic_inst.cordic_inst.y[0] ;
 wire \cordic_inst.cordic_inst.y[10] ;
 wire \cordic_inst.cordic_inst.y[11] ;
 wire \cordic_inst.cordic_inst.y[12] ;
 wire \cordic_inst.cordic_inst.y[13] ;
 wire \cordic_inst.cordic_inst.y[14] ;
 wire \cordic_inst.cordic_inst.y[15] ;
 wire \cordic_inst.cordic_inst.y[16] ;
 wire \cordic_inst.cordic_inst.y[17] ;
 wire \cordic_inst.cordic_inst.y[18] ;
 wire \cordic_inst.cordic_inst.y[19] ;
 wire \cordic_inst.cordic_inst.y[1] ;
 wire \cordic_inst.cordic_inst.y[20] ;
 wire \cordic_inst.cordic_inst.y[21] ;
 wire \cordic_inst.cordic_inst.y[22] ;
 wire \cordic_inst.cordic_inst.y[23] ;
 wire \cordic_inst.cordic_inst.y[24] ;
 wire \cordic_inst.cordic_inst.y[25] ;
 wire \cordic_inst.cordic_inst.y[26] ;
 wire \cordic_inst.cordic_inst.y[27] ;
 wire \cordic_inst.cordic_inst.y[28] ;
 wire \cordic_inst.cordic_inst.y[29] ;
 wire \cordic_inst.cordic_inst.y[2] ;
 wire \cordic_inst.cordic_inst.y[30] ;
 wire \cordic_inst.cordic_inst.y[31] ;
 wire \cordic_inst.cordic_inst.y[3] ;
 wire \cordic_inst.cordic_inst.y[4] ;
 wire \cordic_inst.cordic_inst.y[5] ;
 wire \cordic_inst.cordic_inst.y[6] ;
 wire \cordic_inst.cordic_inst.y[7] ;
 wire \cordic_inst.cordic_inst.y[8] ;
 wire \cordic_inst.cordic_inst.y[9] ;
 wire \cordic_inst.cordic_inst.z[0] ;
 wire \cordic_inst.cordic_inst.z[10] ;
 wire \cordic_inst.cordic_inst.z[11] ;
 wire \cordic_inst.cordic_inst.z[12] ;
 wire \cordic_inst.cordic_inst.z[13] ;
 wire \cordic_inst.cordic_inst.z[14] ;
 wire \cordic_inst.cordic_inst.z[15] ;
 wire \cordic_inst.cordic_inst.z[16] ;
 wire \cordic_inst.cordic_inst.z[17] ;
 wire \cordic_inst.cordic_inst.z[18] ;
 wire \cordic_inst.cordic_inst.z[19] ;
 wire \cordic_inst.cordic_inst.z[1] ;
 wire \cordic_inst.cordic_inst.z[20] ;
 wire \cordic_inst.cordic_inst.z[21] ;
 wire \cordic_inst.cordic_inst.z[22] ;
 wire \cordic_inst.cordic_inst.z[23] ;
 wire \cordic_inst.cordic_inst.z[24] ;
 wire \cordic_inst.cordic_inst.z[25] ;
 wire \cordic_inst.cordic_inst.z[26] ;
 wire \cordic_inst.cordic_inst.z[27] ;
 wire \cordic_inst.cordic_inst.z[28] ;
 wire \cordic_inst.cordic_inst.z[29] ;
 wire \cordic_inst.cordic_inst.z[2] ;
 wire \cordic_inst.cordic_inst.z[30] ;
 wire \cordic_inst.cordic_inst.z[31] ;
 wire \cordic_inst.cordic_inst.z[3] ;
 wire \cordic_inst.cordic_inst.z[4] ;
 wire \cordic_inst.cordic_inst.z[5] ;
 wire \cordic_inst.cordic_inst.z[6] ;
 wire \cordic_inst.cordic_inst.z[7] ;
 wire \cordic_inst.cordic_inst.z[8] ;
 wire \cordic_inst.cordic_inst.z[9] ;
 wire \cordic_inst.deg_handler_inst.isNegative ;
 wire \cordic_inst.deg_handler_inst.kuadran[0] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[0] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[10] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[11] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[12] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[13] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[14] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[15] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[16] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[17] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[18] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[19] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[1] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[20] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[21] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[22] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[23] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[24] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[25] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[26] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[27] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[28] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[29] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[2] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[30] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[31] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[3] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[4] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[5] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[6] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[7] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[8] ;
 wire \cordic_inst.deg_handler_inst.theta_abs[9] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[0] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[10] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[11] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[12] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[13] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[14] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[15] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[16] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[17] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[18] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[19] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[1] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[20] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[21] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[22] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[23] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[24] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[25] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[26] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[27] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[28] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[29] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[2] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[30] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[31] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[3] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[4] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[5] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[6] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[7] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[8] ;
 wire \cordic_inst.deg_handler_inst.theta_norm[9] ;
 wire \cordic_inst.done_d ;
 wire \cordic_inst.sign_handler_inst.done_d ;
 wire \cordic_inst.sign_handler_inst.done_pulse ;
 wire \cordic_inst.state[0] ;
 wire \cordic_inst.state[1] ;
 wire \cordic_inst.state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;

 sky130_fd_sc_hd__inv_2 _2258_ (.A(\cordic_inst.cordic_inst.y[28] ),
    .Y(_0595_));
 sky130_fd_sc_hd__inv_2 _2259_ (.A(\cordic_inst.cordic_inst.y[18] ),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _2260_ (.A(\cordic_inst.cordic_inst.y[10] ),
    .Y(_0597_));
 sky130_fd_sc_hd__inv_2 _2261_ (.A(\cordic_inst.cordic_inst.y[8] ),
    .Y(_0598_));
 sky130_fd_sc_hd__inv_2 _2262_ (.A(\cordic_inst.cordic_inst.y[5] ),
    .Y(_0599_));
 sky130_fd_sc_hd__inv_2 _2263_ (.A(\cordic_inst.cordic_inst.y[0] ),
    .Y(_0600_));
 sky130_fd_sc_hd__inv_2 _2264_ (.A(net264),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_2 _2265_ (.A(\cordic_inst.cordic_inst.x[5] ),
    .Y(_0602_));
 sky130_fd_sc_hd__inv_2 _2266_ (.A(\cordic_inst.cordic_inst.x[0] ),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _2267_ (.A(net270),
    .Y(_0604_));
 sky130_fd_sc_hd__inv_2 _2268_ (.A(\cordic_inst.cordic_inst.cos_out[26] ),
    .Y(_0605_));
 sky130_fd_sc_hd__inv_2 _2269_ (.A(net274),
    .Y(_0606_));
 sky130_fd_sc_hd__inv_2 _2270_ (.A(net282),
    .Y(_0607_));
 sky130_fd_sc_hd__inv_2 _2271_ (.A(net289),
    .Y(_0608_));
 sky130_fd_sc_hd__inv_2 _2272_ (.A(net296),
    .Y(_0609_));
 sky130_fd_sc_hd__inv_2 _2273_ (.A(\axi_controller.state[0] ),
    .Y(_0610_));
 sky130_fd_sc_hd__inv_2 _2274_ (.A(net110),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _2275_ (.A(net315),
    .Y(_0612_));
 sky130_fd_sc_hd__inv_2 _2276_ (.A(net318),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _2277_ (.A(\cordic_inst.deg_handler_inst.kuadran[0] ),
    .Y(_0613_));
 sky130_fd_sc_hd__inv_2 _2278_ (.A(\cordic_inst.cordic_inst.state[1] ),
    .Y(_0614_));
 sky130_fd_sc_hd__inv_2 _2279_ (.A(\cordic_inst.deg_handler_inst.theta_abs[18] ),
    .Y(_0615_));
 sky130_fd_sc_hd__inv_2 _2280_ (.A(\cordic_inst.deg_handler_inst.theta_abs[20] ),
    .Y(_0616_));
 sky130_fd_sc_hd__inv_2 _2281_ (.A(\cordic_inst.deg_handler_inst.theta_abs[22] ),
    .Y(_0617_));
 sky130_fd_sc_hd__inv_2 _2282_ (.A(\cordic_inst.state[0] ),
    .Y(_0618_));
 sky130_fd_sc_hd__inv_2 _2283_ (.A(\axi_controller.state[1] ),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_2 _2284_ (.A(\cordic_inst.state[1] ),
    .Y(_0620_));
 sky130_fd_sc_hd__inv_2 _2285_ (.A(net349),
    .Y(_0621_));
 sky130_fd_sc_hd__inv_2 _2286_ (.A(net107),
    .Y(_0622_));
 sky130_fd_sc_hd__inv_2 _2287_ (.A(\axi_controller.write_addr_reg[4] ),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _2288_ (.A(\axi_controller.state[3] ),
    .Y(_0624_));
 sky130_fd_sc_hd__inv_2 _2289_ (.A(\axi_controller.read_addr_reg[31] ),
    .Y(_0625_));
 sky130_fd_sc_hd__nor2_1 _2290_ (.A(_0614_),
    .B(\cordic_inst.cordic_inst.state[0] ),
    .Y(_0626_));
 sky130_fd_sc_hd__or2_1 _2291_ (.A(_0614_),
    .B(\cordic_inst.cordic_inst.state[0] ),
    .X(_0627_));
 sky130_fd_sc_hd__and2_1 _2292_ (.A(_0614_),
    .B(\cordic_inst.cordic_inst.state[0] ),
    .X(_0628_));
 sky130_fd_sc_hd__nor2_2 _2293_ (.A(net181),
    .B(net174),
    .Y(_0629_));
 sky130_fd_sc_hd__inv_2 _2294_ (.A(net162),
    .Y(\cordic_inst.cordic_inst.next_state[1] ));
 sky130_fd_sc_hd__nor2_1 _2295_ (.A(_0601_),
    .B(net244),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_1 _2296_ (.A(net264),
    .B(net278),
    .Y(_0631_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(\cordic_inst.cordic_inst.x[30] ),
    .A1(net265),
    .S(net304),
    .X(_0632_));
 sky130_fd_sc_hd__and2_1 _2298_ (.A(net264),
    .B(net295),
    .X(_0633_));
 sky130_fd_sc_hd__a21o_1 _2299_ (.A1(_0609_),
    .A2(_0632_),
    .B1(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__and2_1 _2300_ (.A(net264),
    .B(net291),
    .X(_0635_));
 sky130_fd_sc_hd__a21oi_1 _2301_ (.A1(net233),
    .A2(_0634_),
    .B1(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_2 _2302_ (.A(net264),
    .B(net286),
    .Y(_0637_));
 sky130_fd_sc_hd__o21ai_1 _2303_ (.A1(net286),
    .A2(_0636_),
    .B1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__a21o_1 _2304_ (.A1(_0606_),
    .A2(_0638_),
    .B1(net170),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _2305_ (.A0(\cordic_inst.cordic_inst.x[28] ),
    .A1(\cordic_inst.cordic_inst.x[29] ),
    .S(net304),
    .X(_0640_));
 sky130_fd_sc_hd__mux4_1 _2306_ (.A0(\cordic_inst.cordic_inst.x[28] ),
    .A1(\cordic_inst.cordic_inst.x[29] ),
    .A2(\cordic_inst.cordic_inst.x[30] ),
    .A3(net265),
    .S0(net305),
    .S1(net296),
    .X(_0641_));
 sky130_fd_sc_hd__a21o_1 _2307_ (.A1(net234),
    .A2(_0641_),
    .B1(_0635_),
    .X(_0642_));
 sky130_fd_sc_hd__a21bo_1 _2308_ (.A1(net239),
    .A2(_0642_),
    .B1_N(_0637_),
    .X(_0643_));
 sky130_fd_sc_hd__a21o_1 _2309_ (.A1(net242),
    .A2(_0643_),
    .B1(net170),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _2310_ (.A0(\cordic_inst.cordic_inst.x[25] ),
    .A1(\cordic_inst.cordic_inst.x[26] ),
    .S(net307),
    .X(_0645_));
 sky130_fd_sc_hd__mux4_1 _2311_ (.A0(\cordic_inst.cordic_inst.x[23] ),
    .A1(\cordic_inst.cordic_inst.x[24] ),
    .A2(\cordic_inst.cordic_inst.x[25] ),
    .A3(\cordic_inst.cordic_inst.x[26] ),
    .S0(net307),
    .S1(net301),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _2312_ (.A0(\cordic_inst.cordic_inst.x[27] ),
    .A1(\cordic_inst.cordic_inst.x[28] ),
    .S(net304),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _2313_ (.A0(\cordic_inst.cordic_inst.x[29] ),
    .A1(\cordic_inst.cordic_inst.x[30] ),
    .S(net305),
    .X(_0648_));
 sky130_fd_sc_hd__mux4_1 _2314_ (.A0(\cordic_inst.cordic_inst.x[27] ),
    .A1(\cordic_inst.cordic_inst.x[28] ),
    .A2(\cordic_inst.cordic_inst.x[29] ),
    .A3(\cordic_inst.cordic_inst.x[30] ),
    .S0(net305),
    .S1(net296),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _2315_ (.A0(_0646_),
    .A1(_0649_),
    .S(net291),
    .X(_0650_));
 sky130_fd_sc_hd__a21boi_1 _2316_ (.A1(net239),
    .A2(_0650_),
    .B1_N(_0637_),
    .Y(_0651_));
 sky130_fd_sc_hd__nor2_1 _2317_ (.A(net278),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__mux4_1 _2318_ (.A0(\cordic_inst.cordic_inst.x[18] ),
    .A1(\cordic_inst.cordic_inst.x[19] ),
    .A2(\cordic_inst.cordic_inst.x[20] ),
    .A3(\cordic_inst.cordic_inst.x[21] ),
    .S0(net311),
    .S1(net300),
    .X(_0653_));
 sky130_fd_sc_hd__mux4_1 _2319_ (.A0(\cordic_inst.cordic_inst.x[22] ),
    .A1(\cordic_inst.cordic_inst.x[23] ),
    .A2(\cordic_inst.cordic_inst.x[24] ),
    .A3(\cordic_inst.cordic_inst.x[25] ),
    .S0(net307),
    .S1(net301),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _2320_ (.A0(_0653_),
    .A1(_0654_),
    .S(net292),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _2321_ (.A0(\cordic_inst.cordic_inst.x[26] ),
    .A1(\cordic_inst.cordic_inst.x[27] ),
    .S(net304),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _2322_ (.A0(_0640_),
    .A1(_0656_),
    .S(_0609_),
    .X(_0657_));
 sky130_fd_sc_hd__mux4_2 _2323_ (.A0(net265),
    .A1(_0632_),
    .A2(_0640_),
    .A3(_0656_),
    .S0(_0609_),
    .S1(net234),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(_0655_),
    .A1(_0658_),
    .S(net285),
    .X(_0659_));
 sky130_fd_sc_hd__mux4_1 _2325_ (.A0(\cordic_inst.cordic_inst.x[19] ),
    .A1(\cordic_inst.cordic_inst.x[20] ),
    .A2(\cordic_inst.cordic_inst.x[21] ),
    .A3(\cordic_inst.cordic_inst.x[22] ),
    .S0(net311),
    .S1(net300),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(_0646_),
    .A1(_0660_),
    .S(net236),
    .X(_0661_));
 sky130_fd_sc_hd__a21oi_1 _2327_ (.A1(net234),
    .A2(_0649_),
    .B1(_0635_),
    .Y(_0662_));
 sky130_fd_sc_hd__a211o_1 _2328_ (.A1(net234),
    .A2(_0649_),
    .B1(_0635_),
    .C1(net238),
    .X(_0663_));
 sky130_fd_sc_hd__o21ai_1 _2329_ (.A1(net285),
    .A2(_0661_),
    .B1(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__nor2_1 _2330_ (.A(net278),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nor2_1 _2331_ (.A(net170),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__a21o_1 _2332_ (.A1(net245),
    .A2(_0659_),
    .B1(net170),
    .X(_0667_));
 sky130_fd_sc_hd__mux4_1 _2333_ (.A0(\cordic_inst.cordic_inst.x[15] ),
    .A1(\cordic_inst.cordic_inst.x[16] ),
    .A2(\cordic_inst.cordic_inst.x[17] ),
    .A3(\cordic_inst.cordic_inst.x[18] ),
    .S0(net311),
    .S1(net299),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(_0660_),
    .A1(_0668_),
    .S(net236),
    .X(_0669_));
 sky130_fd_sc_hd__nor2_1 _2335_ (.A(net285),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _2336_ (.A(net240),
    .B(_0650_),
    .Y(_0671_));
 sky130_fd_sc_hd__o31a_1 _2337_ (.A1(net278),
    .A2(_0670_),
    .A3(_0671_),
    .B1(_0631_),
    .X(_0672_));
 sky130_fd_sc_hd__mux4_1 _2338_ (.A0(\cordic_inst.cordic_inst.x[10] ),
    .A1(\cordic_inst.cordic_inst.x[11] ),
    .A2(\cordic_inst.cordic_inst.x[12] ),
    .A3(\cordic_inst.cordic_inst.x[13] ),
    .S0(net309),
    .S1(net298),
    .X(_0673_));
 sky130_fd_sc_hd__mux4_1 _2339_ (.A0(\cordic_inst.cordic_inst.x[14] ),
    .A1(\cordic_inst.cordic_inst.x[15] ),
    .A2(\cordic_inst.cordic_inst.x[16] ),
    .A3(\cordic_inst.cordic_inst.x[17] ),
    .S0(net310),
    .S1(net299),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _2340_ (.A0(_0673_),
    .A1(_0674_),
    .S(net292),
    .X(_0675_));
 sky130_fd_sc_hd__a21bo_1 _2341_ (.A1(net239),
    .A2(_0658_),
    .B1_N(_0637_),
    .X(_0676_));
 sky130_fd_sc_hd__mux4_1 _2342_ (.A0(net265),
    .A1(_0655_),
    .A2(_0658_),
    .A3(_0675_),
    .S0(net244),
    .S1(_0607_),
    .X(_0677_));
 sky130_fd_sc_hd__nor2_1 _2343_ (.A(net286),
    .B(net291),
    .Y(_0678_));
 sky130_fd_sc_hd__mux4_1 _2344_ (.A0(\cordic_inst.cordic_inst.x[7] ),
    .A1(\cordic_inst.cordic_inst.x[8] ),
    .A2(\cordic_inst.cordic_inst.x[9] ),
    .A3(\cordic_inst.cordic_inst.x[10] ),
    .S0(net309),
    .S1(net298),
    .X(_0679_));
 sky130_fd_sc_hd__and2b_1 _2345_ (.A_N(net286),
    .B(net291),
    .X(_0680_));
 sky130_fd_sc_hd__mux4_1 _2346_ (.A0(\cordic_inst.cordic_inst.x[11] ),
    .A1(\cordic_inst.cordic_inst.x[12] ),
    .A2(\cordic_inst.cordic_inst.x[13] ),
    .A3(\cordic_inst.cordic_inst.x[14] ),
    .S0(net309),
    .S1(net298),
    .X(_0681_));
 sky130_fd_sc_hd__a221o_1 _2347_ (.A1(net221),
    .A2(_0679_),
    .B1(net219),
    .B2(_0681_),
    .C1(net277),
    .X(_0682_));
 sky130_fd_sc_hd__a21oi_1 _2348_ (.A1(net284),
    .A2(_0669_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a21o_1 _2349_ (.A1(net277),
    .A2(_0651_),
    .B1(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _2350_ (.A0(_0653_),
    .A1(_0674_),
    .S(net235),
    .X(_0685_));
 sky130_fd_sc_hd__inv_2 _2351_ (.A(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__mux4_1 _2352_ (.A0(\cordic_inst.cordic_inst.x[6] ),
    .A1(\cordic_inst.cordic_inst.x[7] ),
    .A2(\cordic_inst.cordic_inst.x[8] ),
    .A3(\cordic_inst.cordic_inst.x[9] ),
    .S0(net309),
    .S1(net297),
    .X(_0687_));
 sky130_fd_sc_hd__a221o_1 _2353_ (.A1(_0673_),
    .A2(net219),
    .B1(_0687_),
    .B2(net221),
    .C1(net277),
    .X(_0688_));
 sky130_fd_sc_hd__a21o_1 _2354_ (.A1(net284),
    .A2(_0685_),
    .B1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__or2_1 _2355_ (.A(net290),
    .B(_0654_),
    .X(_0690_));
 sky130_fd_sc_hd__o21ai_1 _2356_ (.A1(net235),
    .A2(_0657_),
    .B1(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__mux4_2 _2357_ (.A0(net264),
    .A1(_0634_),
    .A2(_0657_),
    .A3(_0654_),
    .S0(net234),
    .S1(net240),
    .X(_0692_));
 sky130_fd_sc_hd__o21ai_2 _2358_ (.A1(net247),
    .A2(_0692_),
    .B1(_0689_),
    .Y(_0693_));
 sky130_fd_sc_hd__mux4_1 _2359_ (.A0(\cordic_inst.cordic_inst.x[16] ),
    .A1(\cordic_inst.cordic_inst.x[17] ),
    .A2(\cordic_inst.cordic_inst.x[18] ),
    .A3(\cordic_inst.cordic_inst.x[19] ),
    .S0(net310),
    .S1(net299),
    .X(_0694_));
 sky130_fd_sc_hd__mux4_1 _2360_ (.A0(\cordic_inst.cordic_inst.x[20] ),
    .A1(\cordic_inst.cordic_inst.x[21] ),
    .A2(\cordic_inst.cordic_inst.x[22] ),
    .A3(\cordic_inst.cordic_inst.x[23] ),
    .S0(net312),
    .S1(net301),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _2361_ (.A0(_0694_),
    .A1(_0695_),
    .S(net292),
    .X(_0696_));
 sky130_fd_sc_hd__mux4_1 _2362_ (.A0(\cordic_inst.cordic_inst.x[24] ),
    .A1(\cordic_inst.cordic_inst.x[25] ),
    .A2(\cordic_inst.cordic_inst.x[26] ),
    .A3(\cordic_inst.cordic_inst.x[27] ),
    .S0(net305),
    .S1(net295),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _2363_ (.A0(_0641_),
    .A1(_0697_),
    .S(net234),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _2364_ (.A0(_0696_),
    .A1(_0698_),
    .S(net285),
    .X(_0699_));
 sky130_fd_sc_hd__mux4_1 _2365_ (.A0(\cordic_inst.cordic_inst.x[8] ),
    .A1(\cordic_inst.cordic_inst.x[9] ),
    .A2(\cordic_inst.cordic_inst.x[10] ),
    .A3(\cordic_inst.cordic_inst.x[11] ),
    .S0(net309),
    .S1(net298),
    .X(_0700_));
 sky130_fd_sc_hd__mux4_1 _2366_ (.A0(\cordic_inst.cordic_inst.x[12] ),
    .A1(\cordic_inst.cordic_inst.x[13] ),
    .A2(\cordic_inst.cordic_inst.x[14] ),
    .A3(\cordic_inst.cordic_inst.x[15] ),
    .S0(net309),
    .S1(net297),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(_0700_),
    .A1(_0701_),
    .S(net292),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(\cordic_inst.cordic_inst.x[4] ),
    .A1(\cordic_inst.cordic_inst.x[5] ),
    .S(net312),
    .X(_0703_));
 sky130_fd_sc_hd__mux4_1 _2369_ (.A0(\cordic_inst.cordic_inst.x[4] ),
    .A1(\cordic_inst.cordic_inst.x[5] ),
    .A2(\cordic_inst.cordic_inst.x[6] ),
    .A3(\cordic_inst.cordic_inst.x[7] ),
    .S0(net311),
    .S1(net300),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_1 _2370_ (.A(net288),
    .B(net294),
    .Y(_0705_));
 sky130_fd_sc_hd__nand2_1 _2371_ (.A(net241),
    .B(net302),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2b_2 _2372_ (.A_N(net294),
    .B(net303),
    .Y(_0707_));
 sky130_fd_sc_hd__nor4b_1 _2373_ (.A(net282),
    .B(net293),
    .C(net295),
    .D_N(net305),
    .Y(_0708_));
 sky130_fd_sc_hd__nor3b_1 _2374_ (.A(net283),
    .B(net290),
    .C_N(net301),
    .Y(_0709_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(\cordic_inst.cordic_inst.x[2] ),
    .A1(\cordic_inst.cordic_inst.x[3] ),
    .S(net312),
    .X(_0710_));
 sky130_fd_sc_hd__nor2_2 _2376_ (.A(net295),
    .B(net305),
    .Y(_0711_));
 sky130_fd_sc_hd__or2_1 _2377_ (.A(net294),
    .B(net302),
    .X(_0712_));
 sky130_fd_sc_hd__and2_2 _2378_ (.A(net232),
    .B(net222),
    .X(_0713_));
 sky130_fd_sc_hd__nand2_1 _2379_ (.A(net222),
    .B(_0711_),
    .Y(_0714_));
 sky130_fd_sc_hd__a221o_1 _2380_ (.A1(\cordic_inst.cordic_inst.x[1] ),
    .A2(net217),
    .B1(net216),
    .B2(_0710_),
    .C1(net276),
    .X(_0715_));
 sky130_fd_sc_hd__a32o_1 _2381_ (.A1(\cordic_inst.cordic_inst.x[0] ),
    .A2(net222),
    .A3(_0711_),
    .B1(_0704_),
    .B2(net219),
    .X(_0716_));
 sky130_fd_sc_hd__a211o_1 _2382_ (.A1(net284),
    .A2(_0702_),
    .B1(_0715_),
    .C1(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__o21a_2 _2383_ (.A1(net247),
    .A2(_0699_),
    .B1(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__mux4_1 _2384_ (.A0(\cordic_inst.cordic_inst.x[17] ),
    .A1(\cordic_inst.cordic_inst.x[18] ),
    .A2(\cordic_inst.cordic_inst.x[19] ),
    .A3(\cordic_inst.cordic_inst.x[20] ),
    .S0(net310),
    .S1(net299),
    .X(_0719_));
 sky130_fd_sc_hd__mux4_1 _2385_ (.A0(\cordic_inst.cordic_inst.x[21] ),
    .A1(\cordic_inst.cordic_inst.x[22] ),
    .A2(\cordic_inst.cordic_inst.x[23] ),
    .A3(\cordic_inst.cordic_inst.x[24] ),
    .S0(net312),
    .S1(net301),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(_0719_),
    .A1(_0720_),
    .S(net290),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(_0645_),
    .A1(_0647_),
    .S(net301),
    .X(_0722_));
 sky130_fd_sc_hd__a21o_1 _2388_ (.A1(net232),
    .A2(_0648_),
    .B1(_0633_),
    .X(_0723_));
 sky130_fd_sc_hd__mux4_2 _2389_ (.A0(net264),
    .A1(_0647_),
    .A2(_0648_),
    .A3(_0645_),
    .S0(net233),
    .S1(net232),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _2390_ (.A0(_0721_),
    .A1(_0724_),
    .S(net285),
    .X(_0725_));
 sky130_fd_sc_hd__mux4_1 _2391_ (.A0(\cordic_inst.cordic_inst.x[9] ),
    .A1(\cordic_inst.cordic_inst.x[10] ),
    .A2(\cordic_inst.cordic_inst.x[11] ),
    .A3(\cordic_inst.cordic_inst.x[12] ),
    .S0(net309),
    .S1(net298),
    .X(_0726_));
 sky130_fd_sc_hd__mux4_2 _2392_ (.A0(\cordic_inst.cordic_inst.x[13] ),
    .A1(\cordic_inst.cordic_inst.x[14] ),
    .A2(\cordic_inst.cordic_inst.x[15] ),
    .A3(\cordic_inst.cordic_inst.x[16] ),
    .S0(net310),
    .S1(net300),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(_0726_),
    .A1(_0727_),
    .S(net290),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _2394_ (.A0(\cordic_inst.cordic_inst.x[5] ),
    .A1(\cordic_inst.cordic_inst.x[6] ),
    .S(net307),
    .X(_0729_));
 sky130_fd_sc_hd__mux4_1 _2395_ (.A0(\cordic_inst.cordic_inst.x[5] ),
    .A1(\cordic_inst.cordic_inst.x[6] ),
    .A2(\cordic_inst.cordic_inst.x[7] ),
    .A3(\cordic_inst.cordic_inst.x[8] ),
    .S0(net308),
    .S1(net297),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(\cordic_inst.cordic_inst.x[3] ),
    .A1(\cordic_inst.cordic_inst.x[4] ),
    .S(net307),
    .X(_0731_));
 sky130_fd_sc_hd__a221o_1 _2397_ (.A1(\cordic_inst.cordic_inst.x[2] ),
    .A2(net217),
    .B1(_0709_),
    .B2(_0731_),
    .C1(net275),
    .X(_0732_));
 sky130_fd_sc_hd__a32o_1 _2398_ (.A1(\cordic_inst.cordic_inst.x[1] ),
    .A2(net222),
    .A3(_0711_),
    .B1(_0730_),
    .B2(net219),
    .X(_0733_));
 sky130_fd_sc_hd__a211o_1 _2399_ (.A1(net284),
    .A2(_0728_),
    .B1(_0732_),
    .C1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__o21a_1 _2400_ (.A1(net243),
    .A2(_0725_),
    .B1(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__a221o_1 _2401_ (.A1(_0703_),
    .A2(net216),
    .B1(_0710_),
    .B2(_0713_),
    .C1(net275),
    .X(_0736_));
 sky130_fd_sc_hd__a22o_1 _2402_ (.A1(net284),
    .A2(_0675_),
    .B1(net218),
    .B2(_0687_),
    .X(_0737_));
 sky130_fd_sc_hd__o22a_1 _2403_ (.A1(net243),
    .A2(_0659_),
    .B1(_0736_),
    .B2(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(_0668_),
    .A1(_0681_),
    .S(net236),
    .X(_0739_));
 sky130_fd_sc_hd__a221o_1 _2405_ (.A1(net216),
    .A2(_0729_),
    .B1(_0731_),
    .B2(_0713_),
    .C1(net275),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _2406_ (.A1(_0679_),
    .A2(net218),
    .B1(_0739_),
    .B2(net284),
    .X(_0741_));
 sky130_fd_sc_hd__a2bb2o_1 _2407_ (.A1_N(_0740_),
    .A2_N(_0741_),
    .B1(net277),
    .B2(_0664_),
    .X(_0742_));
 sky130_fd_sc_hd__nor4b_2 _2408_ (.A(_0718_),
    .B(_0735_),
    .C(_0738_),
    .D_N(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__mux2_1 _2409_ (.A0(_0694_),
    .A1(_0701_),
    .S(net235),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _2410_ (.A1(net218),
    .A2(_0700_),
    .B1(_0704_),
    .B2(net221),
    .X(_0745_));
 sky130_fd_sc_hd__a21oi_1 _2411_ (.A1(net283),
    .A2(_0744_),
    .B1(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__mux2_1 _2412_ (.A0(_0695_),
    .A1(_0697_),
    .S(net290),
    .X(_0747_));
 sky130_fd_sc_hd__a211o_1 _2413_ (.A1(net234),
    .A2(_0641_),
    .B1(_0635_),
    .C1(net238),
    .X(_0748_));
 sky130_fd_sc_hd__o21ai_2 _2414_ (.A1(net285),
    .A2(_0747_),
    .B1(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(_0746_),
    .A1(_0749_),
    .S(net277),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(_0719_),
    .A1(_0727_),
    .S(net235),
    .X(_0751_));
 sky130_fd_sc_hd__a221o_1 _2417_ (.A1(net218),
    .A2(_0726_),
    .B1(_0730_),
    .B2(net221),
    .C1(net277),
    .X(_0752_));
 sky130_fd_sc_hd__a21o_1 _2418_ (.A1(net285),
    .A2(_0751_),
    .B1(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__a21oi_1 _2419_ (.A1(net233),
    .A2(_0723_),
    .B1(_0635_),
    .Y(_0754_));
 sky130_fd_sc_hd__mux4_2 _2420_ (.A0(net265),
    .A1(_0722_),
    .A2(_0723_),
    .A3(_0720_),
    .S0(net240),
    .S1(net235),
    .X(_0755_));
 sky130_fd_sc_hd__o21ai_2 _2421_ (.A1(net244),
    .A2(_0755_),
    .B1(_0753_),
    .Y(_0756_));
 sky130_fd_sc_hd__and2_1 _2422_ (.A(_0750_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__and4_1 _2423_ (.A(_0684_),
    .B(_0693_),
    .C(_0750_),
    .D(_0756_),
    .X(_0758_));
 sky130_fd_sc_hd__a21bo_1 _2424_ (.A1(net239),
    .A2(_0698_),
    .B1_N(_0637_),
    .X(_0759_));
 sky130_fd_sc_hd__mux4_2 _2425_ (.A0(net264),
    .A1(_0696_),
    .A2(_0698_),
    .A3(_0702_),
    .S0(net244),
    .S1(net240),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_1 _2426_ (.A(net238),
    .B(_0724_),
    .Y(_0761_));
 sky130_fd_sc_hd__mux4_1 _2427_ (.A0(net264),
    .A1(_0721_),
    .A2(_0724_),
    .A3(_0728_),
    .S0(net244),
    .S1(_0607_),
    .X(_0762_));
 sky130_fd_sc_hd__or2_1 _2428_ (.A(_0760_),
    .B(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__inv_2 _2429_ (.A(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__nor2_1 _2430_ (.A(_0677_),
    .B(_0763_),
    .Y(_0765_));
 sky130_fd_sc_hd__o21a_1 _2431_ (.A1(net286),
    .A2(_0662_),
    .B1(_0637_),
    .X(_0766_));
 sky130_fd_sc_hd__nand2_1 _2432_ (.A(net287),
    .B(_0661_),
    .Y(_0767_));
 sky130_fd_sc_hd__a21oi_1 _2433_ (.A1(net240),
    .A2(_0739_),
    .B1(net277),
    .Y(_0768_));
 sky130_fd_sc_hd__a22o_1 _2434_ (.A1(net278),
    .A2(_0766_),
    .B1(_0767_),
    .B2(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__and4_1 _2435_ (.A(net154),
    .B(_0758_),
    .C(_0765_),
    .D(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__nand4_2 _2436_ (.A(net154),
    .B(_0758_),
    .C(_0765_),
    .D(_0769_),
    .Y(_0771_));
 sky130_fd_sc_hd__mux4_2 _2437_ (.A0(net264),
    .A1(_0642_),
    .A2(_0747_),
    .A3(_0744_),
    .S0(net240),
    .S1(net245),
    .X(_0772_));
 sky130_fd_sc_hd__inv_2 _2438_ (.A(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__o21a_1 _2439_ (.A1(net286),
    .A2(_0754_),
    .B1(_0637_),
    .X(_0774_));
 sky130_fd_sc_hd__mux4_1 _2440_ (.A0(_0719_),
    .A1(_0722_),
    .A2(_0727_),
    .A3(_0720_),
    .S0(net285),
    .S1(net235),
    .X(_0775_));
 sky130_fd_sc_hd__nor2_1 _2441_ (.A(net277),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__o211a_1 _2442_ (.A1(net286),
    .A2(_0754_),
    .B1(_0637_),
    .C1(net274),
    .X(_0777_));
 sky130_fd_sc_hd__nor2_1 _2443_ (.A(_0776_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__mux4_2 _2444_ (.A0(_0601_),
    .A1(_0636_),
    .A2(_0691_),
    .A3(_0686_),
    .S0(net240),
    .S1(net244),
    .X(_0779_));
 sky130_fd_sc_hd__o211a_1 _2445_ (.A1(_0776_),
    .A2(_0777_),
    .B1(_0779_),
    .C1(_0773_),
    .X(_0780_));
 sky130_fd_sc_hd__nand2_1 _2446_ (.A(_0672_),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__nor2_1 _2447_ (.A(_0771_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__nand2_1 _2448_ (.A(net245),
    .B(_0725_),
    .Y(_0783_));
 sky130_fd_sc_hd__nand2_1 _2449_ (.A(_0631_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__a21oi_1 _2450_ (.A1(net245),
    .A2(_0699_),
    .B1(net170),
    .Y(_0785_));
 sky130_fd_sc_hd__and2_1 _2451_ (.A(_0783_),
    .B(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__nand2_1 _2452_ (.A(_0782_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__or3b_1 _2453_ (.A(_0665_),
    .B(_0667_),
    .C_N(_0786_),
    .X(_0788_));
 sky130_fd_sc_hd__or3_2 _2454_ (.A(_0771_),
    .B(_0781_),
    .C(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__nand2_1 _2455_ (.A(net245),
    .B(_0755_),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_2 _2456_ (.A(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _2457_ (.A(_0631_),
    .B(_0790_),
    .Y(_0792_));
 sky130_fd_sc_hd__o21ai_2 _2458_ (.A1(net278),
    .A2(_0749_),
    .B1(_0631_),
    .Y(_0793_));
 sky130_fd_sc_hd__a21o_1 _2459_ (.A1(net245),
    .A2(_0692_),
    .B1(_0630_),
    .X(_0794_));
 sky130_fd_sc_hd__a21o_1 _2460_ (.A1(net246),
    .A2(_0759_),
    .B1(net170),
    .X(_0795_));
 sky130_fd_sc_hd__a21oi_1 _2461_ (.A1(_0637_),
    .A2(_0761_),
    .B1(net279),
    .Y(_0796_));
 sky130_fd_sc_hd__a21o_1 _2462_ (.A1(net242),
    .A2(_0676_),
    .B1(net170),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_1 _2463_ (.A(net279),
    .B(_0766_),
    .Y(_0798_));
 sky130_fd_sc_hd__o31ai_1 _2464_ (.A1(_0789_),
    .A2(_0791_),
    .A3(_0793_),
    .B1(net271),
    .Y(_0799_));
 sky130_fd_sc_hd__o41a_1 _2465_ (.A1(_0789_),
    .A2(_0791_),
    .A3(_0793_),
    .A4(_0794_),
    .B1(net271),
    .X(_0800_));
 sky130_fd_sc_hd__a21oi_1 _2466_ (.A1(net271),
    .A2(_0652_),
    .B1(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__a21bo_1 _2467_ (.A1(net273),
    .A2(_0795_),
    .B1_N(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__a21o_1 _2468_ (.A1(net273),
    .A2(_0796_),
    .B1(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__a21o_1 _2469_ (.A1(net273),
    .A2(_0797_),
    .B1(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__a21o_1 _2470_ (.A1(net270),
    .A2(_0798_),
    .B1(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__o21a_1 _2471_ (.A1(_0644_),
    .A2(_0805_),
    .B1(net269),
    .X(_0806_));
 sky130_fd_sc_hd__nor2_1 _2472_ (.A(net274),
    .B(_0774_),
    .Y(_0807_));
 sky130_fd_sc_hd__a21oi_1 _2473_ (.A1(net269),
    .A2(_0807_),
    .B1(_0806_),
    .Y(_0808_));
 sky130_fd_sc_hd__xnor2_1 _2474_ (.A(_0639_),
    .B(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(\cordic_inst.cordic_inst.y[30] ),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__or2_1 _2476_ (.A(\cordic_inst.cordic_inst.y[30] ),
    .B(_0809_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2_1 _2477_ (.A(_0810_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__nor2_1 _2478_ (.A(net170),
    .B(_0807_),
    .Y(_0813_));
 sky130_fd_sc_hd__xnor2_1 _2479_ (.A(_0806_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__nor2_1 _2480_ (.A(\cordic_inst.cordic_inst.y[29] ),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__xnor2_1 _2481_ (.A(_0644_),
    .B(_0805_),
    .Y(_0816_));
 sky130_fd_sc_hd__nor2_1 _2482_ (.A(_0595_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__nand2_1 _2483_ (.A(\cordic_inst.cordic_inst.y[29] ),
    .B(_0814_),
    .Y(_0818_));
 sky130_fd_sc_hd__a21oi_1 _2484_ (.A1(\cordic_inst.cordic_inst.y[29] ),
    .A2(_0814_),
    .B1(_0817_),
    .Y(_0819_));
 sky130_fd_sc_hd__and2_1 _2485_ (.A(_0595_),
    .B(_0816_),
    .X(_0820_));
 sky130_fd_sc_hd__or2_1 _2486_ (.A(_0817_),
    .B(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__xnor2_1 _2487_ (.A(_0794_),
    .B(_0799_),
    .Y(_0822_));
 sky130_fd_sc_hd__nand2_1 _2488_ (.A(\cordic_inst.cordic_inst.y[22] ),
    .B(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__or2_1 _2489_ (.A(\cordic_inst.cordic_inst.y[22] ),
    .B(_0822_),
    .X(_0824_));
 sky130_fd_sc_hd__and2_1 _2490_ (.A(_0823_),
    .B(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__nor2_1 _2491_ (.A(_0630_),
    .B(_0652_),
    .Y(_0826_));
 sky130_fd_sc_hd__xnor2_1 _2492_ (.A(_0800_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__nand2_1 _2493_ (.A(\cordic_inst.cordic_inst.y[23] ),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__nor2_1 _2494_ (.A(\cordic_inst.cordic_inst.y[23] ),
    .B(_0827_),
    .Y(_0829_));
 sky130_fd_sc_hd__xnor2_1 _2495_ (.A(\cordic_inst.cordic_inst.y[23] ),
    .B(_0827_),
    .Y(_0830_));
 sky130_fd_sc_hd__inv_2 _2496_ (.A(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__nand2_1 _2497_ (.A(_0825_),
    .B(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_1 _2498_ (.A(net271),
    .B(_0789_),
    .Y(_0833_));
 sky130_fd_sc_hd__xnor2_1 _2499_ (.A(_0793_),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__nand2_1 _2500_ (.A(\cordic_inst.cordic_inst.y[20] ),
    .B(_0834_),
    .Y(_0835_));
 sky130_fd_sc_hd__or2_1 _2501_ (.A(\cordic_inst.cordic_inst.y[20] ),
    .B(_0834_),
    .X(_0836_));
 sky130_fd_sc_hd__nand2_1 _2502_ (.A(_0835_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__o21a_1 _2503_ (.A1(_0789_),
    .A2(_0793_),
    .B1(net271),
    .X(_0838_));
 sky130_fd_sc_hd__xnor2_1 _2504_ (.A(_0792_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__inv_2 _2505_ (.A(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__nand2_1 _2506_ (.A(\cordic_inst.cordic_inst.y[21] ),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__or2_1 _2507_ (.A(\cordic_inst.cordic_inst.y[21] ),
    .B(_0840_),
    .X(_0842_));
 sky130_fd_sc_hd__nand2_1 _2508_ (.A(_0841_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__or3_1 _2509_ (.A(_0832_),
    .B(_0837_),
    .C(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _2510_ (.A(net271),
    .B(_0787_),
    .Y(_0845_));
 sky130_fd_sc_hd__o21a_1 _2511_ (.A1(_0667_),
    .A2(_0787_),
    .B1(net273),
    .X(_0846_));
 sky130_fd_sc_hd__xnor2_1 _2512_ (.A(_0666_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor2_1 _2513_ (.A(\cordic_inst.cordic_inst.y[19] ),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__xor2_1 _2514_ (.A(\cordic_inst.cordic_inst.y[19] ),
    .B(_0847_),
    .X(_0849_));
 sky130_fd_sc_hd__inv_2 _2515_ (.A(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__xor2_1 _2516_ (.A(_0667_),
    .B(_0845_),
    .X(_0851_));
 sky130_fd_sc_hd__or2_1 _2517_ (.A(_0596_),
    .B(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__nand2_1 _2518_ (.A(_0596_),
    .B(_0851_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _2519_ (.A(_0852_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__or2_1 _2520_ (.A(net251),
    .B(_0782_),
    .X(_0855_));
 sky130_fd_sc_hd__a21o_1 _2521_ (.A1(_0782_),
    .A2(_0785_),
    .B1(net251),
    .X(_0856_));
 sky130_fd_sc_hd__xnor2_1 _2522_ (.A(_0784_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__nor2_1 _2523_ (.A(\cordic_inst.cordic_inst.y[17] ),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__xor2_1 _2524_ (.A(_0785_),
    .B(_0855_),
    .X(_0859_));
 sky130_fd_sc_hd__nand2_1 _2525_ (.A(\cordic_inst.cordic_inst.y[16] ),
    .B(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__nand2_1 _2526_ (.A(\cordic_inst.cordic_inst.y[17] ),
    .B(_0857_),
    .Y(_0861_));
 sky130_fd_sc_hd__a21o_1 _2527_ (.A1(_0860_),
    .A2(_0861_),
    .B1(_0858_),
    .X(_0862_));
 sky130_fd_sc_hd__o2bb2a_1 _2528_ (.A1_N(\cordic_inst.cordic_inst.y[19] ),
    .A2_N(_0847_),
    .B1(_0851_),
    .B2(_0596_),
    .X(_0863_));
 sky130_fd_sc_hd__o32a_1 _2529_ (.A1(_0850_),
    .A2(_0854_),
    .A3(_0862_),
    .B1(_0863_),
    .B2(_0848_),
    .X(_0864_));
 sky130_fd_sc_hd__a21bo_1 _2530_ (.A1(_0835_),
    .A2(_0841_),
    .B1_N(_0842_),
    .X(_0865_));
 sky130_fd_sc_hd__a21o_1 _2531_ (.A1(_0823_),
    .A2(_0828_),
    .B1(_0829_),
    .X(_0866_));
 sky130_fd_sc_hd__o221a_1 _2532_ (.A1(_0844_),
    .A2(_0864_),
    .B1(_0865_),
    .B2(_0832_),
    .C1(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__and2b_1 _2533_ (.A_N(_0858_),
    .B(_0861_),
    .X(_0868_));
 sky130_fd_sc_hd__or3b_1 _2534_ (.A(_0850_),
    .B(_0854_),
    .C_N(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__a21oi_1 _2535_ (.A1(_0743_),
    .A2(_0757_),
    .B1(net250),
    .Y(_0870_));
 sky130_fd_sc_hd__a31o_1 _2536_ (.A1(_0693_),
    .A2(_0743_),
    .A3(_0757_),
    .B1(net250),
    .X(_0871_));
 sky130_fd_sc_hd__xor2_1 _2537_ (.A(_0684_),
    .B(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__and2_1 _2538_ (.A(\cordic_inst.cordic_inst.y[7] ),
    .B(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__nor2_1 _2539_ (.A(\cordic_inst.cordic_inst.y[7] ),
    .B(_0872_),
    .Y(_0874_));
 sky130_fd_sc_hd__xnor2_1 _2540_ (.A(_0693_),
    .B(_0870_),
    .Y(_0875_));
 sky130_fd_sc_hd__nor2_1 _2541_ (.A(\cordic_inst.cordic_inst.y[6] ),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__inv_2 _2542_ (.A(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__nand2_1 _2543_ (.A(\cordic_inst.cordic_inst.y[6] ),
    .B(_0875_),
    .Y(_0878_));
 sky130_fd_sc_hd__inv_2 _2544_ (.A(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nor2_1 _2545_ (.A(net250),
    .B(_0743_),
    .Y(_0880_));
 sky130_fd_sc_hd__a21o_1 _2546_ (.A1(_0743_),
    .A2(_0750_),
    .B1(net250),
    .X(_0881_));
 sky130_fd_sc_hd__xnor2_1 _2547_ (.A(_0756_),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__and2_1 _2548_ (.A(_0599_),
    .B(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__nand2_1 _2549_ (.A(_0599_),
    .B(_0882_),
    .Y(_0884_));
 sky130_fd_sc_hd__nor2_1 _2550_ (.A(_0599_),
    .B(_0882_),
    .Y(_0885_));
 sky130_fd_sc_hd__xnor2_1 _2551_ (.A(_0750_),
    .B(_0880_),
    .Y(_0886_));
 sky130_fd_sc_hd__o31a_1 _2552_ (.A1(_0718_),
    .A2(_0735_),
    .A3(_0738_),
    .B1(net272),
    .X(_0887_));
 sky130_fd_sc_hd__xnor2_1 _2553_ (.A(_0742_),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__and2_1 _2554_ (.A(\cordic_inst.cordic_inst.y[3] ),
    .B(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__o21ai_1 _2555_ (.A1(_0718_),
    .A2(_0735_),
    .B1(net272),
    .Y(_0890_));
 sky130_fd_sc_hd__xnor2_1 _2556_ (.A(_0738_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__and2_1 _2557_ (.A(\cordic_inst.cordic_inst.y[2] ),
    .B(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__o211a_1 _2558_ (.A1(net247),
    .A2(_0699_),
    .B1(_0717_),
    .C1(net272),
    .X(_0893_));
 sky130_fd_sc_hd__xor2_1 _2559_ (.A(_0735_),
    .B(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__nand2_1 _2560_ (.A(\cordic_inst.cordic_inst.y[1] ),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand2_1 _2561_ (.A(\cordic_inst.cordic_inst.y[0] ),
    .B(_0718_),
    .Y(_0896_));
 sky130_fd_sc_hd__xnor2_1 _2562_ (.A(\cordic_inst.cordic_inst.y[1] ),
    .B(_0894_),
    .Y(_0897_));
 sky130_fd_sc_hd__or2_1 _2563_ (.A(_0896_),
    .B(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__o21ai_1 _2564_ (.A1(_0896_),
    .A2(_0897_),
    .B1(_0895_),
    .Y(_0899_));
 sky130_fd_sc_hd__xor2_1 _2565_ (.A(\cordic_inst.cordic_inst.y[2] ),
    .B(_0891_),
    .X(_0900_));
 sky130_fd_sc_hd__nand2_1 _2566_ (.A(_0899_),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__a21o_1 _2567_ (.A1(_0899_),
    .A2(_0900_),
    .B1(_0892_),
    .X(_0902_));
 sky130_fd_sc_hd__nor2_1 _2568_ (.A(\cordic_inst.cordic_inst.y[3] ),
    .B(_0888_),
    .Y(_0903_));
 sky130_fd_sc_hd__nor2_1 _2569_ (.A(_0889_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand2_1 _2570_ (.A(_0902_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__a21o_1 _2571_ (.A1(_0902_),
    .A2(_0904_),
    .B1(_0889_),
    .X(_0906_));
 sky130_fd_sc_hd__xor2_1 _2572_ (.A(\cordic_inst.cordic_inst.y[4] ),
    .B(_0886_),
    .X(_0907_));
 sky130_fd_sc_hd__and2_1 _2573_ (.A(_0906_),
    .B(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__inv_2 _2574_ (.A(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21o_1 _2575_ (.A1(\cordic_inst.cordic_inst.y[4] ),
    .A2(_0886_),
    .B1(_0908_),
    .X(_0910_));
 sky130_fd_sc_hd__a31o_1 _2576_ (.A1(\cordic_inst.cordic_inst.y[4] ),
    .A2(_0884_),
    .A3(_0886_),
    .B1(_0885_),
    .X(_0911_));
 sky130_fd_sc_hd__nor2_1 _2577_ (.A(_0883_),
    .B(_0885_),
    .Y(_0912_));
 sky130_fd_sc_hd__a31o_1 _2578_ (.A1(_0906_),
    .A2(_0907_),
    .A3(_0912_),
    .B1(_0911_),
    .X(_0913_));
 sky130_fd_sc_hd__o221a_1 _2579_ (.A1(\cordic_inst.cordic_inst.y[7] ),
    .A2(_0872_),
    .B1(_0879_),
    .B2(_0913_),
    .C1(_0877_),
    .X(_0914_));
 sky130_fd_sc_hd__nor2_1 _2580_ (.A(_0873_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__a21oi_1 _2581_ (.A1(_0770_),
    .A2(_0780_),
    .B1(net251),
    .Y(_0916_));
 sky130_fd_sc_hd__xnor2_2 _2582_ (.A(_0672_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__nand2_1 _2583_ (.A(\cordic_inst.cordic_inst.y[15] ),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__nor2_1 _2584_ (.A(\cordic_inst.cordic_inst.y[15] ),
    .B(_0917_),
    .Y(_0919_));
 sky130_fd_sc_hd__xnor2_1 _2585_ (.A(\cordic_inst.cordic_inst.y[15] ),
    .B(_0917_),
    .Y(_0920_));
 sky130_fd_sc_hd__nor2_1 _2586_ (.A(net250),
    .B(_0770_),
    .Y(_0921_));
 sky130_fd_sc_hd__o31ai_2 _2587_ (.A1(_0771_),
    .A2(_0772_),
    .A3(_0778_),
    .B1(net271),
    .Y(_0922_));
 sky130_fd_sc_hd__xor2_2 _2588_ (.A(_0779_),
    .B(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _2589_ (.A(\cordic_inst.cordic_inst.y[14] ),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__xnor2_1 _2590_ (.A(\cordic_inst.cordic_inst.y[14] ),
    .B(_0923_),
    .Y(_0925_));
 sky130_fd_sc_hd__or2_1 _2591_ (.A(_0920_),
    .B(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__xnor2_1 _2592_ (.A(_0772_),
    .B(_0921_),
    .Y(_0927_));
 sky130_fd_sc_hd__and2b_1 _2593_ (.A_N(_0927_),
    .B(\cordic_inst.cordic_inst.y[12] ),
    .X(_0928_));
 sky130_fd_sc_hd__and2b_1 _2594_ (.A_N(\cordic_inst.cordic_inst.y[12] ),
    .B(_0927_),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_1 _2595_ (.A(_0928_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__a21o_1 _2596_ (.A1(_0770_),
    .A2(_0773_),
    .B1(net250),
    .X(_0931_));
 sky130_fd_sc_hd__xnor2_1 _2597_ (.A(_0778_),
    .B(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__nor2_1 _2598_ (.A(\cordic_inst.cordic_inst.y[13] ),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__and2_1 _2599_ (.A(\cordic_inst.cordic_inst.y[13] ),
    .B(_0932_),
    .X(_0934_));
 sky130_fd_sc_hd__nor2_1 _2600_ (.A(_0933_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__nand3b_1 _2601_ (.A_N(_0926_),
    .B(_0930_),
    .C(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__a31o_1 _2602_ (.A1(net154),
    .A2(_0758_),
    .A3(_0765_),
    .B1(net250),
    .X(_0937_));
 sky130_fd_sc_hd__xnor2_1 _2603_ (.A(_0769_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__nand2b_1 _2604_ (.A_N(\cordic_inst.cordic_inst.y[11] ),
    .B(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__inv_2 _2605_ (.A(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__and2b_1 _2606_ (.A_N(_0938_),
    .B(\cordic_inst.cordic_inst.y[11] ),
    .X(_0941_));
 sky130_fd_sc_hd__nor2_1 _2607_ (.A(_0940_),
    .B(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__a31o_1 _2608_ (.A1(net154),
    .A2(_0758_),
    .A3(_0764_),
    .B1(net250),
    .X(_0943_));
 sky130_fd_sc_hd__xor2_1 _2609_ (.A(_0677_),
    .B(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__nor2_1 _2610_ (.A(_0597_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__and2_1 _2611_ (.A(_0597_),
    .B(_0944_),
    .X(_0946_));
 sky130_fd_sc_hd__or2_1 _2612_ (.A(_0945_),
    .B(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__or3_1 _2613_ (.A(_0940_),
    .B(_0941_),
    .C(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__a21oi_1 _2614_ (.A1(net154),
    .A2(_0758_),
    .B1(net250),
    .Y(_0949_));
 sky130_fd_sc_hd__a21oi_1 _2615_ (.A1(net271),
    .A2(_0760_),
    .B1(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__xnor2_1 _2616_ (.A(_0762_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _2617_ (.A(\cordic_inst.cordic_inst.y[9] ),
    .B(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2_1 _2618_ (.A(\cordic_inst.cordic_inst.y[9] ),
    .B(_0951_),
    .Y(_0953_));
 sky130_fd_sc_hd__inv_2 _2619_ (.A(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__nand2_1 _2620_ (.A(_0952_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__xnor2_1 _2621_ (.A(_0760_),
    .B(_0949_),
    .Y(_0956_));
 sky130_fd_sc_hd__or2_1 _2622_ (.A(_0598_),
    .B(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__nand2_1 _2623_ (.A(_0598_),
    .B(_0956_),
    .Y(_0958_));
 sky130_fd_sc_hd__nand2_1 _2624_ (.A(_0957_),
    .B(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__or4_1 _2625_ (.A(_0936_),
    .B(_0948_),
    .C(_0955_),
    .D(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__or2_1 _2626_ (.A(_0915_),
    .B(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__o21a_1 _2627_ (.A1(_0953_),
    .A2(_0957_),
    .B1(_0952_),
    .X(_0962_));
 sky130_fd_sc_hd__or2_1 _2628_ (.A(_0941_),
    .B(_0945_),
    .X(_0963_));
 sky130_fd_sc_hd__o2bb2a_1 _2629_ (.A1_N(_0939_),
    .A2_N(_0963_),
    .B1(_0962_),
    .B2(_0948_),
    .X(_0964_));
 sky130_fd_sc_hd__a21oi_1 _2630_ (.A1(\cordic_inst.cordic_inst.y[13] ),
    .A2(_0932_),
    .B1(_0928_),
    .Y(_0965_));
 sky130_fd_sc_hd__a21o_1 _2631_ (.A1(_0918_),
    .A2(_0924_),
    .B1(_0919_),
    .X(_0966_));
 sky130_fd_sc_hd__o32a_1 _2632_ (.A1(_0926_),
    .A2(_0933_),
    .A3(_0965_),
    .B1(_0964_),
    .B2(_0936_),
    .X(_0967_));
 sky130_fd_sc_hd__and3_1 _2633_ (.A(_0961_),
    .B(_0966_),
    .C(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__or2_1 _2634_ (.A(\cordic_inst.cordic_inst.y[16] ),
    .B(_0859_),
    .X(_0969_));
 sky130_fd_sc_hd__nand2_1 _2635_ (.A(_0860_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_1 _2636_ (.A(_0968_),
    .B(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__inv_2 _2637_ (.A(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__or3_1 _2638_ (.A(_0869_),
    .B(_0968_),
    .C(_0970_),
    .X(_0973_));
 sky130_fd_sc_hd__o41a_1 _2639_ (.A1(_0844_),
    .A2(_0869_),
    .A3(_0968_),
    .A4(_0970_),
    .B1(_0867_),
    .X(_0974_));
 sky130_fd_sc_hd__xnor2_1 _2640_ (.A(_0795_),
    .B(_0801_),
    .Y(_0975_));
 sky130_fd_sc_hd__and2_1 _2641_ (.A(\cordic_inst.cordic_inst.y[24] ),
    .B(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__nor2_1 _2642_ (.A(\cordic_inst.cordic_inst.y[24] ),
    .B(_0975_),
    .Y(_0977_));
 sky130_fd_sc_hd__or2_1 _2643_ (.A(_0976_),
    .B(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_1 _2644_ (.A(_0974_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__nor2_1 _2645_ (.A(net170),
    .B(_0798_),
    .Y(_0980_));
 sky130_fd_sc_hd__xnor2_1 _2646_ (.A(_0804_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__nor2_1 _2647_ (.A(\cordic_inst.cordic_inst.y[27] ),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_1 _2648_ (.A(\cordic_inst.cordic_inst.y[27] ),
    .B(_0981_),
    .Y(_0983_));
 sky130_fd_sc_hd__and2b_1 _2649_ (.A_N(_0982_),
    .B(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__xor2_1 _2650_ (.A(_0797_),
    .B(_0803_),
    .X(_0985_));
 sky130_fd_sc_hd__xor2_1 _2651_ (.A(\cordic_inst.cordic_inst.y[26] ),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__nor2_1 _2652_ (.A(net170),
    .B(_0796_),
    .Y(_0987_));
 sky130_fd_sc_hd__xnor2_1 _2653_ (.A(_0802_),
    .B(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__or2_1 _2654_ (.A(\cordic_inst.cordic_inst.y[25] ),
    .B(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__nand2_1 _2655_ (.A(\cordic_inst.cordic_inst.y[25] ),
    .B(_0988_),
    .Y(_0990_));
 sky130_fd_sc_hd__and4_1 _2656_ (.A(_0984_),
    .B(_0986_),
    .C(_0989_),
    .D(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_1 _2657_ (.A(_0979_),
    .B(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__a21o_1 _2658_ (.A1(\cordic_inst.cordic_inst.y[25] ),
    .A2(_0988_),
    .B1(_0976_),
    .X(_0993_));
 sky130_fd_sc_hd__nand4_1 _2659_ (.A(_0984_),
    .B(_0986_),
    .C(_0989_),
    .D(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand3b_1 _2660_ (.A_N(_0982_),
    .B(_0985_),
    .C(\cordic_inst.cordic_inst.y[26] ),
    .Y(_0995_));
 sky130_fd_sc_hd__and4_1 _2661_ (.A(_0983_),
    .B(_0992_),
    .C(_0994_),
    .D(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__a41o_1 _2662_ (.A1(_0983_),
    .A2(_0992_),
    .A3(_0994_),
    .A4(_0995_),
    .B1(_0821_),
    .X(_0997_));
 sky130_fd_sc_hd__and2b_1 _2663_ (.A_N(_0815_),
    .B(_0818_),
    .X(_0998_));
 sky130_fd_sc_hd__a21o_1 _2664_ (.A1(_0819_),
    .A2(_0997_),
    .B1(_0815_),
    .X(_0999_));
 sky130_fd_sc_hd__a211o_1 _2665_ (.A1(_0819_),
    .A2(_0997_),
    .B1(_0812_),
    .C1(_0815_),
    .X(_1000_));
 sky130_fd_sc_hd__o31a_1 _2666_ (.A1(_0639_),
    .A2(_0806_),
    .A3(_0807_),
    .B1(net269),
    .X(_1001_));
 sky130_fd_sc_hd__xnor2_2 _2667_ (.A(net263),
    .B(net265),
    .Y(_1002_));
 sky130_fd_sc_hd__xor2_1 _2668_ (.A(_1001_),
    .B(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__a21oi_1 _2669_ (.A1(_0810_),
    .A2(_1000_),
    .B1(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__a31o_1 _2670_ (.A1(_0810_),
    .A2(_1000_),
    .A3(_1003_),
    .B1(net176),
    .X(_1005_));
 sky130_fd_sc_hd__a2bb2o_1 _2671_ (.A1_N(_1004_),
    .A2_N(_1005_),
    .B1(net263),
    .B2(net164),
    .X(_0561_));
 sky130_fd_sc_hd__nand2_1 _2672_ (.A(_0812_),
    .B(_0999_),
    .Y(_1006_));
 sky130_fd_sc_hd__a32o_1 _2673_ (.A1(net181),
    .A2(_1000_),
    .A3(_1006_),
    .B1(net164),
    .B2(\cordic_inst.cordic_inst.y[30] ),
    .X(_0560_));
 sky130_fd_sc_hd__and2b_1 _2674_ (.A_N(_0817_),
    .B(_0997_),
    .X(_1007_));
 sky130_fd_sc_hd__xnor2_1 _2675_ (.A(_0998_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__a22o_1 _2676_ (.A1(\cordic_inst.cordic_inst.y[29] ),
    .A2(net163),
    .B1(_1008_),
    .B2(net182),
    .X(_0559_));
 sky130_fd_sc_hd__nand2_1 _2677_ (.A(_0821_),
    .B(_0996_),
    .Y(_1009_));
 sky130_fd_sc_hd__a32o_1 _2678_ (.A1(net182),
    .A2(_0997_),
    .A3(_1009_),
    .B1(net163),
    .B2(\cordic_inst.cordic_inst.y[28] ),
    .X(_0558_));
 sky130_fd_sc_hd__or2_1 _2679_ (.A(_0976_),
    .B(_0979_),
    .X(_1010_));
 sky130_fd_sc_hd__o21a_1 _2680_ (.A1(_0979_),
    .A2(_0993_),
    .B1(_0989_),
    .X(_1011_));
 sky130_fd_sc_hd__and2_1 _2681_ (.A(_0986_),
    .B(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__a21oi_1 _2682_ (.A1(\cordic_inst.cordic_inst.y[26] ),
    .A2(_0985_),
    .B1(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__xnor2_1 _2683_ (.A(_0984_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__a22o_1 _2684_ (.A1(\cordic_inst.cordic_inst.y[27] ),
    .A2(net163),
    .B1(_1014_),
    .B2(net181),
    .X(_0557_));
 sky130_fd_sc_hd__or2_1 _2685_ (.A(_0986_),
    .B(_1011_),
    .X(_1015_));
 sky130_fd_sc_hd__nor2_1 _2686_ (.A(net176),
    .B(_1012_),
    .Y(_1016_));
 sky130_fd_sc_hd__a22o_1 _2687_ (.A1(\cordic_inst.cordic_inst.y[26] ),
    .A2(net169),
    .B1(_1015_),
    .B2(_1016_),
    .X(_0556_));
 sky130_fd_sc_hd__nand3_1 _2688_ (.A(_0989_),
    .B(_0990_),
    .C(_1010_),
    .Y(_1017_));
 sky130_fd_sc_hd__a21o_1 _2689_ (.A1(_0989_),
    .A2(_0990_),
    .B1(_1010_),
    .X(_1018_));
 sky130_fd_sc_hd__a32o_1 _2690_ (.A1(net186),
    .A2(_1017_),
    .A3(_1018_),
    .B1(net169),
    .B2(\cordic_inst.cordic_inst.y[25] ),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _2691_ (.A(_0974_),
    .B(_0978_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _2692_ (.A(net177),
    .B(_0979_),
    .Y(_1020_));
 sky130_fd_sc_hd__a22o_1 _2693_ (.A1(\cordic_inst.cordic_inst.y[24] ),
    .A2(net169),
    .B1(_1019_),
    .B2(_1020_),
    .X(_0554_));
 sky130_fd_sc_hd__a21o_1 _2694_ (.A1(_0864_),
    .A2(_0973_),
    .B1(_0837_),
    .X(_1021_));
 sky130_fd_sc_hd__nand2_1 _2695_ (.A(_0835_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__a21bo_1 _2696_ (.A1(_0842_),
    .A2(_1022_),
    .B1_N(_0841_),
    .X(_1023_));
 sky130_fd_sc_hd__a21bo_1 _2697_ (.A1(_0825_),
    .A2(_1023_),
    .B1_N(_0823_),
    .X(_1024_));
 sky130_fd_sc_hd__xnor2_1 _2698_ (.A(_0830_),
    .B(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__a22o_1 _2699_ (.A1(\cordic_inst.cordic_inst.y[23] ),
    .A2(net165),
    .B1(_1025_),
    .B2(net186),
    .X(_0553_));
 sky130_fd_sc_hd__xor2_1 _2700_ (.A(_0825_),
    .B(_1023_),
    .X(_1026_));
 sky130_fd_sc_hd__a22o_1 _2701_ (.A1(\cordic_inst.cordic_inst.y[22] ),
    .A2(net165),
    .B1(_1026_),
    .B2(net183),
    .X(_0552_));
 sky130_fd_sc_hd__xnor2_1 _2702_ (.A(_0843_),
    .B(_1022_),
    .Y(_1027_));
 sky130_fd_sc_hd__a22o_1 _2703_ (.A1(\cordic_inst.cordic_inst.y[21] ),
    .A2(net165),
    .B1(_1027_),
    .B2(net183),
    .X(_0551_));
 sky130_fd_sc_hd__nand3_1 _2704_ (.A(_0837_),
    .B(_0864_),
    .C(_0973_),
    .Y(_1028_));
 sky130_fd_sc_hd__a32o_1 _2705_ (.A1(net183),
    .A2(_1021_),
    .A3(_1028_),
    .B1(net167),
    .B2(\cordic_inst.cordic_inst.y[20] ),
    .X(_0550_));
 sky130_fd_sc_hd__and3_1 _2706_ (.A(_0860_),
    .B(_0861_),
    .C(_0972_),
    .X(_1029_));
 sky130_fd_sc_hd__or3_1 _2707_ (.A(_0854_),
    .B(_0858_),
    .C(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__a21oi_1 _2708_ (.A1(_0852_),
    .A2(_1030_),
    .B1(_0850_),
    .Y(_1031_));
 sky130_fd_sc_hd__a31o_1 _2709_ (.A1(_0850_),
    .A2(_0852_),
    .A3(_1030_),
    .B1(net177),
    .X(_1032_));
 sky130_fd_sc_hd__a2bb2o_1 _2710_ (.A1_N(_1031_),
    .A2_N(_1032_),
    .B1(\cordic_inst.cordic_inst.y[19] ),
    .B2(net167),
    .X(_0549_));
 sky130_fd_sc_hd__o21ai_1 _2711_ (.A1(_0858_),
    .A2(_1029_),
    .B1(_0854_),
    .Y(_1033_));
 sky130_fd_sc_hd__a32o_1 _2712_ (.A1(net186),
    .A2(_1030_),
    .A3(_1033_),
    .B1(net167),
    .B2(\cordic_inst.cordic_inst.y[18] ),
    .X(_0548_));
 sky130_fd_sc_hd__nand2_1 _2713_ (.A(_0860_),
    .B(_0972_),
    .Y(_1034_));
 sky130_fd_sc_hd__xor2_1 _2714_ (.A(_0868_),
    .B(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__a22o_1 _2715_ (.A1(\cordic_inst.cordic_inst.y[17] ),
    .A2(net166),
    .B1(_1035_),
    .B2(net184),
    .X(_0547_));
 sky130_fd_sc_hd__nand2_1 _2716_ (.A(_0968_),
    .B(_0970_),
    .Y(_1036_));
 sky130_fd_sc_hd__a32o_1 _2717_ (.A1(net184),
    .A2(_0972_),
    .A3(_1036_),
    .B1(net167),
    .B2(\cordic_inst.cordic_inst.y[16] ),
    .X(_0546_));
 sky130_fd_sc_hd__or2_1 _2718_ (.A(_0915_),
    .B(_0959_),
    .X(_1037_));
 sky130_fd_sc_hd__o21a_1 _2719_ (.A1(_0955_),
    .A2(_1037_),
    .B1(_0962_),
    .X(_1038_));
 sky130_fd_sc_hd__nor2_1 _2720_ (.A(_0947_),
    .B(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__o21a_1 _2721_ (.A1(_0963_),
    .A2(_1039_),
    .B1(_0939_),
    .X(_1040_));
 sky130_fd_sc_hd__o211ai_2 _2722_ (.A1(_0963_),
    .A2(_1039_),
    .B1(_0930_),
    .C1(_0939_),
    .Y(_1041_));
 sky130_fd_sc_hd__a21o_1 _2723_ (.A1(_0965_),
    .A2(_1041_),
    .B1(_0933_),
    .X(_1042_));
 sky130_fd_sc_hd__or2_1 _2724_ (.A(_0925_),
    .B(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__a21bo_1 _2725_ (.A1(\cordic_inst.cordic_inst.y[14] ),
    .A2(_0923_),
    .B1_N(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__xnor2_1 _2726_ (.A(_0920_),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a22o_1 _2727_ (.A1(\cordic_inst.cordic_inst.y[15] ),
    .A2(net166),
    .B1(_1045_),
    .B2(net184),
    .X(_0545_));
 sky130_fd_sc_hd__nand2_1 _2728_ (.A(_0925_),
    .B(_1042_),
    .Y(_1046_));
 sky130_fd_sc_hd__a32o_1 _2729_ (.A1(net184),
    .A2(_1043_),
    .A3(_1046_),
    .B1(net166),
    .B2(\cordic_inst.cordic_inst.y[14] ),
    .X(_0544_));
 sky130_fd_sc_hd__and2b_1 _2730_ (.A_N(_0928_),
    .B(_1041_),
    .X(_1047_));
 sky130_fd_sc_hd__xnor2_1 _2731_ (.A(_0935_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__a22o_1 _2732_ (.A1(\cordic_inst.cordic_inst.y[13] ),
    .A2(net166),
    .B1(_1048_),
    .B2(net184),
    .X(_0543_));
 sky130_fd_sc_hd__or2_1 _2733_ (.A(_0930_),
    .B(_1040_),
    .X(_1049_));
 sky130_fd_sc_hd__a32o_1 _2734_ (.A1(net184),
    .A2(_1041_),
    .A3(_1049_),
    .B1(net166),
    .B2(\cordic_inst.cordic_inst.y[12] ),
    .X(_0542_));
 sky130_fd_sc_hd__o21ai_1 _2735_ (.A1(_0945_),
    .A2(_1039_),
    .B1(_0942_),
    .Y(_1050_));
 sky130_fd_sc_hd__or3_1 _2736_ (.A(_0942_),
    .B(_0945_),
    .C(_1039_),
    .X(_1051_));
 sky130_fd_sc_hd__a32o_1 _2737_ (.A1(net184),
    .A2(_1050_),
    .A3(_1051_),
    .B1(net166),
    .B2(\cordic_inst.cordic_inst.y[11] ),
    .X(_0541_));
 sky130_fd_sc_hd__nand2_1 _2738_ (.A(_0947_),
    .B(_1038_),
    .Y(_1052_));
 sky130_fd_sc_hd__nor2_1 _2739_ (.A(net177),
    .B(_1039_),
    .Y(_1053_));
 sky130_fd_sc_hd__a22o_1 _2740_ (.A1(\cordic_inst.cordic_inst.y[10] ),
    .A2(net166),
    .B1(_1052_),
    .B2(_1053_),
    .X(_0540_));
 sky130_fd_sc_hd__nand3_1 _2741_ (.A(_0955_),
    .B(_0957_),
    .C(_1037_),
    .Y(_1054_));
 sky130_fd_sc_hd__a21o_1 _2742_ (.A1(_0957_),
    .A2(_1037_),
    .B1(_0955_),
    .X(_1055_));
 sky130_fd_sc_hd__a32o_1 _2743_ (.A1(net184),
    .A2(_1054_),
    .A3(_1055_),
    .B1(net166),
    .B2(\cordic_inst.cordic_inst.y[9] ),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_1 _2744_ (.A(_0915_),
    .B(_0959_),
    .Y(_1056_));
 sky130_fd_sc_hd__a32o_1 _2745_ (.A1(net185),
    .A2(_1037_),
    .A3(_1056_),
    .B1(net166),
    .B2(\cordic_inst.cordic_inst.y[8] ),
    .X(_0538_));
 sky130_fd_sc_hd__or3b_1 _2746_ (.A(_0876_),
    .B(_0879_),
    .C_N(_0913_),
    .X(_1057_));
 sky130_fd_sc_hd__o211ai_1 _2747_ (.A1(_0873_),
    .A2(_0874_),
    .B1(_0878_),
    .C1(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__nand2b_1 _2748_ (.A_N(_0873_),
    .B(_0914_),
    .Y(_1059_));
 sky130_fd_sc_hd__a32o_1 _2749_ (.A1(net185),
    .A2(_1058_),
    .A3(_1059_),
    .B1(net168),
    .B2(\cordic_inst.cordic_inst.y[7] ),
    .X(_0537_));
 sky130_fd_sc_hd__a21o_1 _2750_ (.A1(_0877_),
    .A2(_0878_),
    .B1(_0913_),
    .X(_1060_));
 sky130_fd_sc_hd__a32o_1 _2751_ (.A1(net185),
    .A2(_1057_),
    .A3(_1060_),
    .B1(net168),
    .B2(\cordic_inst.cordic_inst.y[6] ),
    .X(_0536_));
 sky130_fd_sc_hd__xor2_1 _2752_ (.A(_0910_),
    .B(_0912_),
    .X(_1061_));
 sky130_fd_sc_hd__a22o_1 _2753_ (.A1(\cordic_inst.cordic_inst.y[5] ),
    .A2(net168),
    .B1(_1061_),
    .B2(net185),
    .X(_0535_));
 sky130_fd_sc_hd__or2_1 _2754_ (.A(_0906_),
    .B(_0907_),
    .X(_1062_));
 sky130_fd_sc_hd__a32o_1 _2755_ (.A1(net185),
    .A2(_0909_),
    .A3(_1062_),
    .B1(net168),
    .B2(\cordic_inst.cordic_inst.y[4] ),
    .X(_0534_));
 sky130_fd_sc_hd__or2_1 _2756_ (.A(_0902_),
    .B(_0904_),
    .X(_1063_));
 sky130_fd_sc_hd__a32o_1 _2757_ (.A1(net185),
    .A2(_0905_),
    .A3(_1063_),
    .B1(net168),
    .B2(\cordic_inst.cordic_inst.y[3] ),
    .X(_0533_));
 sky130_fd_sc_hd__or2_1 _2758_ (.A(_0899_),
    .B(_0900_),
    .X(_1064_));
 sky130_fd_sc_hd__a32o_1 _2759_ (.A1(net183),
    .A2(_0901_),
    .A3(_1064_),
    .B1(net165),
    .B2(\cordic_inst.cordic_inst.y[2] ),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_1 _2760_ (.A(_0896_),
    .B(_0897_),
    .Y(_1065_));
 sky130_fd_sc_hd__a32o_1 _2761_ (.A1(net183),
    .A2(_0898_),
    .A3(_1065_),
    .B1(net165),
    .B2(\cordic_inst.cordic_inst.y[1] ),
    .X(_0531_));
 sky130_fd_sc_hd__nand2_1 _2762_ (.A(net183),
    .B(_0718_),
    .Y(_1066_));
 sky130_fd_sc_hd__nor2_1 _2763_ (.A(_0600_),
    .B(net173),
    .Y(_1067_));
 sky130_fd_sc_hd__mux2_1 _2764_ (.A0(_0600_),
    .A1(_1067_),
    .S(_1066_),
    .X(_0530_));
 sky130_fd_sc_hd__and2_1 _2765_ (.A(net263),
    .B(net274),
    .X(_1068_));
 sky130_fd_sc_hd__nand2_1 _2766_ (.A(net262),
    .B(net276),
    .Y(_1069_));
 sky130_fd_sc_hd__nand2_2 _2767_ (.A(net263),
    .B(net282),
    .Y(_1070_));
 sky130_fd_sc_hd__and2_1 _2768_ (.A(net263),
    .B(net293),
    .X(_1071_));
 sky130_fd_sc_hd__and2_1 _2769_ (.A(net263),
    .B(net295),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _2770_ (.A0(\cordic_inst.cordic_inst.y[30] ),
    .A1(net263),
    .S(net306),
    .X(_1073_));
 sky130_fd_sc_hd__a21o_1 _2771_ (.A1(net232),
    .A2(_1073_),
    .B1(_1072_),
    .X(_1074_));
 sky130_fd_sc_hd__a21o_1 _2772_ (.A1(net237),
    .A2(_1074_),
    .B1(_1071_),
    .X(_1075_));
 sky130_fd_sc_hd__a21bo_1 _2773_ (.A1(net241),
    .A2(_1075_),
    .B1_N(_1070_),
    .X(_1076_));
 sky130_fd_sc_hd__a21o_1 _2774_ (.A1(net242),
    .A2(_1076_),
    .B1(net215),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(\cordic_inst.cordic_inst.y[28] ),
    .A1(\cordic_inst.cordic_inst.y[29] ),
    .S(net306),
    .X(_1078_));
 sky130_fd_sc_hd__mux4_2 _2776_ (.A0(\cordic_inst.cordic_inst.y[28] ),
    .A1(\cordic_inst.cordic_inst.y[29] ),
    .A2(\cordic_inst.cordic_inst.y[30] ),
    .A3(net263),
    .S0(net304),
    .S1(net295),
    .X(_1079_));
 sky130_fd_sc_hd__a21o_1 _2777_ (.A1(net237),
    .A2(_1079_),
    .B1(_1071_),
    .X(_1080_));
 sky130_fd_sc_hd__a21bo_1 _2778_ (.A1(net241),
    .A2(_1080_),
    .B1_N(_1070_),
    .X(_1081_));
 sky130_fd_sc_hd__a21o_1 _2779_ (.A1(net242),
    .A2(_1081_),
    .B1(net215),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _2780_ (.A0(\cordic_inst.cordic_inst.y[25] ),
    .A1(\cordic_inst.cordic_inst.y[26] ),
    .S(net304),
    .X(_1083_));
 sky130_fd_sc_hd__mux4_1 _2781_ (.A0(\cordic_inst.cordic_inst.y[23] ),
    .A1(\cordic_inst.cordic_inst.y[24] ),
    .A2(\cordic_inst.cordic_inst.y[25] ),
    .A3(\cordic_inst.cordic_inst.y[26] ),
    .S0(net307),
    .S1(net301),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _2782_ (.A0(\cordic_inst.cordic_inst.y[27] ),
    .A1(\cordic_inst.cordic_inst.y[28] ),
    .S(net304),
    .X(_1085_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(\cordic_inst.cordic_inst.y[29] ),
    .A1(\cordic_inst.cordic_inst.y[30] ),
    .S(net304),
    .X(_1086_));
 sky130_fd_sc_hd__mux4_1 _2784_ (.A0(\cordic_inst.cordic_inst.y[27] ),
    .A1(\cordic_inst.cordic_inst.y[28] ),
    .A2(\cordic_inst.cordic_inst.y[29] ),
    .A3(\cordic_inst.cordic_inst.y[30] ),
    .S0(net304),
    .S1(net295),
    .X(_1087_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(_1084_),
    .A1(_1087_),
    .S(net291),
    .X(_1088_));
 sky130_fd_sc_hd__a21boi_1 _2786_ (.A1(net238),
    .A2(_1088_),
    .B1_N(_1070_),
    .Y(_1089_));
 sky130_fd_sc_hd__nor2_1 _2787_ (.A(net274),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__a21o_1 _2788_ (.A1(net233),
    .A2(_1087_),
    .B1(_1071_),
    .X(_1091_));
 sky130_fd_sc_hd__nand2_1 _2789_ (.A(net241),
    .B(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__mux4_1 _2790_ (.A0(\cordic_inst.cordic_inst.y[19] ),
    .A1(\cordic_inst.cordic_inst.y[20] ),
    .A2(\cordic_inst.cordic_inst.y[21] ),
    .A3(\cordic_inst.cordic_inst.y[22] ),
    .S0(net307),
    .S1(net300),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(_1084_),
    .A1(_1093_),
    .S(net235),
    .X(_1094_));
 sky130_fd_sc_hd__mux4_1 _2792_ (.A0(\cordic_inst.cordic_inst.y[11] ),
    .A1(\cordic_inst.cordic_inst.y[12] ),
    .A2(\cordic_inst.cordic_inst.y[13] ),
    .A3(\cordic_inst.cordic_inst.y[14] ),
    .S0(net310),
    .S1(net299),
    .X(_1095_));
 sky130_fd_sc_hd__mux4_1 _2793_ (.A0(\cordic_inst.cordic_inst.y[15] ),
    .A1(\cordic_inst.cordic_inst.y[16] ),
    .A2(\cordic_inst.cordic_inst.y[17] ),
    .A3(\cordic_inst.cordic_inst.y[18] ),
    .S0(net310),
    .S1(net299),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(_1095_),
    .A1(_1096_),
    .S(net290),
    .X(_1097_));
 sky130_fd_sc_hd__mux4_1 _2795_ (.A0(\cordic_inst.cordic_inst.y[31] ),
    .A1(_1091_),
    .A2(_1094_),
    .A3(_1097_),
    .S0(net240),
    .S1(net243),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(_1093_),
    .A1(_1096_),
    .S(net235),
    .X(_1099_));
 sky130_fd_sc_hd__mux4_1 _2797_ (.A0(\cordic_inst.cordic_inst.y[7] ),
    .A1(\cordic_inst.cordic_inst.y[8] ),
    .A2(\cordic_inst.cordic_inst.y[9] ),
    .A3(\cordic_inst.cordic_inst.y[10] ),
    .S0(net308),
    .S1(net297),
    .X(_1100_));
 sky130_fd_sc_hd__a221o_1 _2798_ (.A1(net218),
    .A2(_1095_),
    .B1(_1100_),
    .B2(net221),
    .C1(net277),
    .X(_1101_));
 sky130_fd_sc_hd__a21oi_1 _2799_ (.A1(net283),
    .A2(_1099_),
    .B1(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__a21o_1 _2800_ (.A1(net275),
    .A2(_1089_),
    .B1(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__mux4_1 _2801_ (.A0(\cordic_inst.cordic_inst.y[14] ),
    .A1(\cordic_inst.cordic_inst.y[15] ),
    .A2(\cordic_inst.cordic_inst.y[16] ),
    .A3(\cordic_inst.cordic_inst.y[17] ),
    .S0(net310),
    .S1(net299),
    .X(_1104_));
 sky130_fd_sc_hd__mux4_1 _2802_ (.A0(\cordic_inst.cordic_inst.y[18] ),
    .A1(\cordic_inst.cordic_inst.y[19] ),
    .A2(\cordic_inst.cordic_inst.y[20] ),
    .A3(\cordic_inst.cordic_inst.y[21] ),
    .S0(net311),
    .S1(net300),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(_1104_),
    .A1(_1105_),
    .S(net290),
    .X(_1106_));
 sky130_fd_sc_hd__mux4_1 _2804_ (.A0(\cordic_inst.cordic_inst.y[10] ),
    .A1(\cordic_inst.cordic_inst.y[11] ),
    .A2(\cordic_inst.cordic_inst.y[12] ),
    .A3(\cordic_inst.cordic_inst.y[13] ),
    .S0(net308),
    .S1(net297),
    .X(_1107_));
 sky130_fd_sc_hd__mux4_1 _2805_ (.A0(\cordic_inst.cordic_inst.y[6] ),
    .A1(\cordic_inst.cordic_inst.y[7] ),
    .A2(\cordic_inst.cordic_inst.y[8] ),
    .A3(\cordic_inst.cordic_inst.y[9] ),
    .S0(net308),
    .S1(net297),
    .X(_1108_));
 sky130_fd_sc_hd__a221o_1 _2806_ (.A1(net218),
    .A2(_1107_),
    .B1(_1108_),
    .B2(net221),
    .C1(net277),
    .X(_1109_));
 sky130_fd_sc_hd__a21o_1 _2807_ (.A1(net283),
    .A2(_1106_),
    .B1(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__mux4_1 _2808_ (.A0(\cordic_inst.cordic_inst.y[22] ),
    .A1(\cordic_inst.cordic_inst.y[23] ),
    .A2(\cordic_inst.cordic_inst.y[24] ),
    .A3(\cordic_inst.cordic_inst.y[25] ),
    .S0(net307),
    .S1(net301),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(\cordic_inst.cordic_inst.y[26] ),
    .A1(\cordic_inst.cordic_inst.y[27] ),
    .S(net306),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(_1078_),
    .A1(_1112_),
    .S(net232),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(_1111_),
    .A1(_1113_),
    .S(net291),
    .X(_1114_));
 sky130_fd_sc_hd__mux4_1 _2812_ (.A0(net262),
    .A1(_1074_),
    .A2(_1113_),
    .A3(_1111_),
    .S0(net234),
    .S1(net238),
    .X(_1115_));
 sky130_fd_sc_hd__o21ai_2 _2813_ (.A1(net243),
    .A2(_1115_),
    .B1(_1110_),
    .Y(_1116_));
 sky130_fd_sc_hd__mux4_1 _2814_ (.A0(\cordic_inst.cordic_inst.y[13] ),
    .A1(\cordic_inst.cordic_inst.y[14] ),
    .A2(\cordic_inst.cordic_inst.y[15] ),
    .A3(\cordic_inst.cordic_inst.y[16] ),
    .S0(net310),
    .S1(net299),
    .X(_1117_));
 sky130_fd_sc_hd__mux4_1 _2815_ (.A0(\cordic_inst.cordic_inst.y[17] ),
    .A1(\cordic_inst.cordic_inst.y[18] ),
    .A2(\cordic_inst.cordic_inst.y[19] ),
    .A3(\cordic_inst.cordic_inst.y[20] ),
    .S0(net311),
    .S1(net300),
    .X(_1118_));
 sky130_fd_sc_hd__mux2_1 _2816_ (.A0(_1117_),
    .A1(_1118_),
    .S(net290),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(\cordic_inst.cordic_inst.y[5] ),
    .A1(\cordic_inst.cordic_inst.y[6] ),
    .S(net308),
    .X(_1120_));
 sky130_fd_sc_hd__mux4_1 _2818_ (.A0(\cordic_inst.cordic_inst.y[5] ),
    .A1(\cordic_inst.cordic_inst.y[6] ),
    .A2(\cordic_inst.cordic_inst.y[7] ),
    .A3(\cordic_inst.cordic_inst.y[8] ),
    .S0(net308),
    .S1(net297),
    .X(_1121_));
 sky130_fd_sc_hd__mux4_2 _2819_ (.A0(\cordic_inst.cordic_inst.y[9] ),
    .A1(\cordic_inst.cordic_inst.y[10] ),
    .A2(\cordic_inst.cordic_inst.y[11] ),
    .A3(\cordic_inst.cordic_inst.y[12] ),
    .S0(net308),
    .S1(net297),
    .X(_1122_));
 sky130_fd_sc_hd__a221o_1 _2820_ (.A1(net221),
    .A2(_1121_),
    .B1(_1122_),
    .B2(net218),
    .C1(net275),
    .X(_1123_));
 sky130_fd_sc_hd__a21o_1 _2821_ (.A1(net283),
    .A2(_1119_),
    .B1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__mux4_1 _2822_ (.A0(\cordic_inst.cordic_inst.y[21] ),
    .A1(\cordic_inst.cordic_inst.y[22] ),
    .A2(\cordic_inst.cordic_inst.y[23] ),
    .A3(\cordic_inst.cordic_inst.y[24] ),
    .S0(net307),
    .S1(net301),
    .X(_1125_));
 sky130_fd_sc_hd__mux2_1 _2823_ (.A0(_1083_),
    .A1(_1085_),
    .S(net295),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(_1125_),
    .A1(_1126_),
    .S(net291),
    .X(_1127_));
 sky130_fd_sc_hd__a21o_1 _2825_ (.A1(net232),
    .A2(_1086_),
    .B1(_1072_),
    .X(_1128_));
 sky130_fd_sc_hd__a21o_1 _2826_ (.A1(net237),
    .A2(_1128_),
    .B1(_1071_),
    .X(_1129_));
 sky130_fd_sc_hd__mux4_2 _2827_ (.A0(net262),
    .A1(_1126_),
    .A2(_1128_),
    .A3(_1125_),
    .S0(net239),
    .S1(net233),
    .X(_1130_));
 sky130_fd_sc_hd__o21ai_2 _2828_ (.A1(net243),
    .A2(_1130_),
    .B1(_1124_),
    .Y(_1131_));
 sky130_fd_sc_hd__mux4_2 _2829_ (.A0(\cordic_inst.cordic_inst.y[16] ),
    .A1(\cordic_inst.cordic_inst.y[17] ),
    .A2(\cordic_inst.cordic_inst.y[18] ),
    .A3(\cordic_inst.cordic_inst.y[19] ),
    .S0(net310),
    .S1(net299),
    .X(_1132_));
 sky130_fd_sc_hd__mux4_1 _2830_ (.A0(\cordic_inst.cordic_inst.y[20] ),
    .A1(\cordic_inst.cordic_inst.y[21] ),
    .A2(\cordic_inst.cordic_inst.y[22] ),
    .A3(\cordic_inst.cordic_inst.y[23] ),
    .S0(net307),
    .S1(net301),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _2831_ (.A0(_1132_),
    .A1(_1133_),
    .S(net291),
    .X(_1134_));
 sky130_fd_sc_hd__mux4_1 _2832_ (.A0(\cordic_inst.cordic_inst.y[24] ),
    .A1(\cordic_inst.cordic_inst.y[25] ),
    .A2(\cordic_inst.cordic_inst.y[26] ),
    .A3(\cordic_inst.cordic_inst.y[27] ),
    .S0(net304),
    .S1(net295),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _2833_ (.A0(_1079_),
    .A1(_1135_),
    .S(net233),
    .X(_1136_));
 sky130_fd_sc_hd__mux4_2 _2834_ (.A0(_1079_),
    .A1(_1133_),
    .A2(_1135_),
    .A3(_1132_),
    .S0(net239),
    .S1(net233),
    .X(_1137_));
 sky130_fd_sc_hd__or2_1 _2835_ (.A(net242),
    .B(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__mux4_2 _2836_ (.A0(\cordic_inst.cordic_inst.y[8] ),
    .A1(\cordic_inst.cordic_inst.y[9] ),
    .A2(\cordic_inst.cordic_inst.y[10] ),
    .A3(\cordic_inst.cordic_inst.y[11] ),
    .S0(net308),
    .S1(net297),
    .X(_1139_));
 sky130_fd_sc_hd__mux4_2 _2837_ (.A0(\cordic_inst.cordic_inst.y[12] ),
    .A1(\cordic_inst.cordic_inst.y[13] ),
    .A2(\cordic_inst.cordic_inst.y[14] ),
    .A3(\cordic_inst.cordic_inst.y[15] ),
    .S0(net310),
    .S1(net299),
    .X(_1140_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(_1139_),
    .A1(_1140_),
    .S(net291),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(\cordic_inst.cordic_inst.y[4] ),
    .A1(\cordic_inst.cordic_inst.y[5] ),
    .S(net308),
    .X(_1142_));
 sky130_fd_sc_hd__mux4_2 _2840_ (.A0(\cordic_inst.cordic_inst.y[4] ),
    .A1(\cordic_inst.cordic_inst.y[5] ),
    .A2(\cordic_inst.cordic_inst.y[6] ),
    .A3(\cordic_inst.cordic_inst.y[7] ),
    .S0(net308),
    .S1(net297),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(\cordic_inst.cordic_inst.y[2] ),
    .A1(\cordic_inst.cordic_inst.y[3] ),
    .S(net311),
    .X(_1144_));
 sky130_fd_sc_hd__a221o_1 _2842_ (.A1(\cordic_inst.cordic_inst.y[1] ),
    .A2(net217),
    .B1(_0709_),
    .B2(_1144_),
    .C1(net275),
    .X(_1145_));
 sky130_fd_sc_hd__a32o_1 _2843_ (.A1(\cordic_inst.cordic_inst.y[0] ),
    .A2(net221),
    .A3(_0711_),
    .B1(_1143_),
    .B2(net219),
    .X(_1146_));
 sky130_fd_sc_hd__a211o_1 _2844_ (.A1(net286),
    .A2(_1141_),
    .B1(_1145_),
    .C1(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__and2_1 _2845_ (.A(_1138_),
    .B(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(_1118_),
    .A1(_1125_),
    .S(net290),
    .X(_1149_));
 sky130_fd_sc_hd__mux4_2 _2847_ (.A0(net262),
    .A1(_1085_),
    .A2(_1086_),
    .A3(_1083_),
    .S0(net233),
    .S1(net232),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(_1149_),
    .A1(_1150_),
    .S(net283),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(_1117_),
    .A1(_1122_),
    .S(net235),
    .X(_1152_));
 sky130_fd_sc_hd__and2_1 _2850_ (.A(net283),
    .B(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\cordic_inst.cordic_inst.y[3] ),
    .A1(\cordic_inst.cordic_inst.y[4] ),
    .S(net311),
    .X(_1154_));
 sky130_fd_sc_hd__a221o_1 _2852_ (.A1(\cordic_inst.cordic_inst.y[2] ),
    .A2(net217),
    .B1(net216),
    .B2(_1154_),
    .C1(net275),
    .X(_1155_));
 sky130_fd_sc_hd__a32o_1 _2853_ (.A1(\cordic_inst.cordic_inst.y[1] ),
    .A2(net221),
    .A3(_0711_),
    .B1(_1121_),
    .B2(net218),
    .X(_1156_));
 sky130_fd_sc_hd__o32a_1 _2854_ (.A1(_1153_),
    .A2(_1155_),
    .A3(_1156_),
    .B1(_1151_),
    .B2(net243),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(_1104_),
    .A1(_1107_),
    .S(net235),
    .X(_1158_));
 sky130_fd_sc_hd__a221o_1 _2856_ (.A1(net216),
    .A2(_1142_),
    .B1(_1144_),
    .B2(_0713_),
    .C1(net275),
    .X(_1159_));
 sky130_fd_sc_hd__a22o_1 _2857_ (.A1(net218),
    .A2(_1108_),
    .B1(_1158_),
    .B2(net283),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_1 _2858_ (.A0(_1105_),
    .A1(_1111_),
    .S(net290),
    .X(_1161_));
 sky130_fd_sc_hd__mux4_2 _2859_ (.A0(net263),
    .A1(_1073_),
    .A2(_1078_),
    .A3(_1112_),
    .S0(net232),
    .S1(net237),
    .X(_1162_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(_1161_),
    .A1(_1162_),
    .S(net283),
    .X(_1163_));
 sky130_fd_sc_hd__o22a_1 _2861_ (.A1(_1159_),
    .A2(_1160_),
    .B1(_1163_),
    .B2(net243),
    .X(_1164_));
 sky130_fd_sc_hd__a221o_1 _2862_ (.A1(net216),
    .A2(_1120_),
    .B1(_1154_),
    .B2(_0713_),
    .C1(net276),
    .X(_1165_));
 sky130_fd_sc_hd__a22o_1 _2863_ (.A1(net283),
    .A2(_1097_),
    .B1(_1100_),
    .B2(net218),
    .X(_1166_));
 sky130_fd_sc_hd__a211o_1 _2864_ (.A1(net233),
    .A2(_1087_),
    .B1(_1071_),
    .C1(net238),
    .X(_1167_));
 sky130_fd_sc_hd__o21ai_1 _2865_ (.A1(net285),
    .A2(_1094_),
    .B1(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__a2bb2o_1 _2866_ (.A1_N(_1165_),
    .A2_N(_1166_),
    .B1(_1168_),
    .B2(net275),
    .X(_1169_));
 sky130_fd_sc_hd__or4b_1 _2867_ (.A(_1148_),
    .B(_1157_),
    .C(_1164_),
    .D_N(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(_1132_),
    .A1(_1140_),
    .S(net234),
    .X(_1171_));
 sky130_fd_sc_hd__a22o_1 _2869_ (.A1(net219),
    .A2(_1139_),
    .B1(_1143_),
    .B2(net221),
    .X(_1172_));
 sky130_fd_sc_hd__a21oi_1 _2870_ (.A1(net286),
    .A2(_1171_),
    .B1(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(_1133_),
    .A1(_1135_),
    .S(net291),
    .X(_1174_));
 sky130_fd_sc_hd__a211o_1 _2872_ (.A1(net233),
    .A2(_1079_),
    .B1(_1071_),
    .C1(net238),
    .X(_1175_));
 sky130_fd_sc_hd__o21ai_1 _2873_ (.A1(net286),
    .A2(_1174_),
    .B1(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(_1173_),
    .A1(_1176_),
    .S(net275),
    .X(_1177_));
 sky130_fd_sc_hd__and2b_1 _2875_ (.A_N(_1170_),
    .B(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__nand4_1 _2876_ (.A(_1103_),
    .B(_1116_),
    .C(_1131_),
    .D(_1177_),
    .Y(_1179_));
 sky130_fd_sc_hd__or2_1 _2877_ (.A(_1170_),
    .B(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__nand2_1 _2878_ (.A(net241),
    .B(_1150_),
    .Y(_1181_));
 sky130_fd_sc_hd__mux4_1 _2879_ (.A0(net262),
    .A1(_1149_),
    .A2(_1150_),
    .A3(_1152_),
    .S0(net243),
    .S1(net240),
    .X(_1182_));
 sky130_fd_sc_hd__a21bo_1 _2880_ (.A1(net239),
    .A2(_1136_),
    .B1_N(_1070_),
    .X(_1183_));
 sky130_fd_sc_hd__mux4_2 _2881_ (.A0(net262),
    .A1(_1134_),
    .A2(_1136_),
    .A3(_1141_),
    .S0(net242),
    .S1(net239),
    .X(_1184_));
 sky130_fd_sc_hd__or2_1 _2882_ (.A(_1182_),
    .B(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__a21bo_1 _2883_ (.A1(net241),
    .A2(_1162_),
    .B1_N(_1070_),
    .X(_1186_));
 sky130_fd_sc_hd__mux4_1 _2884_ (.A0(net262),
    .A1(_1161_),
    .A2(_1162_),
    .A3(_1158_),
    .S0(net243),
    .S1(net240),
    .X(_1187_));
 sky130_fd_sc_hd__or3_1 _2885_ (.A(_1098_),
    .B(_1185_),
    .C(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__or2_1 _2886_ (.A(_1180_),
    .B(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__mux4_2 _2887_ (.A0(net262),
    .A1(_1080_),
    .A2(_1174_),
    .A3(_1171_),
    .S0(net238),
    .S1(net242),
    .X(_1190_));
 sky130_fd_sc_hd__a21boi_1 _2888_ (.A1(net241),
    .A2(_1129_),
    .B1_N(_1070_),
    .Y(_1191_));
 sky130_fd_sc_hd__mux4_2 _2889_ (.A0(net262),
    .A1(_1127_),
    .A2(_1129_),
    .A3(_1119_),
    .S0(net242),
    .S1(net239),
    .X(_1192_));
 sky130_fd_sc_hd__mux4_2 _2890_ (.A0(net262),
    .A1(_1075_),
    .A2(_1114_),
    .A3(_1106_),
    .S0(net238),
    .S1(net243),
    .X(_1193_));
 sky130_fd_sc_hd__or3_1 _2891_ (.A(_1190_),
    .B(_1192_),
    .C(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__or4_2 _2892_ (.A(_1170_),
    .B(_1179_),
    .C(_1188_),
    .D(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__or2_1 _2893_ (.A(net285),
    .B(_1099_),
    .X(_1196_));
 sky130_fd_sc_hd__or2_1 _2894_ (.A(net238),
    .B(_1088_),
    .X(_1197_));
 sky130_fd_sc_hd__a31o_1 _2895_ (.A1(net244),
    .A2(_1196_),
    .A3(_1197_),
    .B1(net215),
    .X(_1198_));
 sky130_fd_sc_hd__nand2_1 _2896_ (.A(net244),
    .B(_1151_),
    .Y(_1199_));
 sky130_fd_sc_hd__nand2_1 _2897_ (.A(_1069_),
    .B(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__a21oi_4 _2898_ (.A1(net246),
    .A2(_1137_),
    .B1(net215),
    .Y(_1201_));
 sky130_fd_sc_hd__nand2_1 _2899_ (.A(_1199_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__o21ai_2 _2900_ (.A1(net276),
    .A2(_1168_),
    .B1(_1069_),
    .Y(_1203_));
 sky130_fd_sc_hd__a21o_1 _2901_ (.A1(net244),
    .A2(_1163_),
    .B1(net215),
    .X(_1204_));
 sky130_fd_sc_hd__a211o_1 _2902_ (.A1(net244),
    .A2(_1163_),
    .B1(_1202_),
    .C1(_1203_),
    .X(_1205_));
 sky130_fd_sc_hd__nand2_1 _2903_ (.A(net246),
    .B(_1130_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand2_1 _2904_ (.A(_1069_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__o21a_1 _2905_ (.A1(net276),
    .A2(_1176_),
    .B1(_1069_),
    .X(_1208_));
 sky130_fd_sc_hd__nand2_1 _2906_ (.A(_1206_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__a21o_1 _2907_ (.A1(net246),
    .A2(_1115_),
    .B1(_1068_),
    .X(_1210_));
 sky130_fd_sc_hd__a21o_1 _2908_ (.A1(net242),
    .A2(_1183_),
    .B1(net215),
    .X(_1211_));
 sky130_fd_sc_hd__a21oi_1 _2909_ (.A1(_1070_),
    .A2(_1181_),
    .B1(net274),
    .Y(_1212_));
 sky130_fd_sc_hd__a21o_1 _2910_ (.A1(net242),
    .A2(_1186_),
    .B1(net215),
    .X(_1213_));
 sky130_fd_sc_hd__a21oi_1 _2911_ (.A1(_1070_),
    .A2(_1092_),
    .B1(net274),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _2912_ (.A(net272),
    .B(_1189_),
    .Y(_1215_));
 sky130_fd_sc_hd__and2_1 _2913_ (.A(net271),
    .B(_1195_),
    .X(_1216_));
 sky130_fd_sc_hd__o21a_1 _2914_ (.A1(_1195_),
    .A2(_1198_),
    .B1(net271),
    .X(_1217_));
 sky130_fd_sc_hd__o31a_1 _2915_ (.A1(_1195_),
    .A2(_1198_),
    .A3(_1205_),
    .B1(net270),
    .X(_1218_));
 sky130_fd_sc_hd__a21o_1 _2916_ (.A1(net270),
    .A2(_1209_),
    .B1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__a21o_1 _2917_ (.A1(net270),
    .A2(_1210_),
    .B1(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__a21o_1 _2918_ (.A1(net270),
    .A2(_1090_),
    .B1(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__a21o_1 _2919_ (.A1(net269),
    .A2(_1211_),
    .B1(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__a21o_1 _2920_ (.A1(net269),
    .A2(_1212_),
    .B1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__a21o_1 _2921_ (.A1(net269),
    .A2(_1213_),
    .B1(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__a21o_1 _2922_ (.A1(net269),
    .A2(_1214_),
    .B1(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__o21a_1 _2923_ (.A1(_1082_),
    .A2(_1225_),
    .B1(net269),
    .X(_1226_));
 sky130_fd_sc_hd__nor2_1 _2924_ (.A(net274),
    .B(_1191_),
    .Y(_1227_));
 sky130_fd_sc_hd__a21oi_1 _2925_ (.A1(net269),
    .A2(_1227_),
    .B1(_1226_),
    .Y(_1228_));
 sky130_fd_sc_hd__xnor2_1 _2926_ (.A(_1077_),
    .B(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__and2b_1 _2927_ (.A_N(_1229_),
    .B(\cordic_inst.cordic_inst.x[30] ),
    .X(_1230_));
 sky130_fd_sc_hd__xor2_1 _2928_ (.A(\cordic_inst.cordic_inst.x[30] ),
    .B(_1229_),
    .X(_1231_));
 sky130_fd_sc_hd__or2_1 _2929_ (.A(net215),
    .B(_1227_),
    .X(_1232_));
 sky130_fd_sc_hd__xnor2_1 _2930_ (.A(_1226_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__nor2_1 _2931_ (.A(\cordic_inst.cordic_inst.x[29] ),
    .B(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__xnor2_1 _2932_ (.A(_1082_),
    .B(_1225_),
    .Y(_1235_));
 sky130_fd_sc_hd__nand2_1 _2933_ (.A(\cordic_inst.cordic_inst.x[28] ),
    .B(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__and2_1 _2934_ (.A(\cordic_inst.cordic_inst.x[29] ),
    .B(_1233_),
    .X(_1237_));
 sky130_fd_sc_hd__nand2_1 _2935_ (.A(\cordic_inst.cordic_inst.x[29] ),
    .B(_1233_),
    .Y(_1238_));
 sky130_fd_sc_hd__or2_1 _2936_ (.A(\cordic_inst.cordic_inst.x[28] ),
    .B(_1235_),
    .X(_1239_));
 sky130_fd_sc_hd__and2_1 _2937_ (.A(_1236_),
    .B(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__a31o_1 _2938_ (.A1(_1116_),
    .A2(_1131_),
    .A3(_1178_),
    .B1(net251),
    .X(_1241_));
 sky130_fd_sc_hd__xnor2_1 _2939_ (.A(_1103_),
    .B(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__nor2_1 _2940_ (.A(\cordic_inst.cordic_inst.x[7] ),
    .B(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__nand2_1 _2941_ (.A(\cordic_inst.cordic_inst.x[7] ),
    .B(_1242_),
    .Y(_1244_));
 sky130_fd_sc_hd__a21o_1 _2942_ (.A1(_1131_),
    .A2(_1178_),
    .B1(net251),
    .X(_1245_));
 sky130_fd_sc_hd__xor2_1 _2943_ (.A(_1116_),
    .B(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__nand2b_2 _2944_ (.A_N(_1246_),
    .B(\cordic_inst.cordic_inst.x[6] ),
    .Y(_1247_));
 sky130_fd_sc_hd__nand2b_1 _2945_ (.A_N(\cordic_inst.cordic_inst.x[6] ),
    .B(_1246_),
    .Y(_1248_));
 sky130_fd_sc_hd__nand2_1 _2946_ (.A(_1247_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__or2_1 _2947_ (.A(net251),
    .B(_1178_),
    .X(_1250_));
 sky130_fd_sc_hd__xor2_1 _2948_ (.A(_1131_),
    .B(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__and2_1 _2949_ (.A(_0602_),
    .B(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__nor2_1 _2950_ (.A(_0602_),
    .B(_1251_),
    .Y(_1253_));
 sky130_fd_sc_hd__inv_2 _2951_ (.A(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _2952_ (.A(net270),
    .B(_1170_),
    .Y(_1255_));
 sky130_fd_sc_hd__xnor2_1 _2953_ (.A(_1177_),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__and2_1 _2954_ (.A(\cordic_inst.cordic_inst.x[4] ),
    .B(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__inv_2 _2955_ (.A(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__nor2_1 _2956_ (.A(\cordic_inst.cordic_inst.x[4] ),
    .B(_1256_),
    .Y(_1259_));
 sky130_fd_sc_hd__or2_1 _2957_ (.A(_1257_),
    .B(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__o31a_1 _2958_ (.A1(_1148_),
    .A2(_1157_),
    .A3(_1164_),
    .B1(net270),
    .X(_1261_));
 sky130_fd_sc_hd__xor2_1 _2959_ (.A(_1169_),
    .B(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__nand2_1 _2960_ (.A(\cordic_inst.cordic_inst.x[3] ),
    .B(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__o21a_1 _2961_ (.A1(_1148_),
    .A2(_1157_),
    .B1(net270),
    .X(_1264_));
 sky130_fd_sc_hd__xnor2_1 _2962_ (.A(_1164_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__nand2_1 _2963_ (.A(\cordic_inst.cordic_inst.x[2] ),
    .B(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__and3_1 _2964_ (.A(net270),
    .B(_1138_),
    .C(_1147_),
    .X(_1267_));
 sky130_fd_sc_hd__xnor2_1 _2965_ (.A(_1157_),
    .B(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__nand2_1 _2966_ (.A(\cordic_inst.cordic_inst.x[1] ),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__and3_1 _2967_ (.A(_0603_),
    .B(_1138_),
    .C(_1147_),
    .X(_1270_));
 sky130_fd_sc_hd__xor2_1 _2968_ (.A(\cordic_inst.cordic_inst.x[1] ),
    .B(_1268_),
    .X(_1271_));
 sky130_fd_sc_hd__nand2b_1 _2969_ (.A_N(_1270_),
    .B(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__xnor2_1 _2970_ (.A(\cordic_inst.cordic_inst.x[2] ),
    .B(_1265_),
    .Y(_1273_));
 sky130_fd_sc_hd__a21o_1 _2971_ (.A1(_1269_),
    .A2(_1272_),
    .B1(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__or2_1 _2972_ (.A(\cordic_inst.cordic_inst.x[3] ),
    .B(_1262_),
    .X(_1275_));
 sky130_fd_sc_hd__nand2_1 _2973_ (.A(_1263_),
    .B(_1275_),
    .Y(_1276_));
 sky130_fd_sc_hd__a21o_1 _2974_ (.A1(_1266_),
    .A2(_1274_),
    .B1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__a21o_1 _2975_ (.A1(_1263_),
    .A2(_1277_),
    .B1(_1260_),
    .X(_1278_));
 sky130_fd_sc_hd__nand2_1 _2976_ (.A(_1258_),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__or2_1 _2977_ (.A(_1252_),
    .B(_1253_),
    .X(_1280_));
 sky130_fd_sc_hd__a31o_1 _2978_ (.A1(_1254_),
    .A2(_1258_),
    .A3(_1278_),
    .B1(_1252_),
    .X(_1281_));
 sky130_fd_sc_hd__a311o_2 _2979_ (.A1(_1254_),
    .A2(_1258_),
    .A3(_1278_),
    .B1(_1252_),
    .C1(_1249_),
    .X(_1282_));
 sky130_fd_sc_hd__nand2b_1 _2980_ (.A_N(_1243_),
    .B(_1244_),
    .Y(_1283_));
 sky130_fd_sc_hd__a31o_1 _2981_ (.A1(_1244_),
    .A2(_1247_),
    .A3(_1282_),
    .B1(_1243_),
    .X(_1284_));
 sky130_fd_sc_hd__nand2_1 _2982_ (.A(net272),
    .B(_1180_),
    .Y(_1285_));
 sky130_fd_sc_hd__xor2_1 _2983_ (.A(_1184_),
    .B(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__nand2_1 _2984_ (.A(\cordic_inst.cordic_inst.x[8] ),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__or2_1 _2985_ (.A(\cordic_inst.cordic_inst.x[8] ),
    .B(_1286_),
    .X(_1288_));
 sky130_fd_sc_hd__nand2_1 _2986_ (.A(_1287_),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__a311o_1 _2987_ (.A1(_1244_),
    .A2(_1247_),
    .A3(_1282_),
    .B1(_1289_),
    .C1(_1243_),
    .X(_1290_));
 sky130_fd_sc_hd__o21ai_1 _2988_ (.A1(_1180_),
    .A2(_1184_),
    .B1(net272),
    .Y(_1291_));
 sky130_fd_sc_hd__xnor2_1 _2989_ (.A(_1182_),
    .B(_1291_),
    .Y(_1292_));
 sky130_fd_sc_hd__and2b_1 _2990_ (.A_N(\cordic_inst.cordic_inst.x[9] ),
    .B(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__nand2b_1 _2991_ (.A_N(_1292_),
    .B(\cordic_inst.cordic_inst.x[9] ),
    .Y(_1294_));
 sky130_fd_sc_hd__nand2b_1 _2992_ (.A_N(_1293_),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__xnor2_1 _2993_ (.A(_1198_),
    .B(_1216_),
    .Y(_1296_));
 sky130_fd_sc_hd__nor2_1 _2994_ (.A(\cordic_inst.cordic_inst.x[15] ),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__nand2_1 _2995_ (.A(\cordic_inst.cordic_inst.x[15] ),
    .B(_1296_),
    .Y(_1298_));
 sky130_fd_sc_hd__and2b_1 _2996_ (.A_N(_1297_),
    .B(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__o31a_1 _2997_ (.A1(_1189_),
    .A2(_1190_),
    .A3(_1192_),
    .B1(net272),
    .X(_1300_));
 sky130_fd_sc_hd__xnor2_1 _2998_ (.A(_1193_),
    .B(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__nand2_1 _2999_ (.A(\cordic_inst.cordic_inst.x[14] ),
    .B(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__xor2_1 _3000_ (.A(\cordic_inst.cordic_inst.x[14] ),
    .B(_1301_),
    .X(_1303_));
 sky130_fd_sc_hd__and2_1 _3001_ (.A(_1299_),
    .B(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__o21a_1 _3002_ (.A1(_1189_),
    .A2(_1190_),
    .B1(net272),
    .X(_1305_));
 sky130_fd_sc_hd__xnor2_1 _3003_ (.A(_1192_),
    .B(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__or2_1 _3004_ (.A(\cordic_inst.cordic_inst.x[13] ),
    .B(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__nand2_1 _3005_ (.A(\cordic_inst.cordic_inst.x[13] ),
    .B(_1306_),
    .Y(_1308_));
 sky130_fd_sc_hd__and2_1 _3006_ (.A(_1307_),
    .B(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__xor2_2 _3007_ (.A(_1190_),
    .B(_1215_),
    .X(_1310_));
 sky130_fd_sc_hd__xnor2_1 _3008_ (.A(\cordic_inst.cordic_inst.x[12] ),
    .B(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__inv_2 _3009_ (.A(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__and3_1 _3010_ (.A(_1304_),
    .B(_1309_),
    .C(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__o31a_1 _3011_ (.A1(_1180_),
    .A2(_1185_),
    .A3(_1187_),
    .B1(net272),
    .X(_1314_));
 sky130_fd_sc_hd__xnor2_1 _3012_ (.A(_1098_),
    .B(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__nor2_1 _3013_ (.A(\cordic_inst.cordic_inst.x[11] ),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2_1 _3014_ (.A(\cordic_inst.cordic_inst.x[11] ),
    .B(_1315_),
    .Y(_1317_));
 sky130_fd_sc_hd__nand2b_1 _3015_ (.A_N(_1316_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__o21ai_1 _3016_ (.A1(_1180_),
    .A2(_1185_),
    .B1(net272),
    .Y(_1319_));
 sky130_fd_sc_hd__xor2_1 _3017_ (.A(_1187_),
    .B(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__nand2_1 _3018_ (.A(\cordic_inst.cordic_inst.x[10] ),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__or2_1 _3019_ (.A(\cordic_inst.cordic_inst.x[10] ),
    .B(_1320_),
    .X(_1322_));
 sky130_fd_sc_hd__nand2_1 _3020_ (.A(_1321_),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__nor2_1 _3021_ (.A(_1318_),
    .B(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__or4bb_1 _3022_ (.A(_1290_),
    .B(_1295_),
    .C_N(_1313_),
    .D_N(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__a22o_1 _3023_ (.A1(\cordic_inst.cordic_inst.x[13] ),
    .A2(_1306_),
    .B1(_1310_),
    .B2(\cordic_inst.cordic_inst.x[12] ),
    .X(_1326_));
 sky130_fd_sc_hd__a21oi_1 _3024_ (.A1(_1298_),
    .A2(_1302_),
    .B1(_1297_),
    .Y(_1327_));
 sky130_fd_sc_hd__a31o_1 _3025_ (.A1(_1304_),
    .A2(_1307_),
    .A3(_1326_),
    .B1(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__a21o_1 _3026_ (.A1(_1317_),
    .A2(_1321_),
    .B1(_1316_),
    .X(_1329_));
 sky130_fd_sc_hd__a2111o_1 _3027_ (.A1(_1287_),
    .A2(_1294_),
    .B1(_1318_),
    .C1(_1323_),
    .D1(_1293_),
    .X(_1330_));
 sky130_fd_sc_hd__a21bo_1 _3028_ (.A1(_1329_),
    .A2(_1330_),
    .B1_N(_1313_),
    .X(_1331_));
 sky130_fd_sc_hd__nand3b_2 _3029_ (.A_N(_1328_),
    .B(_1331_),
    .C(_1325_),
    .Y(_1332_));
 sky130_fd_sc_hd__or2_1 _3030_ (.A(_1068_),
    .B(_1090_),
    .X(_1333_));
 sky130_fd_sc_hd__xnor2_1 _3031_ (.A(_1220_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__xnor2_1 _3032_ (.A(\cordic_inst.cordic_inst.x[23] ),
    .B(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__xnor2_1 _3033_ (.A(_1210_),
    .B(_1219_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand2_1 _3034_ (.A(\cordic_inst.cordic_inst.x[22] ),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__or2_1 _3035_ (.A(\cordic_inst.cordic_inst.x[22] ),
    .B(_1336_),
    .X(_1338_));
 sky130_fd_sc_hd__nand2_1 _3036_ (.A(_1337_),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__xor2_1 _3037_ (.A(_1208_),
    .B(_1218_),
    .X(_1340_));
 sky130_fd_sc_hd__nand2_1 _3038_ (.A(\cordic_inst.cordic_inst.x[20] ),
    .B(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__or2_1 _3039_ (.A(\cordic_inst.cordic_inst.x[20] ),
    .B(_1340_),
    .X(_1342_));
 sky130_fd_sc_hd__nand2_1 _3040_ (.A(_1341_),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__o21bai_1 _3041_ (.A1(net251),
    .A2(_1208_),
    .B1_N(_1218_),
    .Y(_1344_));
 sky130_fd_sc_hd__xnor2_1 _3042_ (.A(_1207_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__nor2_1 _3043_ (.A(\cordic_inst.cordic_inst.x[21] ),
    .B(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__nand2_1 _3044_ (.A(\cordic_inst.cordic_inst.x[21] ),
    .B(_1345_),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2b_1 _3045_ (.A_N(_1346_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__or4_1 _3046_ (.A(_1335_),
    .B(_1339_),
    .C(_1343_),
    .D(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__a21oi_1 _3047_ (.A1(net273),
    .A2(_1202_),
    .B1(_1217_),
    .Y(_1350_));
 sky130_fd_sc_hd__o41a_1 _3048_ (.A1(_1195_),
    .A2(_1198_),
    .A3(_1202_),
    .A4(_1204_),
    .B1(net273),
    .X(_1351_));
 sky130_fd_sc_hd__xnor2_1 _3049_ (.A(_1203_),
    .B(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__nor2_1 _3050_ (.A(\cordic_inst.cordic_inst.x[19] ),
    .B(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand2_1 _3051_ (.A(\cordic_inst.cordic_inst.x[19] ),
    .B(_1352_),
    .Y(_1354_));
 sky130_fd_sc_hd__nand2b_1 _3052_ (.A_N(_1353_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__xor2_1 _3053_ (.A(_1204_),
    .B(_1350_),
    .X(_1356_));
 sky130_fd_sc_hd__nand2_1 _3054_ (.A(\cordic_inst.cordic_inst.x[18] ),
    .B(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__xnor2_1 _3055_ (.A(\cordic_inst.cordic_inst.x[18] ),
    .B(_1356_),
    .Y(_1358_));
 sky130_fd_sc_hd__or2_1 _3056_ (.A(_1355_),
    .B(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__xor2_2 _3057_ (.A(_1201_),
    .B(_1217_),
    .X(_1360_));
 sky130_fd_sc_hd__xor2_1 _3058_ (.A(\cordic_inst.cordic_inst.x[16] ),
    .B(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__xnor2_1 _3059_ (.A(\cordic_inst.cordic_inst.x[16] ),
    .B(_1360_),
    .Y(_1362_));
 sky130_fd_sc_hd__o21bai_1 _3060_ (.A1(net250),
    .A2(_1201_),
    .B1_N(_1217_),
    .Y(_1363_));
 sky130_fd_sc_hd__xnor2_1 _3061_ (.A(_1200_),
    .B(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__nor2_1 _3062_ (.A(\cordic_inst.cordic_inst.x[17] ),
    .B(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__and2_1 _3063_ (.A(\cordic_inst.cordic_inst.x[17] ),
    .B(_1364_),
    .X(_1366_));
 sky130_fd_sc_hd__or2_1 _3064_ (.A(_1365_),
    .B(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__nor4_1 _3065_ (.A(_1349_),
    .B(_1359_),
    .C(_1362_),
    .D(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__and2_1 _3066_ (.A(_1341_),
    .B(_1347_),
    .X(_1369_));
 sky130_fd_sc_hd__or4_1 _3067_ (.A(_1335_),
    .B(_1339_),
    .C(_1346_),
    .D(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__o21ba_1 _3068_ (.A1(\cordic_inst.cordic_inst.x[23] ),
    .A2(_1334_),
    .B1_N(_1337_),
    .X(_1371_));
 sky130_fd_sc_hd__a21oi_1 _3069_ (.A1(\cordic_inst.cordic_inst.x[23] ),
    .A2(_1334_),
    .B1(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__a22oi_1 _3070_ (.A1(\cordic_inst.cordic_inst.x[16] ),
    .A2(_1360_),
    .B1(_1364_),
    .B2(\cordic_inst.cordic_inst.x[17] ),
    .Y(_1373_));
 sky130_fd_sc_hd__a21o_1 _3071_ (.A1(_1354_),
    .A2(_1357_),
    .B1(_1353_),
    .X(_1374_));
 sky130_fd_sc_hd__o31a_1 _3072_ (.A1(_1359_),
    .A2(_1365_),
    .A3(_1373_),
    .B1(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__o211a_1 _3073_ (.A1(_1349_),
    .A2(_1375_),
    .B1(_1372_),
    .C1(_1370_),
    .X(_1376_));
 sky130_fd_sc_hd__a21bo_1 _3074_ (.A1(_1332_),
    .A2(_1368_),
    .B1_N(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__xnor2_1 _3075_ (.A(_1211_),
    .B(_1221_),
    .Y(_1378_));
 sky130_fd_sc_hd__and2_1 _3076_ (.A(\cordic_inst.cordic_inst.x[24] ),
    .B(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__nor2_1 _3077_ (.A(\cordic_inst.cordic_inst.x[24] ),
    .B(_1378_),
    .Y(_1380_));
 sky130_fd_sc_hd__nor2_1 _3078_ (.A(_1379_),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _3079_ (.A(_1377_),
    .B(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__or2_1 _3080_ (.A(net215),
    .B(_1214_),
    .X(_1383_));
 sky130_fd_sc_hd__xnor2_1 _3081_ (.A(_1224_),
    .B(_1383_),
    .Y(_1384_));
 sky130_fd_sc_hd__xor2_1 _3082_ (.A(\cordic_inst.cordic_inst.x[27] ),
    .B(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__xnor2_1 _3083_ (.A(_1213_),
    .B(_1223_),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_1 _3084_ (.A(\cordic_inst.cordic_inst.x[26] ),
    .B(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__or2_1 _3085_ (.A(\cordic_inst.cordic_inst.x[26] ),
    .B(_1386_),
    .X(_1388_));
 sky130_fd_sc_hd__and2_1 _3086_ (.A(_1387_),
    .B(_1388_),
    .X(_1389_));
 sky130_fd_sc_hd__inv_2 _3087_ (.A(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__or2_1 _3088_ (.A(net215),
    .B(_1212_),
    .X(_1391_));
 sky130_fd_sc_hd__xnor2_1 _3089_ (.A(_1222_),
    .B(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__and2_1 _3090_ (.A(\cordic_inst.cordic_inst.x[25] ),
    .B(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__nor2_1 _3091_ (.A(\cordic_inst.cordic_inst.x[25] ),
    .B(_1392_),
    .Y(_1394_));
 sky130_fd_sc_hd__nor2_1 _3092_ (.A(_1393_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__and4b_1 _3093_ (.A_N(_1382_),
    .B(_1385_),
    .C(_1389_),
    .D(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__nor2_1 _3094_ (.A(_1379_),
    .B(_1393_),
    .Y(_1397_));
 sky130_fd_sc_hd__and4bb_1 _3095_ (.A_N(_1394_),
    .B_N(_1397_),
    .C(_1385_),
    .D(_1389_),
    .X(_1398_));
 sky130_fd_sc_hd__o21ba_1 _3096_ (.A1(\cordic_inst.cordic_inst.x[27] ),
    .A2(_1384_),
    .B1_N(_1387_),
    .X(_1399_));
 sky130_fd_sc_hd__a21o_1 _3097_ (.A1(\cordic_inst.cordic_inst.x[27] ),
    .A2(_1384_),
    .B1(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__o31ai_4 _3098_ (.A1(_1396_),
    .A2(_1398_),
    .A3(_1400_),
    .B1(_1240_),
    .Y(_1401_));
 sky130_fd_sc_hd__a31o_1 _3099_ (.A1(_1236_),
    .A2(_1238_),
    .A3(_1401_),
    .B1(_1234_),
    .X(_1402_));
 sky130_fd_sc_hd__a311oi_1 _3100_ (.A1(_1236_),
    .A2(_1238_),
    .A3(_1401_),
    .B1(_1234_),
    .C1(_1231_),
    .Y(_1403_));
 sky130_fd_sc_hd__o31a_1 _3101_ (.A1(_1077_),
    .A2(_1226_),
    .A3(_1227_),
    .B1(net269),
    .X(_1404_));
 sky130_fd_sc_hd__xor2_1 _3102_ (.A(_1002_),
    .B(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__o21ai_1 _3103_ (.A1(_1230_),
    .A2(_1403_),
    .B1(_1405_),
    .Y(_1406_));
 sky130_fd_sc_hd__or3_1 _3104_ (.A(_1230_),
    .B(_1403_),
    .C(_1405_),
    .X(_1407_));
 sky130_fd_sc_hd__a32o_1 _3105_ (.A1(net179),
    .A2(_1406_),
    .A3(_1407_),
    .B1(net163),
    .B2(net265),
    .X(_0529_));
 sky130_fd_sc_hd__xor2_1 _3106_ (.A(_1231_),
    .B(_1402_),
    .X(_1408_));
 sky130_fd_sc_hd__a22o_1 _3107_ (.A1(\cordic_inst.cordic_inst.x[30] ),
    .A2(net163),
    .B1(_1408_),
    .B2(net179),
    .X(_0528_));
 sky130_fd_sc_hd__o211ai_1 _3108_ (.A1(_1234_),
    .A2(_1237_),
    .B1(_1401_),
    .C1(_1236_),
    .Y(_1409_));
 sky130_fd_sc_hd__a211o_1 _3109_ (.A1(_1236_),
    .A2(_1401_),
    .B1(_1237_),
    .C1(_1234_),
    .X(_1410_));
 sky130_fd_sc_hd__a32o_1 _3110_ (.A1(net179),
    .A2(_1409_),
    .A3(_1410_),
    .B1(net163),
    .B2(\cordic_inst.cordic_inst.x[29] ),
    .X(_0527_));
 sky130_fd_sc_hd__or4_1 _3111_ (.A(_1240_),
    .B(_1396_),
    .C(_1398_),
    .D(_1400_),
    .X(_1411_));
 sky130_fd_sc_hd__a32o_1 _3112_ (.A1(net181),
    .A2(_1401_),
    .A3(_1411_),
    .B1(net163),
    .B2(\cordic_inst.cordic_inst.x[28] ),
    .X(_0526_));
 sky130_fd_sc_hd__a21o_1 _3113_ (.A1(_1382_),
    .A2(_1397_),
    .B1(_1394_),
    .X(_1412_));
 sky130_fd_sc_hd__or2_1 _3114_ (.A(_1390_),
    .B(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__nand2_1 _3115_ (.A(_1387_),
    .B(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__xnor2_1 _3116_ (.A(_1385_),
    .B(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__o2bb2ai_1 _3117_ (.A1_N(\cordic_inst.cordic_inst.x[27] ),
    .A2_N(net163),
    .B1(_1415_),
    .B2(net176),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_1 _3118_ (.A(_1390_),
    .B(_1412_),
    .Y(_1416_));
 sky130_fd_sc_hd__a32o_1 _3119_ (.A1(net181),
    .A2(_1413_),
    .A3(_1416_),
    .B1(net163),
    .B2(\cordic_inst.cordic_inst.x[26] ),
    .X(_0524_));
 sky130_fd_sc_hd__a21oi_1 _3120_ (.A1(_1377_),
    .A2(_1381_),
    .B1(_1379_),
    .Y(_1417_));
 sky130_fd_sc_hd__xnor2_1 _3121_ (.A(_1395_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__a22o_1 _3122_ (.A1(\cordic_inst.cordic_inst.x[25] ),
    .A2(net163),
    .B1(_1418_),
    .B2(net181),
    .X(_0523_));
 sky130_fd_sc_hd__or2_1 _3123_ (.A(_1377_),
    .B(_1381_),
    .X(_1419_));
 sky130_fd_sc_hd__a32o_1 _3124_ (.A1(net181),
    .A2(_1382_),
    .A3(_1419_),
    .B1(net164),
    .B2(\cordic_inst.cordic_inst.x[24] ),
    .X(_0522_));
 sky130_fd_sc_hd__or4b_1 _3125_ (.A(_1359_),
    .B(_1362_),
    .C(_1367_),
    .D_N(_1332_),
    .X(_1420_));
 sky130_fd_sc_hd__a21o_1 _3126_ (.A1(_1375_),
    .A2(_1420_),
    .B1(_1343_),
    .X(_1421_));
 sky130_fd_sc_hd__a21o_1 _3127_ (.A1(_1369_),
    .A2(_1421_),
    .B1(_1346_),
    .X(_1422_));
 sky130_fd_sc_hd__or2_1 _3128_ (.A(_1339_),
    .B(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__a21oi_1 _3129_ (.A1(_1337_),
    .A2(_1423_),
    .B1(_1335_),
    .Y(_1424_));
 sky130_fd_sc_hd__a31o_1 _3130_ (.A1(_1335_),
    .A2(_1337_),
    .A3(_1423_),
    .B1(net177),
    .X(_1425_));
 sky130_fd_sc_hd__a2bb2o_1 _3131_ (.A1_N(_1424_),
    .A2_N(_1425_),
    .B1(\cordic_inst.cordic_inst.x[23] ),
    .B2(net169),
    .X(_0521_));
 sky130_fd_sc_hd__nand2_1 _3132_ (.A(_1339_),
    .B(_1422_),
    .Y(_1426_));
 sky130_fd_sc_hd__a32o_1 _3133_ (.A1(net183),
    .A2(_1423_),
    .A3(_1426_),
    .B1(net165),
    .B2(\cordic_inst.cordic_inst.x[22] ),
    .X(_0520_));
 sky130_fd_sc_hd__a21oi_1 _3134_ (.A1(_1341_),
    .A2(_1421_),
    .B1(_1348_),
    .Y(_1427_));
 sky130_fd_sc_hd__a31o_1 _3135_ (.A1(_1341_),
    .A2(_1348_),
    .A3(_1421_),
    .B1(net177),
    .X(_1428_));
 sky130_fd_sc_hd__a2bb2o_1 _3136_ (.A1_N(_1427_),
    .A2_N(_1428_),
    .B1(\cordic_inst.cordic_inst.x[21] ),
    .B2(net165),
    .X(_0519_));
 sky130_fd_sc_hd__nand3_1 _3137_ (.A(_1343_),
    .B(_1375_),
    .C(_1420_),
    .Y(_1429_));
 sky130_fd_sc_hd__a32o_1 _3138_ (.A1(net183),
    .A2(_1421_),
    .A3(_1429_),
    .B1(net165),
    .B2(\cordic_inst.cordic_inst.x[20] ),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_1 _3139_ (.A(_1332_),
    .B(_1361_),
    .Y(_1430_));
 sky130_fd_sc_hd__a21o_1 _3140_ (.A1(_1373_),
    .A2(_1430_),
    .B1(_1365_),
    .X(_1431_));
 sky130_fd_sc_hd__or2_1 _3141_ (.A(_1358_),
    .B(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a21oi_1 _3142_ (.A1(_1357_),
    .A2(_1432_),
    .B1(_1355_),
    .Y(_1433_));
 sky130_fd_sc_hd__a31o_1 _3143_ (.A1(_1355_),
    .A2(_1357_),
    .A3(_1432_),
    .B1(net177),
    .X(_1434_));
 sky130_fd_sc_hd__a2bb2o_1 _3144_ (.A1_N(_1433_),
    .A2_N(_1434_),
    .B1(\cordic_inst.cordic_inst.x[19] ),
    .B2(net167),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_1 _3145_ (.A(_1358_),
    .B(_1431_),
    .Y(_1435_));
 sky130_fd_sc_hd__a32o_1 _3146_ (.A1(net185),
    .A2(_1432_),
    .A3(_1435_),
    .B1(net167),
    .B2(\cordic_inst.cordic_inst.x[18] ),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _3147_ (.A1(\cordic_inst.cordic_inst.x[16] ),
    .A2(_1360_),
    .B1(_1361_),
    .B2(_1332_),
    .X(_1436_));
 sky130_fd_sc_hd__xnor2_1 _3148_ (.A(_1367_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__a22o_1 _3149_ (.A1(\cordic_inst.cordic_inst.x[17] ),
    .A2(net166),
    .B1(_1437_),
    .B2(net184),
    .X(_0515_));
 sky130_fd_sc_hd__or2_1 _3150_ (.A(_1332_),
    .B(_1361_),
    .X(_1438_));
 sky130_fd_sc_hd__a32o_1 _3151_ (.A1(net184),
    .A2(_1430_),
    .A3(_1438_),
    .B1(net167),
    .B2(\cordic_inst.cordic_inst.x[16] ),
    .X(_0514_));
 sky130_fd_sc_hd__nand2_1 _3152_ (.A(_1287_),
    .B(_1290_),
    .Y(_1439_));
 sky130_fd_sc_hd__and3_1 _3153_ (.A(_1287_),
    .B(_1290_),
    .C(_1294_),
    .X(_1440_));
 sky130_fd_sc_hd__or3_1 _3154_ (.A(_1293_),
    .B(_1323_),
    .C(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__o21a_1 _3155_ (.A1(_1318_),
    .A2(_1441_),
    .B1(_1329_),
    .X(_1442_));
 sky130_fd_sc_hd__nor2_1 _3156_ (.A(_1311_),
    .B(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__o21a_1 _3157_ (.A1(_1326_),
    .A2(_1443_),
    .B1(_1307_),
    .X(_1444_));
 sky130_fd_sc_hd__nand2_1 _3158_ (.A(_1303_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__a21oi_1 _3159_ (.A1(_1302_),
    .A2(_1445_),
    .B1(_1299_),
    .Y(_1446_));
 sky130_fd_sc_hd__a31o_1 _3160_ (.A1(_1299_),
    .A2(_1302_),
    .A3(_1445_),
    .B1(net177),
    .X(_1447_));
 sky130_fd_sc_hd__o22a_1 _3161_ (.A1(\cordic_inst.cordic_inst.x[15] ),
    .A2(\cordic_inst.cordic_inst.next_state[1] ),
    .B1(_1446_),
    .B2(_1447_),
    .X(_0513_));
 sky130_fd_sc_hd__or2_1 _3162_ (.A(_1303_),
    .B(_1444_),
    .X(_1448_));
 sky130_fd_sc_hd__a32o_1 _3163_ (.A1(net185),
    .A2(_1445_),
    .A3(_1448_),
    .B1(net168),
    .B2(\cordic_inst.cordic_inst.x[14] ),
    .X(_0512_));
 sky130_fd_sc_hd__a21oi_1 _3164_ (.A1(\cordic_inst.cordic_inst.x[12] ),
    .A2(_1310_),
    .B1(_1443_),
    .Y(_1449_));
 sky130_fd_sc_hd__xnor2_1 _3165_ (.A(_1309_),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__a22o_1 _3166_ (.A1(\cordic_inst.cordic_inst.x[13] ),
    .A2(net168),
    .B1(_1450_),
    .B2(net185),
    .X(_0511_));
 sky130_fd_sc_hd__xnor2_1 _3167_ (.A(_1312_),
    .B(_1442_),
    .Y(_1451_));
 sky130_fd_sc_hd__o22a_1 _3168_ (.A1(\cordic_inst.cordic_inst.x[12] ),
    .A2(\cordic_inst.cordic_inst.next_state[1] ),
    .B1(_1451_),
    .B2(net178),
    .X(_0510_));
 sky130_fd_sc_hd__a21boi_1 _3169_ (.A1(_1321_),
    .A2(_1441_),
    .B1_N(_1318_),
    .Y(_1452_));
 sky130_fd_sc_hd__and3b_1 _3170_ (.A_N(_1318_),
    .B(_1321_),
    .C(_1441_),
    .X(_1453_));
 sky130_fd_sc_hd__o32a_1 _3171_ (.A1(net178),
    .A2(_1452_),
    .A3(_1453_),
    .B1(\cordic_inst.cordic_inst.next_state[1] ),
    .B2(\cordic_inst.cordic_inst.x[11] ),
    .X(_0509_));
 sky130_fd_sc_hd__o21ai_1 _3172_ (.A1(_1293_),
    .A2(_1440_),
    .B1(_1323_),
    .Y(_1454_));
 sky130_fd_sc_hd__a32o_1 _3173_ (.A1(net185),
    .A2(_1441_),
    .A3(_1454_),
    .B1(net168),
    .B2(\cordic_inst.cordic_inst.x[10] ),
    .X(_0508_));
 sky130_fd_sc_hd__nor2_1 _3174_ (.A(_1295_),
    .B(_1439_),
    .Y(_1455_));
 sky130_fd_sc_hd__a21o_1 _3175_ (.A1(_1295_),
    .A2(_1439_),
    .B1(net178),
    .X(_1456_));
 sky130_fd_sc_hd__o22a_1 _3176_ (.A1(\cordic_inst.cordic_inst.x[9] ),
    .A2(net158),
    .B1(_1455_),
    .B2(_1456_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _3177_ (.A(_1284_),
    .B(_1289_),
    .Y(_1457_));
 sky130_fd_sc_hd__and2_1 _3178_ (.A(_1290_),
    .B(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__o22a_1 _3179_ (.A1(\cordic_inst.cordic_inst.x[8] ),
    .A2(net158),
    .B1(_1458_),
    .B2(net178),
    .X(_0506_));
 sky130_fd_sc_hd__a21oi_1 _3180_ (.A1(_1247_),
    .A2(_1282_),
    .B1(_1283_),
    .Y(_1459_));
 sky130_fd_sc_hd__a31o_1 _3181_ (.A1(_1247_),
    .A2(_1282_),
    .A3(_1283_),
    .B1(net177),
    .X(_1460_));
 sky130_fd_sc_hd__a2bb2o_1 _3182_ (.A1_N(_1459_),
    .A2_N(_1460_),
    .B1(\cordic_inst.cordic_inst.x[7] ),
    .B2(net168),
    .X(_0505_));
 sky130_fd_sc_hd__xnor2_1 _3183_ (.A(_1249_),
    .B(_1281_),
    .Y(_1461_));
 sky130_fd_sc_hd__o2bb2a_1 _3184_ (.A1_N(net183),
    .A2_N(_1461_),
    .B1(net158),
    .B2(\cordic_inst.cordic_inst.x[6] ),
    .X(_0504_));
 sky130_fd_sc_hd__nor2_1 _3185_ (.A(_1279_),
    .B(_1280_),
    .Y(_1462_));
 sky130_fd_sc_hd__a21o_1 _3186_ (.A1(_1279_),
    .A2(_1280_),
    .B1(net177),
    .X(_1463_));
 sky130_fd_sc_hd__o22a_1 _3187_ (.A1(\cordic_inst.cordic_inst.x[5] ),
    .A2(net158),
    .B1(_1462_),
    .B2(_1463_),
    .X(_0503_));
 sky130_fd_sc_hd__nand3_1 _3188_ (.A(_1260_),
    .B(_1263_),
    .C(_1277_),
    .Y(_1464_));
 sky130_fd_sc_hd__and2_1 _3189_ (.A(_1278_),
    .B(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__o22a_1 _3190_ (.A1(\cordic_inst.cordic_inst.x[4] ),
    .A2(net158),
    .B1(_1465_),
    .B2(net177),
    .X(_0502_));
 sky130_fd_sc_hd__nand3_1 _3191_ (.A(_1266_),
    .B(_1274_),
    .C(_1276_),
    .Y(_1466_));
 sky130_fd_sc_hd__a32o_1 _3192_ (.A1(net183),
    .A2(_1277_),
    .A3(_1466_),
    .B1(net165),
    .B2(\cordic_inst.cordic_inst.x[3] ),
    .X(_0501_));
 sky130_fd_sc_hd__nand3_1 _3193_ (.A(_1269_),
    .B(_1272_),
    .C(_1273_),
    .Y(_1467_));
 sky130_fd_sc_hd__and2_1 _3194_ (.A(_1274_),
    .B(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__o22a_1 _3195_ (.A1(\cordic_inst.cordic_inst.x[2] ),
    .A2(net158),
    .B1(_1468_),
    .B2(net176),
    .X(_0500_));
 sky130_fd_sc_hd__nand2b_1 _3196_ (.A_N(_1271_),
    .B(_1270_),
    .Y(_1469_));
 sky130_fd_sc_hd__a32o_1 _3197_ (.A1(net181),
    .A2(_1272_),
    .A3(_1469_),
    .B1(net165),
    .B2(\cordic_inst.cordic_inst.x[1] ),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_1 _3198_ (.A(net180),
    .B(_1148_),
    .Y(_1470_));
 sky130_fd_sc_hd__nor2_1 _3199_ (.A(_0603_),
    .B(net174),
    .Y(_1471_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(_0603_),
    .A1(_1471_),
    .S(_1470_),
    .X(_0498_));
 sky130_fd_sc_hd__nand2_1 _3201_ (.A(\cordic_inst.cordic_inst.state[1] ),
    .B(\cordic_inst.cordic_inst.state[0] ),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(net263),
    .A1(\cordic_inst.cordic_inst.sin_out[31] ),
    .S(net207),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(\cordic_inst.cordic_inst.y[30] ),
    .A1(\cordic_inst.cordic_inst.sin_out[30] ),
    .S(net209),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(\cordic_inst.cordic_inst.y[29] ),
    .A1(\cordic_inst.cordic_inst.sin_out[29] ),
    .S(net207),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(\cordic_inst.cordic_inst.y[28] ),
    .A1(\cordic_inst.cordic_inst.sin_out[28] ),
    .S(net207),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(\cordic_inst.cordic_inst.y[27] ),
    .A1(\cordic_inst.cordic_inst.sin_out[27] ),
    .S(net209),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(\cordic_inst.cordic_inst.y[26] ),
    .A1(\cordic_inst.cordic_inst.sin_out[26] ),
    .S(net209),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(\cordic_inst.cordic_inst.y[25] ),
    .A1(\cordic_inst.cordic_inst.sin_out[25] ),
    .S(net209),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(\cordic_inst.cordic_inst.y[24] ),
    .A1(\cordic_inst.cordic_inst.sin_out[24] ),
    .S(net208),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _3210_ (.A0(\cordic_inst.cordic_inst.y[23] ),
    .A1(\cordic_inst.cordic_inst.sin_out[23] ),
    .S(net208),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(\cordic_inst.cordic_inst.y[22] ),
    .A1(\cordic_inst.cordic_inst.sin_out[22] ),
    .S(net208),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(\cordic_inst.cordic_inst.y[21] ),
    .A1(\cordic_inst.cordic_inst.sin_out[21] ),
    .S(net214),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(\cordic_inst.cordic_inst.y[20] ),
    .A1(\cordic_inst.cordic_inst.sin_out[20] ),
    .S(net214),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(\cordic_inst.cordic_inst.y[19] ),
    .A1(\cordic_inst.cordic_inst.sin_out[19] ),
    .S(net214),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\cordic_inst.cordic_inst.y[18] ),
    .A1(\cordic_inst.cordic_inst.sin_out[18] ),
    .S(net212),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(\cordic_inst.cordic_inst.y[17] ),
    .A1(\cordic_inst.cordic_inst.sin_out[17] ),
    .S(net212),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(\cordic_inst.cordic_inst.y[16] ),
    .A1(\cordic_inst.cordic_inst.sin_out[16] ),
    .S(net213),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(\cordic_inst.cordic_inst.y[15] ),
    .A1(\cordic_inst.cordic_inst.sin_out[15] ),
    .S(net213),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(\cordic_inst.cordic_inst.y[14] ),
    .A1(\cordic_inst.cordic_inst.sin_out[14] ),
    .S(net212),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(\cordic_inst.cordic_inst.y[13] ),
    .A1(\cordic_inst.cordic_inst.sin_out[13] ),
    .S(net213),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(\cordic_inst.cordic_inst.y[12] ),
    .A1(\cordic_inst.cordic_inst.sin_out[12] ),
    .S(net210),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(\cordic_inst.cordic_inst.y[11] ),
    .A1(\cordic_inst.cordic_inst.sin_out[11] ),
    .S(net210),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(\cordic_inst.cordic_inst.y[10] ),
    .A1(\cordic_inst.cordic_inst.sin_out[10] ),
    .S(net211),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(\cordic_inst.cordic_inst.y[9] ),
    .A1(\cordic_inst.cordic_inst.sin_out[9] ),
    .S(net210),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(\cordic_inst.cordic_inst.y[8] ),
    .A1(\cordic_inst.cordic_inst.sin_out[8] ),
    .S(net210),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(\cordic_inst.cordic_inst.y[7] ),
    .A1(\cordic_inst.cordic_inst.sin_out[7] ),
    .S(net210),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(\cordic_inst.cordic_inst.y[6] ),
    .A1(\cordic_inst.cordic_inst.sin_out[6] ),
    .S(net211),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(\cordic_inst.cordic_inst.y[5] ),
    .A1(\cordic_inst.cordic_inst.sin_out[5] ),
    .S(net211),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(\cordic_inst.cordic_inst.y[4] ),
    .A1(\cordic_inst.cordic_inst.sin_out[4] ),
    .S(net211),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(\cordic_inst.cordic_inst.y[3] ),
    .A1(\cordic_inst.cordic_inst.sin_out[3] ),
    .S(net214),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(\cordic_inst.cordic_inst.y[2] ),
    .A1(\cordic_inst.cordic_inst.sin_out[2] ),
    .S(net214),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(\cordic_inst.cordic_inst.y[1] ),
    .A1(\cordic_inst.cordic_inst.sin_out[1] ),
    .S(net214),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(\cordic_inst.cordic_inst.y[0] ),
    .A1(\cordic_inst.cordic_inst.sin_out[0] ),
    .S(net208),
    .X(_0466_));
 sky130_fd_sc_hd__nand2_1 _3234_ (.A(net249),
    .B(\cordic_inst.cordic_inst.z[30] ),
    .Y(_1473_));
 sky130_fd_sc_hd__xnor2_1 _3235_ (.A(net268),
    .B(\cordic_inst.cordic_inst.z[30] ),
    .Y(_1474_));
 sky130_fd_sc_hd__xnor2_1 _3236_ (.A(net268),
    .B(\cordic_inst.cordic_inst.z[29] ),
    .Y(_1475_));
 sky130_fd_sc_hd__inv_2 _3237_ (.A(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__xor2_1 _3238_ (.A(net268),
    .B(\cordic_inst.cordic_inst.z[28] ),
    .X(_1477_));
 sky130_fd_sc_hd__nand2_1 _3239_ (.A(net248),
    .B(\cordic_inst.cordic_inst.z[24] ),
    .Y(_1478_));
 sky130_fd_sc_hd__or2_1 _3240_ (.A(net248),
    .B(\cordic_inst.cordic_inst.z[24] ),
    .X(_1479_));
 sky130_fd_sc_hd__nand2_1 _3241_ (.A(_1478_),
    .B(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2_2 _3242_ (.A(net268),
    .B(_0714_),
    .Y(_1481_));
 sky130_fd_sc_hd__nor2_1 _3243_ (.A(net268),
    .B(_0714_),
    .Y(_1482_));
 sky130_fd_sc_hd__inv_2 _3244_ (.A(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__and3_1 _3245_ (.A(\cordic_inst.cordic_inst.z[21] ),
    .B(_1481_),
    .C(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__a21oi_1 _3246_ (.A1(_1481_),
    .A2(_1483_),
    .B1(\cordic_inst.cordic_inst.z[21] ),
    .Y(_1485_));
 sky130_fd_sc_hd__or2_1 _3247_ (.A(_1484_),
    .B(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__xnor2_1 _3248_ (.A(net268),
    .B(_0708_),
    .Y(_1487_));
 sky130_fd_sc_hd__nand2_1 _3249_ (.A(\cordic_inst.cordic_inst.z[20] ),
    .B(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__or2_1 _3250_ (.A(\cordic_inst.cordic_inst.z[20] ),
    .B(_1487_),
    .X(_1489_));
 sky130_fd_sc_hd__nand2_1 _3251_ (.A(_1488_),
    .B(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__and2_1 _3252_ (.A(net248),
    .B(\cordic_inst.cordic_inst.z[22] ),
    .X(_1491_));
 sky130_fd_sc_hd__nor2_1 _3253_ (.A(net248),
    .B(\cordic_inst.cordic_inst.z[22] ),
    .Y(_1492_));
 sky130_fd_sc_hd__or2_1 _3254_ (.A(_1491_),
    .B(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__xnor2_1 _3255_ (.A(net268),
    .B(\cordic_inst.cordic_inst.z[23] ),
    .Y(_1494_));
 sky130_fd_sc_hd__or3b_1 _3256_ (.A(_1491_),
    .B(_1492_),
    .C_N(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__or3_1 _3257_ (.A(_1486_),
    .B(_1490_),
    .C(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__o21ba_1 _3258_ (.A1(_1485_),
    .A2(_1488_),
    .B1_N(_1484_),
    .X(_1497_));
 sky130_fd_sc_hd__nor2_1 _3259_ (.A(net237),
    .B(net232),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2_1 _3260_ (.A(net288),
    .B(net294),
    .Y(_1499_));
 sky130_fd_sc_hd__nand2_1 _3261_ (.A(net294),
    .B(net303),
    .Y(_1500_));
 sky130_fd_sc_hd__a21oi_1 _3262_ (.A1(_1499_),
    .A2(_1500_),
    .B1(net281),
    .Y(_1501_));
 sky130_fd_sc_hd__nor3_1 _3263_ (.A(net288),
    .B(net294),
    .C(net302),
    .Y(_1502_));
 sky130_fd_sc_hd__a21oi_1 _3264_ (.A1(net280),
    .A2(net206),
    .B1(_1501_),
    .Y(_1503_));
 sky130_fd_sc_hd__or2_1 _3265_ (.A(net248),
    .B(net206),
    .X(_1504_));
 sky130_fd_sc_hd__o22a_1 _3266_ (.A1(net267),
    .A2(_1503_),
    .B1(_1504_),
    .B2(_1501_),
    .X(_1505_));
 sky130_fd_sc_hd__and2_1 _3267_ (.A(\cordic_inst.cordic_inst.z[13] ),
    .B(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__or2_1 _3268_ (.A(net248),
    .B(_0705_),
    .X(_1507_));
 sky130_fd_sc_hd__nand2_1 _3269_ (.A(net222),
    .B(_0707_),
    .Y(_1508_));
 sky130_fd_sc_hd__xor2_1 _3270_ (.A(net294),
    .B(net303),
    .X(_1509_));
 sky130_fd_sc_hd__a22o_1 _3271_ (.A1(net222),
    .A2(_0707_),
    .B1(_1509_),
    .B2(net220),
    .X(_1510_));
 sky130_fd_sc_hd__o21ai_1 _3272_ (.A1(net289),
    .A2(net294),
    .B1(net280),
    .Y(_1511_));
 sky130_fd_sc_hd__nand2b_1 _3273_ (.A_N(_1510_),
    .B(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(net267),
    .A1(_1507_),
    .S(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__nand2_1 _3275_ (.A(\cordic_inst.cordic_inst.z[12] ),
    .B(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__and2b_1 _3276_ (.A_N(_1506_),
    .B(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__nand2_1 _3277_ (.A(net220),
    .B(_0712_),
    .Y(_1516_));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(net267),
    .A1(_1481_),
    .S(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__and2_1 _3279_ (.A(\cordic_inst.cordic_inst.z[14] ),
    .B(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__nor2_1 _3280_ (.A(\cordic_inst.cordic_inst.z[14] ),
    .B(_1517_),
    .Y(_1519_));
 sky130_fd_sc_hd__or2_1 _3281_ (.A(_1518_),
    .B(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__or2_1 _3282_ (.A(net237),
    .B(net303),
    .X(_1521_));
 sky130_fd_sc_hd__inv_2 _3283_ (.A(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__a21o_1 _3284_ (.A1(_0707_),
    .A2(_1521_),
    .B1(net280),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _3285_ (.A0(net267),
    .A1(_1481_),
    .S(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__or2_1 _3286_ (.A(\cordic_inst.cordic_inst.z[15] ),
    .B(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__nand2_1 _3287_ (.A(\cordic_inst.cordic_inst.z[15] ),
    .B(_1524_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _3288_ (.A(_1525_),
    .B(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__nor2_1 _3289_ (.A(_1520_),
    .B(_1527_),
    .Y(_1528_));
 sky130_fd_sc_hd__inv_2 _3290_ (.A(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__nor2_1 _3291_ (.A(\cordic_inst.cordic_inst.z[13] ),
    .B(_1505_),
    .Y(_1530_));
 sky130_fd_sc_hd__nand2_1 _3292_ (.A(_1518_),
    .B(_1525_),
    .Y(_1531_));
 sky130_fd_sc_hd__o311a_1 _3293_ (.A1(_1515_),
    .A2(_1529_),
    .A3(_1530_),
    .B1(_1531_),
    .C1(_1526_),
    .X(_1532_));
 sky130_fd_sc_hd__or2_1 _3294_ (.A(_1506_),
    .B(_1530_),
    .X(_1533_));
 sky130_fd_sc_hd__or2_1 _3295_ (.A(\cordic_inst.cordic_inst.z[12] ),
    .B(_1513_),
    .X(_1534_));
 sky130_fd_sc_hd__nand2_1 _3296_ (.A(_1514_),
    .B(_1534_),
    .Y(_1535_));
 sky130_fd_sc_hd__a221o_1 _3297_ (.A1(net294),
    .A2(net302),
    .B1(_0706_),
    .B2(net288),
    .C1(_0713_),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(net266),
    .A1(_1504_),
    .S(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__or2_1 _3299_ (.A(\cordic_inst.cordic_inst.z[11] ),
    .B(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__nand2_1 _3300_ (.A(\cordic_inst.cordic_inst.z[11] ),
    .B(_1537_),
    .Y(_1539_));
 sky130_fd_sc_hd__nand2_1 _3301_ (.A(_1538_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__nand2_1 _3302_ (.A(net280),
    .B(net288),
    .Y(_1541_));
 sky130_fd_sc_hd__and4b_1 _3303_ (.A_N(net222),
    .B(_0706_),
    .C(_0712_),
    .D(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _3304_ (.A0(_1481_),
    .A1(net266),
    .S(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__and2_1 _3305_ (.A(\cordic_inst.cordic_inst.z[10] ),
    .B(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__or2_1 _3306_ (.A(\cordic_inst.cordic_inst.z[10] ),
    .B(_1543_),
    .X(_1545_));
 sky130_fd_sc_hd__nand2b_1 _3307_ (.A_N(_1544_),
    .B(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__nor2_1 _3308_ (.A(_1540_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__a311o_1 _3309_ (.A1(net288),
    .A2(_0706_),
    .A3(_0712_),
    .B1(net222),
    .C1(_0705_),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _3310_ (.A0(net266),
    .A1(_1481_),
    .S(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__or2_1 _3311_ (.A(\cordic_inst.cordic_inst.z[9] ),
    .B(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__inv_2 _3312_ (.A(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__a31o_1 _3313_ (.A1(net281),
    .A2(_0707_),
    .A3(_1521_),
    .B1(_1510_),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(net266),
    .A1(_1481_),
    .S(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__and2_1 _3315_ (.A(\cordic_inst.cordic_inst.z[7] ),
    .B(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__nor2_1 _3316_ (.A(\cordic_inst.cordic_inst.z[7] ),
    .B(_1553_),
    .Y(_1555_));
 sky130_fd_sc_hd__or2_1 _3317_ (.A(_1554_),
    .B(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__a21oi_1 _3318_ (.A1(net280),
    .A2(net237),
    .B1(_0712_),
    .Y(_1557_));
 sky130_fd_sc_hd__and2_1 _3319_ (.A(net237),
    .B(net302),
    .X(_1558_));
 sky130_fd_sc_hd__or3_1 _3320_ (.A(net220),
    .B(_1557_),
    .C(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(net266),
    .A1(_1504_),
    .S(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__and2_1 _3322_ (.A(\cordic_inst.cordic_inst.z[6] ),
    .B(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__nor2_1 _3323_ (.A(\cordic_inst.cordic_inst.z[6] ),
    .B(_1560_),
    .Y(_1562_));
 sky130_fd_sc_hd__or2_1 _3324_ (.A(_1561_),
    .B(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__or2_1 _3325_ (.A(net281),
    .B(_0707_),
    .X(_1564_));
 sky130_fd_sc_hd__o21ai_1 _3326_ (.A1(_1498_),
    .A2(_1558_),
    .B1(_0706_),
    .Y(_1565_));
 sky130_fd_sc_hd__and2_1 _3327_ (.A(_1564_),
    .B(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(net266),
    .A1(_1481_),
    .S(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__and2_1 _3329_ (.A(\cordic_inst.cordic_inst.z[5] ),
    .B(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__nor2_1 _3330_ (.A(\cordic_inst.cordic_inst.z[5] ),
    .B(_1567_),
    .Y(_1569_));
 sky130_fd_sc_hd__nor2_1 _3331_ (.A(_1568_),
    .B(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__nor2_1 _3332_ (.A(net302),
    .B(_0705_),
    .Y(_1571_));
 sky130_fd_sc_hd__o211a_1 _3333_ (.A1(net241),
    .A2(net294),
    .B1(net302),
    .C1(net288),
    .X(_1572_));
 sky130_fd_sc_hd__a31o_1 _3334_ (.A1(net280),
    .A2(_1499_),
    .A3(_1571_),
    .B1(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _3335_ (.A0(_1481_),
    .A1(net266),
    .S(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__nand2_1 _3336_ (.A(\cordic_inst.cordic_inst.z[4] ),
    .B(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__a21o_1 _3337_ (.A1(net296),
    .A2(net303),
    .B1(net289),
    .X(_1576_));
 sky130_fd_sc_hd__nor2_1 _3338_ (.A(_0711_),
    .B(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__nor2_1 _3339_ (.A(_1498_),
    .B(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__a32o_1 _3340_ (.A1(net281),
    .A2(_1521_),
    .A3(_1578_),
    .B1(net220),
    .B2(_1500_),
    .X(_1579_));
 sky130_fd_sc_hd__and3_1 _3341_ (.A(net293),
    .B(net295),
    .C(net306),
    .X(_1580_));
 sky130_fd_sc_hd__inv_2 _3342_ (.A(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__o32a_1 _3343_ (.A1(net281),
    .A2(_1577_),
    .A3(_1580_),
    .B1(_1511_),
    .B2(_1522_),
    .X(_1582_));
 sky130_fd_sc_hd__a211o_1 _3344_ (.A1(net288),
    .A2(_1509_),
    .B1(net206),
    .C1(net280),
    .X(_1583_));
 sky130_fd_sc_hd__nand2b_1 _3345_ (.A_N(_1511_),
    .B(_0707_),
    .Y(_1584_));
 sky130_fd_sc_hd__a21oi_1 _3346_ (.A1(_1583_),
    .A2(_1584_),
    .B1(net248),
    .Y(_1585_));
 sky130_fd_sc_hd__o21a_1 _3347_ (.A1(net241),
    .A2(net302),
    .B1(net288),
    .X(_1586_));
 sky130_fd_sc_hd__a21o_1 _3348_ (.A1(_1564_),
    .A2(_1586_),
    .B1(_1577_),
    .X(_1587_));
 sky130_fd_sc_hd__a21oi_1 _3349_ (.A1(net267),
    .A2(_1587_),
    .B1(_1585_),
    .Y(_1588_));
 sky130_fd_sc_hd__a21boi_1 _3350_ (.A1(net267),
    .A2(_1582_),
    .B1_N(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__xor2_1 _3351_ (.A(_1579_),
    .B(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__and2_1 _3352_ (.A(\cordic_inst.cordic_inst.z[3] ),
    .B(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__xnor2_1 _3353_ (.A(\cordic_inst.cordic_inst.z[3] ),
    .B(_1590_),
    .Y(_1592_));
 sky130_fd_sc_hd__xor2_1 _3354_ (.A(_1582_),
    .B(_1588_),
    .X(_1593_));
 sky130_fd_sc_hd__nand2_1 _3355_ (.A(\cordic_inst.cordic_inst.z[2] ),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__xnor2_1 _3356_ (.A(_1585_),
    .B(_1587_),
    .Y(_1595_));
 sky130_fd_sc_hd__and2_1 _3357_ (.A(\cordic_inst.cordic_inst.z[1] ),
    .B(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__a21oi_1 _3358_ (.A1(_1583_),
    .A2(_1584_),
    .B1(\cordic_inst.cordic_inst.z[0] ),
    .Y(_1597_));
 sky130_fd_sc_hd__xnor2_1 _3359_ (.A(\cordic_inst.cordic_inst.z[1] ),
    .B(_1595_),
    .Y(_1598_));
 sky130_fd_sc_hd__nor2_1 _3360_ (.A(_1597_),
    .B(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__xor2_1 _3361_ (.A(\cordic_inst.cordic_inst.z[2] ),
    .B(_1593_),
    .X(_1600_));
 sky130_fd_sc_hd__o21ai_1 _3362_ (.A1(_1596_),
    .A2(_1599_),
    .B1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__a21oi_1 _3363_ (.A1(_1594_),
    .A2(_1601_),
    .B1(_1592_),
    .Y(_1602_));
 sky130_fd_sc_hd__or2_1 _3364_ (.A(\cordic_inst.cordic_inst.z[4] ),
    .B(_1574_),
    .X(_1603_));
 sky130_fd_sc_hd__and2_1 _3365_ (.A(_1575_),
    .B(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__o21ai_1 _3366_ (.A1(_1591_),
    .A2(_1602_),
    .B1(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__a21boi_1 _3367_ (.A1(_1575_),
    .A2(_1605_),
    .B1_N(_1570_),
    .Y(_1606_));
 sky130_fd_sc_hd__nor2_1 _3368_ (.A(_1568_),
    .B(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__o21ba_1 _3369_ (.A1(_1568_),
    .A2(_1606_),
    .B1_N(_1563_),
    .X(_1608_));
 sky130_fd_sc_hd__nor2_1 _3370_ (.A(_1561_),
    .B(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__o21ba_1 _3371_ (.A1(_1561_),
    .A2(_1608_),
    .B1_N(_1556_),
    .X(_1610_));
 sky130_fd_sc_hd__or2_1 _3372_ (.A(_1554_),
    .B(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__or2_1 _3373_ (.A(net280),
    .B(net302),
    .X(_1612_));
 sky130_fd_sc_hd__o32a_1 _3374_ (.A1(_1498_),
    .A2(_1510_),
    .A3(_1577_),
    .B1(_1612_),
    .B2(net232),
    .X(_1613_));
 sky130_fd_sc_hd__nand2_1 _3375_ (.A(net266),
    .B(_0712_),
    .Y(_1614_));
 sky130_fd_sc_hd__mux2_1 _3376_ (.A0(net266),
    .A1(_1614_),
    .S(_1613_),
    .X(_1615_));
 sky130_fd_sc_hd__and2_1 _3377_ (.A(\cordic_inst.cordic_inst.z[8] ),
    .B(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__nor2_1 _3378_ (.A(\cordic_inst.cordic_inst.z[8] ),
    .B(_1615_),
    .Y(_1617_));
 sky130_fd_sc_hd__nor2_1 _3379_ (.A(_1616_),
    .B(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__and2_1 _3380_ (.A(_1611_),
    .B(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__and2_1 _3381_ (.A(\cordic_inst.cordic_inst.z[9] ),
    .B(_1549_),
    .X(_1620_));
 sky130_fd_sc_hd__a21oi_1 _3382_ (.A1(_1550_),
    .A2(_1616_),
    .B1(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__nor2_1 _3383_ (.A(_1551_),
    .B(_1620_),
    .Y(_1622_));
 sky130_fd_sc_hd__o31a_1 _3384_ (.A1(_1616_),
    .A2(_1619_),
    .A3(_1620_),
    .B1(_1550_),
    .X(_1623_));
 sky130_fd_sc_hd__nand2_1 _3385_ (.A(_1538_),
    .B(_1544_),
    .Y(_1624_));
 sky130_fd_sc_hd__o311a_1 _3386_ (.A1(_1540_),
    .A2(_1546_),
    .A3(_1621_),
    .B1(_1624_),
    .C1(_1539_),
    .X(_1625_));
 sky130_fd_sc_hd__o2111ai_2 _3387_ (.A1(_1554_),
    .A2(_1610_),
    .B1(_1618_),
    .C1(_1622_),
    .D1(_1547_),
    .Y(_1626_));
 sky130_fd_sc_hd__a21o_1 _3388_ (.A1(_1625_),
    .A2(_1626_),
    .B1(_1535_),
    .X(_1627_));
 sky130_fd_sc_hd__a2111o_1 _3389_ (.A1(_1625_),
    .A2(_1626_),
    .B1(_1529_),
    .C1(_1533_),
    .D1(_1535_),
    .X(_1628_));
 sky130_fd_sc_hd__nand2_1 _3390_ (.A(_1532_),
    .B(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__nand2_1 _3391_ (.A(net241),
    .B(_1578_),
    .Y(_1630_));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(_1507_),
    .A1(net266),
    .S(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__and2b_1 _3393_ (.A_N(_1631_),
    .B(\cordic_inst.cordic_inst.z[16] ),
    .X(_1632_));
 sky130_fd_sc_hd__and2b_1 _3394_ (.A_N(\cordic_inst.cordic_inst.z[16] ),
    .B(_1631_),
    .X(_1633_));
 sky130_fd_sc_hd__nor2_1 _3395_ (.A(_1632_),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__nor2_1 _3396_ (.A(net280),
    .B(_1576_),
    .Y(_1635_));
 sky130_fd_sc_hd__xnor2_1 _3397_ (.A(net267),
    .B(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__or2_1 _3398_ (.A(\cordic_inst.cordic_inst.z[19] ),
    .B(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__nand2_1 _3399_ (.A(\cordic_inst.cordic_inst.z[19] ),
    .B(_1636_),
    .Y(_1638_));
 sky130_fd_sc_hd__and2_1 _3400_ (.A(_1637_),
    .B(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__xnor2_1 _3401_ (.A(net249),
    .B(_1508_),
    .Y(_1640_));
 sky130_fd_sc_hd__xor2_1 _3402_ (.A(\cordic_inst.cordic_inst.z[18] ),
    .B(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__nand2_1 _3403_ (.A(_1639_),
    .B(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__a2111o_1 _3404_ (.A1(net288),
    .A2(net302),
    .B1(_1498_),
    .C1(_1502_),
    .D1(net280),
    .X(_1643_));
 sky130_fd_sc_hd__xnor2_1 _3405_ (.A(net248),
    .B(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__or2_1 _3406_ (.A(\cordic_inst.cordic_inst.z[17] ),
    .B(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__inv_2 _3407_ (.A(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__and2_1 _3408_ (.A(\cordic_inst.cordic_inst.z[17] ),
    .B(_1644_),
    .X(_1647_));
 sky130_fd_sc_hd__nor2_1 _3409_ (.A(_1646_),
    .B(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__or4bb_1 _3410_ (.A(_1647_),
    .B(_1642_),
    .C_N(_1634_),
    .D_N(_1645_),
    .X(_1649_));
 sky130_fd_sc_hd__a21o_1 _3411_ (.A1(_1532_),
    .A2(_1628_),
    .B1(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__o21a_1 _3412_ (.A1(_1632_),
    .A2(_1647_),
    .B1(_1645_),
    .X(_1651_));
 sky130_fd_sc_hd__inv_2 _3413_ (.A(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__a22o_1 _3414_ (.A1(\cordic_inst.cordic_inst.z[19] ),
    .A2(_1636_),
    .B1(_1640_),
    .B2(\cordic_inst.cordic_inst.z[18] ),
    .X(_1653_));
 sky130_fd_sc_hd__o2bb2a_1 _3415_ (.A1_N(_1637_),
    .A2_N(_1653_),
    .B1(_1652_),
    .B2(_1642_),
    .X(_1654_));
 sky130_fd_sc_hd__a211o_1 _3416_ (.A1(_1532_),
    .A2(_1628_),
    .B1(_1649_),
    .C1(_1496_),
    .X(_1655_));
 sky130_fd_sc_hd__o22ai_1 _3417_ (.A1(_1495_),
    .A2(_1497_),
    .B1(_1654_),
    .B2(_1496_),
    .Y(_1656_));
 sky130_fd_sc_hd__a211oi_1 _3418_ (.A1(net248),
    .A2(\cordic_inst.cordic_inst.z[23] ),
    .B1(_1491_),
    .C1(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__a21o_1 _3419_ (.A1(_1655_),
    .A2(_1657_),
    .B1(_1480_),
    .X(_1658_));
 sky130_fd_sc_hd__xor2_1 _3420_ (.A(net267),
    .B(\cordic_inst.cordic_inst.z[25] ),
    .X(_1659_));
 sky130_fd_sc_hd__xnor2_1 _3421_ (.A(net268),
    .B(\cordic_inst.cordic_inst.z[27] ),
    .Y(_1660_));
 sky130_fd_sc_hd__xnor2_1 _3422_ (.A(net268),
    .B(\cordic_inst.cordic_inst.z[26] ),
    .Y(_1661_));
 sky130_fd_sc_hd__nand2_1 _3423_ (.A(_1660_),
    .B(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__o21a_1 _3424_ (.A1(\cordic_inst.cordic_inst.z[25] ),
    .A2(\cordic_inst.cordic_inst.z[24] ),
    .B1(net248),
    .X(_1663_));
 sky130_fd_sc_hd__o21a_1 _3425_ (.A1(\cordic_inst.cordic_inst.z[27] ),
    .A2(\cordic_inst.cordic_inst.z[26] ),
    .B1(net249),
    .X(_1664_));
 sky130_fd_sc_hd__nor2_1 _3426_ (.A(_1663_),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__o31a_1 _3427_ (.A1(_1658_),
    .A2(_1659_),
    .A3(_1662_),
    .B1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__nor2_1 _3428_ (.A(_1477_),
    .B(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__o21ai_1 _3429_ (.A1(\cordic_inst.cordic_inst.z[29] ),
    .A2(\cordic_inst.cordic_inst.z[28] ),
    .B1(net249),
    .Y(_1668_));
 sky130_fd_sc_hd__o31ai_1 _3430_ (.A1(_1476_),
    .A2(_1477_),
    .A3(_1666_),
    .B1(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__a21oi_1 _3431_ (.A1(_1474_),
    .A2(_1669_),
    .B1(net176),
    .Y(_1670_));
 sky130_fd_sc_hd__a221o_1 _3432_ (.A1(_0614_),
    .A2(\cordic_inst.cordic_inst.angle[31] ),
    .B1(_1473_),
    .B2(_1670_),
    .C1(net162),
    .X(_1671_));
 sky130_fd_sc_hd__o21a_1 _3433_ (.A1(net268),
    .A2(net158),
    .B1(_1671_),
    .X(_0465_));
 sky130_fd_sc_hd__or2_1 _3434_ (.A(_1474_),
    .B(_1669_),
    .X(_1672_));
 sky130_fd_sc_hd__a221o_1 _3435_ (.A1(\cordic_inst.cordic_inst.angle[30] ),
    .A2(net176),
    .B1(_1670_),
    .B2(_1672_),
    .C1(net162),
    .X(_1673_));
 sky130_fd_sc_hd__o21a_1 _3436_ (.A1(\cordic_inst.cordic_inst.z[30] ),
    .A2(net158),
    .B1(_1673_),
    .X(_0464_));
 sky130_fd_sc_hd__a21oi_1 _3437_ (.A1(net249),
    .A2(\cordic_inst.cordic_inst.z[28] ),
    .B1(_1667_),
    .Y(_1674_));
 sky130_fd_sc_hd__xnor2_1 _3438_ (.A(_1475_),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__a22o_1 _3439_ (.A1(\cordic_inst.cordic_inst.angle[29] ),
    .A2(net174),
    .B1(net162),
    .B2(\cordic_inst.cordic_inst.z[29] ),
    .X(_1676_));
 sky130_fd_sc_hd__a21o_1 _3440_ (.A1(net181),
    .A2(_1675_),
    .B1(_1676_),
    .X(_0463_));
 sky130_fd_sc_hd__or2_1 _3441_ (.A(net176),
    .B(_1667_),
    .X(_1677_));
 sky130_fd_sc_hd__a21oi_1 _3442_ (.A1(_1477_),
    .A2(_1666_),
    .B1(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__a221o_1 _3443_ (.A1(\cordic_inst.cordic_inst.angle[28] ),
    .A2(net174),
    .B1(net162),
    .B2(\cordic_inst.cordic_inst.z[28] ),
    .C1(_1678_),
    .X(_0462_));
 sky130_fd_sc_hd__nor2_1 _3444_ (.A(_1658_),
    .B(_1659_),
    .Y(_1679_));
 sky130_fd_sc_hd__o21ai_1 _3445_ (.A1(_1663_),
    .A2(_1679_),
    .B1(_1661_),
    .Y(_1680_));
 sky130_fd_sc_hd__a21boi_1 _3446_ (.A1(net249),
    .A2(\cordic_inst.cordic_inst.z[26] ),
    .B1_N(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__xnor2_1 _3447_ (.A(_1660_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__a22o_1 _3448_ (.A1(\cordic_inst.cordic_inst.angle[27] ),
    .A2(net173),
    .B1(net161),
    .B2(\cordic_inst.cordic_inst.z[27] ),
    .X(_1683_));
 sky130_fd_sc_hd__a21o_1 _3449_ (.A1(net180),
    .A2(_1682_),
    .B1(_1683_),
    .X(_0461_));
 sky130_fd_sc_hd__or3_1 _3450_ (.A(_1661_),
    .B(_1663_),
    .C(_1679_),
    .X(_1684_));
 sky130_fd_sc_hd__a22o_1 _3451_ (.A1(\cordic_inst.cordic_inst.angle[26] ),
    .A2(net173),
    .B1(net161),
    .B2(\cordic_inst.cordic_inst.z[26] ),
    .X(_1685_));
 sky130_fd_sc_hd__a31o_1 _3452_ (.A1(net180),
    .A2(_1680_),
    .A3(_1684_),
    .B1(_1685_),
    .X(_0460_));
 sky130_fd_sc_hd__a21oi_1 _3453_ (.A1(_1478_),
    .A2(_1658_),
    .B1(_1659_),
    .Y(_1686_));
 sky130_fd_sc_hd__a31o_1 _3454_ (.A1(_1478_),
    .A2(_1658_),
    .A3(_1659_),
    .B1(net176),
    .X(_1687_));
 sky130_fd_sc_hd__nor2_1 _3455_ (.A(_1686_),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__a221o_1 _3456_ (.A1(\cordic_inst.cordic_inst.angle[25] ),
    .A2(net173),
    .B1(net161),
    .B2(\cordic_inst.cordic_inst.z[25] ),
    .C1(_1688_),
    .X(_0459_));
 sky130_fd_sc_hd__and3_1 _3457_ (.A(_1480_),
    .B(_1655_),
    .C(_1657_),
    .X(_1689_));
 sky130_fd_sc_hd__and3b_1 _3458_ (.A_N(_1689_),
    .B(net180),
    .C(_1658_),
    .X(_1690_));
 sky130_fd_sc_hd__a221o_1 _3459_ (.A1(\cordic_inst.cordic_inst.angle[24] ),
    .A2(net173),
    .B1(net161),
    .B2(\cordic_inst.cordic_inst.z[24] ),
    .C1(_1690_),
    .X(_0458_));
 sky130_fd_sc_hd__a21o_1 _3460_ (.A1(_1650_),
    .A2(_1654_),
    .B1(_1490_),
    .X(_1691_));
 sky130_fd_sc_hd__o21a_1 _3461_ (.A1(_1486_),
    .A2(_1691_),
    .B1(_1497_),
    .X(_1692_));
 sky130_fd_sc_hd__nor2_1 _3462_ (.A(_1493_),
    .B(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__o21ai_1 _3463_ (.A1(_1491_),
    .A2(_1693_),
    .B1(_1494_),
    .Y(_1694_));
 sky130_fd_sc_hd__or3_1 _3464_ (.A(_1491_),
    .B(_1494_),
    .C(_1693_),
    .X(_1695_));
 sky130_fd_sc_hd__a22o_1 _3465_ (.A1(\cordic_inst.cordic_inst.angle[23] ),
    .A2(net173),
    .B1(net161),
    .B2(\cordic_inst.cordic_inst.z[23] ),
    .X(_1696_));
 sky130_fd_sc_hd__a31o_1 _3466_ (.A1(net180),
    .A2(_1694_),
    .A3(_1695_),
    .B1(_1696_),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_1 _3467_ (.A(_1493_),
    .B(_1692_),
    .Y(_1697_));
 sky130_fd_sc_hd__and3b_1 _3468_ (.A_N(_1693_),
    .B(_1697_),
    .C(net180),
    .X(_1698_));
 sky130_fd_sc_hd__a221o_1 _3469_ (.A1(\cordic_inst.cordic_inst.angle[22] ),
    .A2(net173),
    .B1(net161),
    .B2(\cordic_inst.cordic_inst.z[22] ),
    .C1(_1698_),
    .X(_0456_));
 sky130_fd_sc_hd__nand3_1 _3470_ (.A(_1486_),
    .B(_1488_),
    .C(_1691_),
    .Y(_1699_));
 sky130_fd_sc_hd__a21o_1 _3471_ (.A1(_1488_),
    .A2(_1691_),
    .B1(_1486_),
    .X(_1700_));
 sky130_fd_sc_hd__a22o_1 _3472_ (.A1(\cordic_inst.cordic_inst.angle[21] ),
    .A2(net173),
    .B1(net162),
    .B2(\cordic_inst.cordic_inst.z[21] ),
    .X(_1701_));
 sky130_fd_sc_hd__a31o_1 _3473_ (.A1(net180),
    .A2(_1699_),
    .A3(_1700_),
    .B1(_1701_),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(net180),
    .B(_1691_),
    .Y(_1702_));
 sky130_fd_sc_hd__a31o_1 _3475_ (.A1(_1490_),
    .A2(_1650_),
    .A3(_1654_),
    .B1(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__a22oi_1 _3476_ (.A1(\cordic_inst.cordic_inst.angle[20] ),
    .A2(net173),
    .B1(net161),
    .B2(\cordic_inst.cordic_inst.z[20] ),
    .Y(_1704_));
 sky130_fd_sc_hd__nand2_1 _3477_ (.A(_1703_),
    .B(_1704_),
    .Y(_0454_));
 sky130_fd_sc_hd__and2_1 _3478_ (.A(_1629_),
    .B(_1634_),
    .X(_1705_));
 sky130_fd_sc_hd__o311a_1 _3479_ (.A1(_1632_),
    .A2(_1647_),
    .A3(_1705_),
    .B1(_1641_),
    .C1(_1645_),
    .X(_1706_));
 sky130_fd_sc_hd__a21o_1 _3480_ (.A1(\cordic_inst.cordic_inst.z[18] ),
    .A2(_1640_),
    .B1(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__a21oi_1 _3481_ (.A1(_1639_),
    .A2(_1707_),
    .B1(net175),
    .Y(_1708_));
 sky130_fd_sc_hd__o21a_1 _3482_ (.A1(_1639_),
    .A2(_1707_),
    .B1(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__a221o_1 _3483_ (.A1(\cordic_inst.cordic_inst.angle[19] ),
    .A2(net173),
    .B1(net162),
    .B2(\cordic_inst.cordic_inst.z[19] ),
    .C1(_1709_),
    .X(_0453_));
 sky130_fd_sc_hd__a211o_1 _3484_ (.A1(_1648_),
    .A2(_1705_),
    .B1(_1651_),
    .C1(_1641_),
    .X(_1710_));
 sky130_fd_sc_hd__and3b_1 _3485_ (.A_N(_1706_),
    .B(_1710_),
    .C(net179),
    .X(_1711_));
 sky130_fd_sc_hd__a221o_1 _3486_ (.A1(\cordic_inst.cordic_inst.angle[18] ),
    .A2(net172),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[18] ),
    .C1(_1711_),
    .X(_0452_));
 sky130_fd_sc_hd__o21ai_1 _3487_ (.A1(_1632_),
    .A2(_1705_),
    .B1(_1648_),
    .Y(_1712_));
 sky130_fd_sc_hd__or3_1 _3488_ (.A(_1632_),
    .B(_1648_),
    .C(_1705_),
    .X(_1713_));
 sky130_fd_sc_hd__a22o_1 _3489_ (.A1(\cordic_inst.cordic_inst.angle[17] ),
    .A2(net172),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[17] ),
    .X(_1714_));
 sky130_fd_sc_hd__a31o_1 _3490_ (.A1(net179),
    .A2(_1712_),
    .A3(_1713_),
    .B1(_1714_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_1 _3491_ (.A(net175),
    .B(_1705_),
    .Y(_1715_));
 sky130_fd_sc_hd__o21a_1 _3492_ (.A1(_1629_),
    .A2(_1634_),
    .B1(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__a221o_1 _3493_ (.A1(\cordic_inst.cordic_inst.angle[16] ),
    .A2(net172),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[16] ),
    .C1(_1716_),
    .X(_0450_));
 sky130_fd_sc_hd__a21o_1 _3494_ (.A1(_1515_),
    .A2(_1627_),
    .B1(_1530_),
    .X(_1717_));
 sky130_fd_sc_hd__nor2_1 _3495_ (.A(_1520_),
    .B(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__nor2_1 _3496_ (.A(_1518_),
    .B(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__o21ai_1 _3497_ (.A1(_1527_),
    .A2(_1719_),
    .B1(net179),
    .Y(_1720_));
 sky130_fd_sc_hd__a21oi_1 _3498_ (.A1(_1527_),
    .A2(_1719_),
    .B1(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__a221o_1 _3499_ (.A1(\cordic_inst.cordic_inst.angle[15] ),
    .A2(net172),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[15] ),
    .C1(_1721_),
    .X(_0449_));
 sky130_fd_sc_hd__nor2_1 _3500_ (.A(net175),
    .B(_1718_),
    .Y(_1722_));
 sky130_fd_sc_hd__a21boi_1 _3501_ (.A1(_1520_),
    .A2(_1717_),
    .B1_N(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__a221o_1 _3502_ (.A1(\cordic_inst.cordic_inst.angle[14] ),
    .A2(net172),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[14] ),
    .C1(_1723_),
    .X(_0448_));
 sky130_fd_sc_hd__nand3_1 _3503_ (.A(_1514_),
    .B(_1533_),
    .C(_1627_),
    .Y(_1724_));
 sky130_fd_sc_hd__a21o_1 _3504_ (.A1(_1514_),
    .A2(_1627_),
    .B1(_1533_),
    .X(_1725_));
 sky130_fd_sc_hd__a22o_1 _3505_ (.A1(\cordic_inst.cordic_inst.angle[13] ),
    .A2(net172),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[13] ),
    .X(_1726_));
 sky130_fd_sc_hd__a31o_1 _3506_ (.A1(net179),
    .A2(_1724_),
    .A3(_1725_),
    .B1(_1726_),
    .X(_0447_));
 sky130_fd_sc_hd__and3_1 _3507_ (.A(_1535_),
    .B(_1625_),
    .C(_1626_),
    .X(_1727_));
 sky130_fd_sc_hd__and3b_1 _3508_ (.A_N(_1727_),
    .B(net179),
    .C(_1627_),
    .X(_1728_));
 sky130_fd_sc_hd__a221o_1 _3509_ (.A1(\cordic_inst.cordic_inst.angle[12] ),
    .A2(net172),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[12] ),
    .C1(_1728_),
    .X(_0446_));
 sky130_fd_sc_hd__a21oi_1 _3510_ (.A1(_1545_),
    .A2(_1623_),
    .B1(_1544_),
    .Y(_1729_));
 sky130_fd_sc_hd__a21o_1 _3511_ (.A1(_1540_),
    .A2(_1729_),
    .B1(net175),
    .X(_1730_));
 sky130_fd_sc_hd__o21ba_1 _3512_ (.A1(_1540_),
    .A2(_1729_),
    .B1_N(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__a221o_1 _3513_ (.A1(\cordic_inst.cordic_inst.angle[11] ),
    .A2(net171),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[11] ),
    .C1(_1731_),
    .X(_0445_));
 sky130_fd_sc_hd__xor2_1 _3514_ (.A(_1546_),
    .B(_1623_),
    .X(_1732_));
 sky130_fd_sc_hd__nor2_1 _3515_ (.A(net175),
    .B(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__a221o_1 _3516_ (.A1(\cordic_inst.cordic_inst.angle[10] ),
    .A2(net171),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[10] ),
    .C1(_1733_),
    .X(_0444_));
 sky130_fd_sc_hd__or3_1 _3517_ (.A(_1616_),
    .B(_1619_),
    .C(_1622_),
    .X(_1734_));
 sky130_fd_sc_hd__o21ai_1 _3518_ (.A1(_1616_),
    .A2(_1619_),
    .B1(_1622_),
    .Y(_1735_));
 sky130_fd_sc_hd__a22o_1 _3519_ (.A1(\cordic_inst.cordic_inst.angle[9] ),
    .A2(net171),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[9] ),
    .X(_1736_));
 sky130_fd_sc_hd__a31o_1 _3520_ (.A1(net182),
    .A2(_1734_),
    .A3(_1735_),
    .B1(_1736_),
    .X(_0443_));
 sky130_fd_sc_hd__nor2_1 _3521_ (.A(net176),
    .B(_1619_),
    .Y(_1737_));
 sky130_fd_sc_hd__o21a_1 _3522_ (.A1(_1611_),
    .A2(_1618_),
    .B1(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__a221o_1 _3523_ (.A1(\cordic_inst.cordic_inst.angle[8] ),
    .A2(net171),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[8] ),
    .C1(_1738_),
    .X(_0442_));
 sky130_fd_sc_hd__or2_1 _3524_ (.A(net175),
    .B(_1610_),
    .X(_1739_));
 sky130_fd_sc_hd__a21oi_1 _3525_ (.A1(_1556_),
    .A2(_1609_),
    .B1(_1739_),
    .Y(_1740_));
 sky130_fd_sc_hd__a221o_1 _3526_ (.A1(\cordic_inst.cordic_inst.angle[7] ),
    .A2(net171),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[7] ),
    .C1(_1740_),
    .X(_0441_));
 sky130_fd_sc_hd__or2_1 _3527_ (.A(net175),
    .B(_1608_),
    .X(_1741_));
 sky130_fd_sc_hd__a21oi_1 _3528_ (.A1(_1563_),
    .A2(_1607_),
    .B1(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__a221o_1 _3529_ (.A1(\cordic_inst.cordic_inst.angle[6] ),
    .A2(net171),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[6] ),
    .C1(_1742_),
    .X(_0440_));
 sky130_fd_sc_hd__and3b_1 _3530_ (.A_N(_1570_),
    .B(_1575_),
    .C(_1605_),
    .X(_1743_));
 sky130_fd_sc_hd__nor3_1 _3531_ (.A(net175),
    .B(_1606_),
    .C(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__a221o_1 _3532_ (.A1(\cordic_inst.cordic_inst.angle[5] ),
    .A2(net171),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[5] ),
    .C1(_1744_),
    .X(_0439_));
 sky130_fd_sc_hd__or3_1 _3533_ (.A(_1591_),
    .B(_1602_),
    .C(_1604_),
    .X(_1745_));
 sky130_fd_sc_hd__a22o_1 _3534_ (.A1(\cordic_inst.cordic_inst.angle[4] ),
    .A2(net171),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[4] ),
    .X(_1746_));
 sky130_fd_sc_hd__a31o_1 _3535_ (.A1(net182),
    .A2(_1605_),
    .A3(_1745_),
    .B1(_1746_),
    .X(_0438_));
 sky130_fd_sc_hd__and3_1 _3536_ (.A(_1592_),
    .B(_1594_),
    .C(_1601_),
    .X(_1747_));
 sky130_fd_sc_hd__a22oi_1 _3537_ (.A1(\cordic_inst.cordic_inst.angle[3] ),
    .A2(net171),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[3] ),
    .Y(_1748_));
 sky130_fd_sc_hd__o31ai_1 _3538_ (.A1(net175),
    .A2(_1602_),
    .A3(_1747_),
    .B1(_1748_),
    .Y(_0437_));
 sky130_fd_sc_hd__or3_1 _3539_ (.A(_1596_),
    .B(_1599_),
    .C(_1600_),
    .X(_1749_));
 sky130_fd_sc_hd__a22o_1 _3540_ (.A1(\cordic_inst.cordic_inst.angle[2] ),
    .A2(net172),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[2] ),
    .X(_1750_));
 sky130_fd_sc_hd__a31o_1 _3541_ (.A1(net182),
    .A2(_1601_),
    .A3(_1749_),
    .B1(_1750_),
    .X(_0436_));
 sky130_fd_sc_hd__or2_1 _3542_ (.A(net175),
    .B(_1599_),
    .X(_1751_));
 sky130_fd_sc_hd__a21oi_1 _3543_ (.A1(_1597_),
    .A2(_1598_),
    .B1(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__a221o_1 _3544_ (.A1(\cordic_inst.cordic_inst.angle[1] ),
    .A2(net172),
    .B1(net160),
    .B2(\cordic_inst.cordic_inst.z[1] ),
    .C1(_1752_),
    .X(_0435_));
 sky130_fd_sc_hd__and3_1 _3545_ (.A(\cordic_inst.cordic_inst.z[0] ),
    .B(_1583_),
    .C(_1584_),
    .X(_1753_));
 sky130_fd_sc_hd__o21a_1 _3546_ (.A1(_1597_),
    .A2(_1753_),
    .B1(net182),
    .X(_1754_));
 sky130_fd_sc_hd__a221o_1 _3547_ (.A1(\cordic_inst.cordic_inst.angle[0] ),
    .A2(net171),
    .B1(net159),
    .B2(\cordic_inst.cordic_inst.z[0] ),
    .C1(_1754_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(net265),
    .A1(\cordic_inst.cordic_inst.cos_out[31] ),
    .S(net207),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(\cordic_inst.cordic_inst.x[30] ),
    .A1(\cordic_inst.cordic_inst.cos_out[30] ),
    .S(net207),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(\cordic_inst.cordic_inst.x[29] ),
    .A1(\cordic_inst.cordic_inst.cos_out[29] ),
    .S(net207),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(\cordic_inst.cordic_inst.x[28] ),
    .A1(\cordic_inst.cordic_inst.cos_out[28] ),
    .S(net207),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(\cordic_inst.cordic_inst.x[27] ),
    .A1(\cordic_inst.cordic_inst.cos_out[27] ),
    .S(net207),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3553_ (.A0(\cordic_inst.cordic_inst.x[26] ),
    .A1(\cordic_inst.cordic_inst.cos_out[26] ),
    .S(net207),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _3554_ (.A0(\cordic_inst.cordic_inst.x[25] ),
    .A1(\cordic_inst.cordic_inst.cos_out[25] ),
    .S(net207),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(\cordic_inst.cordic_inst.x[24] ),
    .A1(\cordic_inst.cordic_inst.cos_out[24] ),
    .S(net209),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(\cordic_inst.cordic_inst.x[23] ),
    .A1(\cordic_inst.cordic_inst.cos_out[23] ),
    .S(net208),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(\cordic_inst.cordic_inst.x[22] ),
    .A1(\cordic_inst.cordic_inst.cos_out[22] ),
    .S(net208),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(\cordic_inst.cordic_inst.x[21] ),
    .A1(\cordic_inst.cordic_inst.cos_out[21] ),
    .S(net214),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(\cordic_inst.cordic_inst.x[20] ),
    .A1(\cordic_inst.cordic_inst.cos_out[20] ),
    .S(net214),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(\cordic_inst.cordic_inst.x[19] ),
    .A1(\cordic_inst.cordic_inst.cos_out[19] ),
    .S(net212),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(\cordic_inst.cordic_inst.x[18] ),
    .A1(\cordic_inst.cordic_inst.cos_out[18] ),
    .S(net212),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3562_ (.A0(\cordic_inst.cordic_inst.x[17] ),
    .A1(\cordic_inst.cordic_inst.cos_out[17] ),
    .S(net212),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(\cordic_inst.cordic_inst.x[16] ),
    .A1(\cordic_inst.cordic_inst.cos_out[16] ),
    .S(net212),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(\cordic_inst.cordic_inst.x[15] ),
    .A1(\cordic_inst.cordic_inst.cos_out[15] ),
    .S(net212),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(\cordic_inst.cordic_inst.x[14] ),
    .A1(\cordic_inst.cordic_inst.cos_out[14] ),
    .S(net212),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(\cordic_inst.cordic_inst.x[13] ),
    .A1(\cordic_inst.cordic_inst.cos_out[13] ),
    .S(net212),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3567_ (.A0(\cordic_inst.cordic_inst.x[12] ),
    .A1(\cordic_inst.cordic_inst.cos_out[12] ),
    .S(net210),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(\cordic_inst.cordic_inst.x[11] ),
    .A1(\cordic_inst.cordic_inst.cos_out[11] ),
    .S(net211),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3569_ (.A0(\cordic_inst.cordic_inst.x[10] ),
    .A1(\cordic_inst.cordic_inst.cos_out[10] ),
    .S(net211),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(\cordic_inst.cordic_inst.x[9] ),
    .A1(\cordic_inst.cordic_inst.cos_out[9] ),
    .S(net210),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _3571_ (.A0(\cordic_inst.cordic_inst.x[8] ),
    .A1(\cordic_inst.cordic_inst.cos_out[8] ),
    .S(net210),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(\cordic_inst.cordic_inst.x[7] ),
    .A1(\cordic_inst.cordic_inst.cos_out[7] ),
    .S(net210),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3573_ (.A0(\cordic_inst.cordic_inst.x[6] ),
    .A1(\cordic_inst.cordic_inst.cos_out[6] ),
    .S(net210),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\cordic_inst.cordic_inst.x[5] ),
    .A1(\cordic_inst.cordic_inst.cos_out[5] ),
    .S(net211),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(\cordic_inst.cordic_inst.x[4] ),
    .A1(\cordic_inst.cordic_inst.cos_out[4] ),
    .S(net211),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(\cordic_inst.cordic_inst.x[3] ),
    .A1(\cordic_inst.cordic_inst.cos_out[3] ),
    .S(net208),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(\cordic_inst.cordic_inst.x[2] ),
    .A1(\cordic_inst.cordic_inst.cos_out[2] ),
    .S(net208),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(\cordic_inst.cordic_inst.x[1] ),
    .A1(\cordic_inst.cordic_inst.cos_out[1] ),
    .S(net208),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(\cordic_inst.cordic_inst.x[0] ),
    .A1(\cordic_inst.cordic_inst.cos_out[0] ),
    .S(net208),
    .X(_0402_));
 sky130_fd_sc_hd__o21a_1 _3580_ (.A1(\cordic_inst.cordic_inst.done ),
    .A2(\cordic_inst.cordic_inst.state[0] ),
    .B1(\cordic_inst.cordic_inst.state[1] ),
    .X(_0401_));
 sky130_fd_sc_hd__o211a_1 _3581_ (.A1(\cordic_inst.cordic_inst.start ),
    .A2(\cordic_inst.state[2] ),
    .B1(_0620_),
    .C1(_0618_),
    .X(_0400_));
 sky130_fd_sc_hd__and3_1 _3582_ (.A(net282),
    .B(net180),
    .C(_1580_),
    .X(_1755_));
 sky130_fd_sc_hd__nor2_1 _3583_ (.A(net174),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(_1755_),
    .A1(_1756_),
    .S(net274),
    .X(_0390_));
 sky130_fd_sc_hd__a21o_1 _3585_ (.A1(net158),
    .A2(_1580_),
    .B1(net282),
    .X(_1757_));
 sky130_fd_sc_hd__and2_1 _3586_ (.A(_1756_),
    .B(_1757_),
    .X(_0389_));
 sky130_fd_sc_hd__a32o_1 _3587_ (.A1(net179),
    .A2(_1576_),
    .A3(_1581_),
    .B1(net161),
    .B2(net289),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _3588_ (.A1(net296),
    .A2(net161),
    .B1(_1509_),
    .B2(net179),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _3589_ (.A0(net180),
    .A1(net161),
    .S(net303),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _3590_ (.A(\cordic_inst.deg_handler_inst.theta_abs[0] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[1] ),
    .X(_1758_));
 sky130_fd_sc_hd__or3_1 _3591_ (.A(\cordic_inst.deg_handler_inst.theta_abs[0] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[1] ),
    .C(\cordic_inst.deg_handler_inst.theta_abs[2] ),
    .X(_1759_));
 sky130_fd_sc_hd__or2_1 _3592_ (.A(\cordic_inst.deg_handler_inst.theta_abs[3] ),
    .B(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__or2_1 _3593_ (.A(\cordic_inst.deg_handler_inst.theta_abs[4] ),
    .B(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__or2_1 _3594_ (.A(\cordic_inst.deg_handler_inst.theta_abs[5] ),
    .B(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__or2_1 _3595_ (.A(\cordic_inst.deg_handler_inst.theta_abs[6] ),
    .B(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__or2_1 _3596_ (.A(\cordic_inst.deg_handler_inst.theta_abs[7] ),
    .B(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__or2_1 _3597_ (.A(\cordic_inst.deg_handler_inst.theta_abs[8] ),
    .B(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__or2_1 _3598_ (.A(\cordic_inst.deg_handler_inst.theta_abs[9] ),
    .B(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__or2_1 _3599_ (.A(\cordic_inst.deg_handler_inst.theta_abs[10] ),
    .B(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__or2_1 _3600_ (.A(\cordic_inst.deg_handler_inst.theta_abs[11] ),
    .B(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__or2_1 _3601_ (.A(\cordic_inst.deg_handler_inst.theta_abs[12] ),
    .B(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__or2_1 _3602_ (.A(\cordic_inst.deg_handler_inst.theta_abs[13] ),
    .B(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__or2_1 _3603_ (.A(\cordic_inst.deg_handler_inst.theta_abs[14] ),
    .B(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__or2_1 _3604_ (.A(\cordic_inst.deg_handler_inst.theta_abs[15] ),
    .B(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__or2_1 _3605_ (.A(\cordic_inst.deg_handler_inst.theta_abs[16] ),
    .B(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(\cordic_inst.deg_handler_inst.theta_abs[17] ),
    .B(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__nand2_1 _3607_ (.A(_0615_),
    .B(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__a31o_1 _3608_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[19] ),
    .A2(\cordic_inst.deg_handler_inst.theta_abs[20] ),
    .A3(_1775_),
    .B1(\cordic_inst.deg_handler_inst.theta_abs[21] ),
    .X(_1776_));
 sky130_fd_sc_hd__or4_1 _3609_ (.A(\cordic_inst.deg_handler_inst.theta_abs[28] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[29] ),
    .C(\cordic_inst.deg_handler_inst.theta_abs[30] ),
    .D(\cordic_inst.deg_handler_inst.theta_abs[31] ),
    .X(_1777_));
 sky130_fd_sc_hd__or4_1 _3610_ (.A(\cordic_inst.deg_handler_inst.theta_abs[24] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[25] ),
    .C(\cordic_inst.deg_handler_inst.theta_abs[26] ),
    .D(\cordic_inst.deg_handler_inst.theta_abs[27] ),
    .X(_1778_));
 sky130_fd_sc_hd__or2_1 _3611_ (.A(_1777_),
    .B(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__a211oi_1 _3612_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[22] ),
    .A2(_1776_),
    .B1(_1779_),
    .C1(\cordic_inst.deg_handler_inst.theta_abs[23] ),
    .Y(_1780_));
 sky130_fd_sc_hd__or2_1 _3613_ (.A(\cordic_inst.deg_handler_inst.theta_abs[31] ),
    .B(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__nor2_1 _3614_ (.A(\cordic_inst.deg_handler_inst.theta_abs[18] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[19] ),
    .Y(_1782_));
 sky130_fd_sc_hd__nand2_1 _3615_ (.A(\cordic_inst.deg_handler_inst.theta_abs[20] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[21] ),
    .Y(_1783_));
 sky130_fd_sc_hd__o21ai_1 _3616_ (.A1(_1782_),
    .A2(_1783_),
    .B1(_0617_),
    .Y(_1784_));
 sky130_fd_sc_hd__a21o_1 _3617_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[23] ),
    .A2(_1784_),
    .B1(_1779_),
    .X(_1785_));
 sky130_fd_sc_hd__inv_2 _3618_ (.A(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__o21a_1 _3619_ (.A1(net153),
    .A2(_1786_),
    .B1(\cordic_inst.deg_handler_inst.theta_abs[0] ),
    .X(_0053_));
 sky130_fd_sc_hd__or2_2 _3620_ (.A(\cordic_inst.deg_handler_inst.theta_abs[17] ),
    .B(_1773_),
    .X(_1787_));
 sky130_fd_sc_hd__or4b_1 _3621_ (.A(_0615_),
    .B(\cordic_inst.deg_handler_inst.theta_abs[19] ),
    .C(\cordic_inst.deg_handler_inst.theta_abs[22] ),
    .D_N(\cordic_inst.deg_handler_inst.theta_abs[23] ),
    .X(_1788_));
 sky130_fd_sc_hd__or4_1 _3622_ (.A(_1779_),
    .B(_1783_),
    .C(_1787_),
    .D(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__a21oi_1 _3623_ (.A1(_1785_),
    .A2(_1789_),
    .B1(_1780_),
    .Y(_1790_));
 sky130_fd_sc_hd__inv_2 _3624_ (.A(net149),
    .Y(_0005_));
 sky130_fd_sc_hd__nand2_1 _3625_ (.A(\cordic_inst.deg_handler_inst.theta_abs[0] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[1] ),
    .Y(_1791_));
 sky130_fd_sc_hd__a32o_1 _3626_ (.A1(_1758_),
    .A2(net148),
    .A3(_1791_),
    .B1(net151),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[1] ),
    .X(_0064_));
 sky130_fd_sc_hd__nand2_1 _3627_ (.A(\cordic_inst.deg_handler_inst.theta_abs[2] ),
    .B(_1758_),
    .Y(_1792_));
 sky130_fd_sc_hd__a32o_1 _3628_ (.A1(_1759_),
    .A2(net148),
    .A3(_1792_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[2] ),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_1 _3629_ (.A(\cordic_inst.deg_handler_inst.theta_abs[3] ),
    .B(_1759_),
    .Y(_1793_));
 sky130_fd_sc_hd__a32o_1 _3630_ (.A1(_1760_),
    .A2(net148),
    .A3(_1793_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[3] ),
    .X(_0078_));
 sky130_fd_sc_hd__nand2_1 _3631_ (.A(\cordic_inst.deg_handler_inst.theta_abs[4] ),
    .B(_1760_),
    .Y(_1794_));
 sky130_fd_sc_hd__a32o_1 _3632_ (.A1(_1761_),
    .A2(net148),
    .A3(_1794_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[4] ),
    .X(_0079_));
 sky130_fd_sc_hd__nand2_1 _3633_ (.A(\cordic_inst.deg_handler_inst.theta_abs[5] ),
    .B(_1761_),
    .Y(_1795_));
 sky130_fd_sc_hd__a32o_1 _3634_ (.A1(_1762_),
    .A2(net147),
    .A3(_1795_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[5] ),
    .X(_0080_));
 sky130_fd_sc_hd__nand2_1 _3635_ (.A(\cordic_inst.deg_handler_inst.theta_abs[6] ),
    .B(_1762_),
    .Y(_1796_));
 sky130_fd_sc_hd__a32o_1 _3636_ (.A1(_1763_),
    .A2(net147),
    .A3(_1796_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[6] ),
    .X(_0081_));
 sky130_fd_sc_hd__nand2_1 _3637_ (.A(\cordic_inst.deg_handler_inst.theta_abs[7] ),
    .B(_1763_),
    .Y(_1797_));
 sky130_fd_sc_hd__a32o_1 _3638_ (.A1(_1764_),
    .A2(net147),
    .A3(_1797_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[7] ),
    .X(_0082_));
 sky130_fd_sc_hd__nand2_1 _3639_ (.A(\cordic_inst.deg_handler_inst.theta_abs[8] ),
    .B(_1764_),
    .Y(_1798_));
 sky130_fd_sc_hd__a32o_1 _3640_ (.A1(_1765_),
    .A2(net148),
    .A3(_1798_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[8] ),
    .X(_0083_));
 sky130_fd_sc_hd__nand2_1 _3641_ (.A(\cordic_inst.deg_handler_inst.theta_abs[9] ),
    .B(_1765_),
    .Y(_1799_));
 sky130_fd_sc_hd__a32o_1 _3642_ (.A1(_1766_),
    .A2(net148),
    .A3(_1799_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[9] ),
    .X(_0084_));
 sky130_fd_sc_hd__nand2_1 _3643_ (.A(\cordic_inst.deg_handler_inst.theta_abs[10] ),
    .B(_1766_),
    .Y(_1800_));
 sky130_fd_sc_hd__a32o_1 _3644_ (.A1(_1767_),
    .A2(net147),
    .A3(_1800_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[10] ),
    .X(_0054_));
 sky130_fd_sc_hd__nand2_1 _3645_ (.A(\cordic_inst.deg_handler_inst.theta_abs[11] ),
    .B(_1767_),
    .Y(_1801_));
 sky130_fd_sc_hd__a32o_1 _3646_ (.A1(_1768_),
    .A2(net147),
    .A3(_1801_),
    .B1(net150),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[11] ),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_1 _3647_ (.A(\cordic_inst.deg_handler_inst.theta_abs[12] ),
    .B(_1768_),
    .Y(_1802_));
 sky130_fd_sc_hd__a32o_1 _3648_ (.A1(_1769_),
    .A2(net147),
    .A3(_1802_),
    .B1(net151),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[12] ),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _3649_ (.A(\cordic_inst.deg_handler_inst.theta_abs[13] ),
    .B(_1769_),
    .Y(_1803_));
 sky130_fd_sc_hd__a32o_1 _3650_ (.A1(_1770_),
    .A2(net147),
    .A3(_1803_),
    .B1(net151),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[13] ),
    .X(_0057_));
 sky130_fd_sc_hd__nand2_1 _3651_ (.A(\cordic_inst.deg_handler_inst.theta_abs[14] ),
    .B(_1770_),
    .Y(_1804_));
 sky130_fd_sc_hd__a32o_1 _3652_ (.A1(_1771_),
    .A2(net147),
    .A3(_1804_),
    .B1(net151),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[14] ),
    .X(_0058_));
 sky130_fd_sc_hd__nand2_1 _3653_ (.A(\cordic_inst.deg_handler_inst.theta_abs[15] ),
    .B(_1771_),
    .Y(_1805_));
 sky130_fd_sc_hd__a32o_1 _3654_ (.A1(_1772_),
    .A2(net147),
    .A3(_1805_),
    .B1(net151),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[15] ),
    .X(_0059_));
 sky130_fd_sc_hd__nand2_1 _3655_ (.A(\cordic_inst.deg_handler_inst.theta_abs[16] ),
    .B(_1772_),
    .Y(_1806_));
 sky130_fd_sc_hd__a32o_1 _3656_ (.A1(_1773_),
    .A2(net147),
    .A3(_1806_),
    .B1(net151),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[16] ),
    .X(_0060_));
 sky130_fd_sc_hd__a32o_1 _3657_ (.A1(_1774_),
    .A2(_1787_),
    .A3(net149),
    .B1(net151),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[17] ),
    .X(_0061_));
 sky130_fd_sc_hd__xnor2_1 _3658_ (.A(\cordic_inst.deg_handler_inst.theta_abs[18] ),
    .B(_1787_),
    .Y(_1807_));
 sky130_fd_sc_hd__a22o_1 _3659_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[18] ),
    .A2(net152),
    .B1(net149),
    .B2(_1807_),
    .X(_0062_));
 sky130_fd_sc_hd__a21oi_2 _3660_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[18] ),
    .A2(_1787_),
    .B1(\cordic_inst.deg_handler_inst.theta_abs[19] ),
    .Y(_1808_));
 sky130_fd_sc_hd__and3_1 _3661_ (.A(\cordic_inst.deg_handler_inst.theta_abs[18] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[19] ),
    .C(_1787_),
    .X(_1809_));
 sky130_fd_sc_hd__nor2_1 _3662_ (.A(_1808_),
    .B(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__a22o_1 _3663_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[19] ),
    .A2(net152),
    .B1(net149),
    .B2(_1810_),
    .X(_0063_));
 sky130_fd_sc_hd__xnor2_1 _3664_ (.A(_0616_),
    .B(_1808_),
    .Y(_1811_));
 sky130_fd_sc_hd__a22o_1 _3665_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[20] ),
    .A2(net152),
    .B1(net149),
    .B2(_1811_),
    .X(_0065_));
 sky130_fd_sc_hd__o21bai_1 _3666_ (.A1(_0616_),
    .A2(_1808_),
    .B1_N(\cordic_inst.deg_handler_inst.theta_abs[21] ),
    .Y(_1812_));
 sky130_fd_sc_hd__o21ai_1 _3667_ (.A1(_1783_),
    .A2(_1808_),
    .B1(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__a22o_1 _3668_ (.A1(\cordic_inst.deg_handler_inst.theta_abs[21] ),
    .A2(net152),
    .B1(net149),
    .B2(_1813_),
    .X(_0066_));
 sky130_fd_sc_hd__or3_1 _3669_ (.A(_0617_),
    .B(_1783_),
    .C(_1808_),
    .X(_1814_));
 sky130_fd_sc_hd__o21ai_1 _3670_ (.A1(_1783_),
    .A2(_1808_),
    .B1(_0617_),
    .Y(_1815_));
 sky130_fd_sc_hd__a32o_1 _3671_ (.A1(net149),
    .A2(_1814_),
    .A3(_1815_),
    .B1(net152),
    .B2(\cordic_inst.deg_handler_inst.theta_abs[22] ),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _3672_ (.A(\cordic_inst.deg_handler_inst.theta_abs[23] ),
    .B(\cordic_inst.deg_handler_inst.theta_abs[31] ),
    .X(_0068_));
 sky130_fd_sc_hd__and2_1 _3673_ (.A(\cordic_inst.deg_handler_inst.theta_abs[24] ),
    .B(net152),
    .X(_0069_));
 sky130_fd_sc_hd__and2_1 _3674_ (.A(\cordic_inst.deg_handler_inst.theta_abs[25] ),
    .B(net153),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _3675_ (.A(\cordic_inst.deg_handler_inst.theta_abs[26] ),
    .B(net152),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _3676_ (.A(\cordic_inst.deg_handler_inst.theta_abs[27] ),
    .B(net152),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _3677_ (.A(\cordic_inst.deg_handler_inst.theta_abs[28] ),
    .B(net152),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _3678_ (.A(\cordic_inst.deg_handler_inst.theta_abs[29] ),
    .B(net153),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _3679_ (.A(\cordic_inst.deg_handler_inst.theta_abs[30] ),
    .B(net152),
    .X(_0076_));
 sky130_fd_sc_hd__nand2_1 _3680_ (.A(\cordic_inst.deg_handler_inst.theta_norm[0] ),
    .B(net255),
    .Y(_1816_));
 sky130_fd_sc_hd__xnor2_1 _3681_ (.A(\cordic_inst.deg_handler_inst.theta_norm[1] ),
    .B(_1816_),
    .Y(_0019_));
 sky130_fd_sc_hd__o21ai_1 _3682_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[0] ),
    .A2(\cordic_inst.deg_handler_inst.theta_norm[1] ),
    .B1(net252),
    .Y(_1817_));
 sky130_fd_sc_hd__xnor2_1 _3683_ (.A(\cordic_inst.deg_handler_inst.theta_norm[2] ),
    .B(_1817_),
    .Y(_0030_));
 sky130_fd_sc_hd__o31a_1 _3684_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[0] ),
    .A2(\cordic_inst.deg_handler_inst.theta_norm[1] ),
    .A3(\cordic_inst.deg_handler_inst.theta_norm[2] ),
    .B1(net252),
    .X(_1818_));
 sky130_fd_sc_hd__xor2_1 _3685_ (.A(\cordic_inst.deg_handler_inst.theta_norm[3] ),
    .B(_1818_),
    .X(_0033_));
 sky130_fd_sc_hd__or4_1 _3686_ (.A(\cordic_inst.deg_handler_inst.theta_norm[0] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[1] ),
    .C(\cordic_inst.deg_handler_inst.theta_norm[3] ),
    .D(\cordic_inst.deg_handler_inst.theta_norm[2] ),
    .X(_1819_));
 sky130_fd_sc_hd__nand2_1 _3687_ (.A(net252),
    .B(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__xnor2_1 _3688_ (.A(\cordic_inst.deg_handler_inst.theta_norm[4] ),
    .B(_1820_),
    .Y(_0034_));
 sky130_fd_sc_hd__o21ai_1 _3689_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[4] ),
    .A2(_1819_),
    .B1(net252),
    .Y(_1821_));
 sky130_fd_sc_hd__xnor2_1 _3690_ (.A(\cordic_inst.deg_handler_inst.theta_norm[5] ),
    .B(_1821_),
    .Y(_0035_));
 sky130_fd_sc_hd__or3_1 _3691_ (.A(\cordic_inst.deg_handler_inst.theta_norm[5] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[4] ),
    .C(_1819_),
    .X(_1822_));
 sky130_fd_sc_hd__nand2_1 _3692_ (.A(net252),
    .B(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__xnor2_1 _3693_ (.A(\cordic_inst.deg_handler_inst.theta_norm[6] ),
    .B(_1823_),
    .Y(_0036_));
 sky130_fd_sc_hd__or2_1 _3694_ (.A(\cordic_inst.deg_handler_inst.theta_norm[6] ),
    .B(_1822_),
    .X(_1824_));
 sky130_fd_sc_hd__nand2_1 _3695_ (.A(net252),
    .B(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__xnor2_1 _3696_ (.A(\cordic_inst.deg_handler_inst.theta_norm[7] ),
    .B(_1825_),
    .Y(_0037_));
 sky130_fd_sc_hd__o21ai_1 _3697_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[7] ),
    .A2(_1824_),
    .B1(net252),
    .Y(_1826_));
 sky130_fd_sc_hd__xnor2_1 _3698_ (.A(\cordic_inst.deg_handler_inst.theta_norm[8] ),
    .B(_1826_),
    .Y(_0038_));
 sky130_fd_sc_hd__or3_1 _3699_ (.A(\cordic_inst.deg_handler_inst.theta_norm[8] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[7] ),
    .C(_1824_),
    .X(_1827_));
 sky130_fd_sc_hd__nand2_1 _3700_ (.A(net252),
    .B(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__xnor2_1 _3701_ (.A(\cordic_inst.deg_handler_inst.theta_norm[9] ),
    .B(_1828_),
    .Y(_0039_));
 sky130_fd_sc_hd__or2_1 _3702_ (.A(\cordic_inst.deg_handler_inst.theta_norm[9] ),
    .B(_1827_),
    .X(_1829_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(net252),
    .B(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__xnor2_1 _3704_ (.A(\cordic_inst.deg_handler_inst.theta_norm[10] ),
    .B(_1830_),
    .Y(_0009_));
 sky130_fd_sc_hd__o21ai_1 _3705_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[10] ),
    .A2(_1829_),
    .B1(net252),
    .Y(_1831_));
 sky130_fd_sc_hd__xnor2_1 _3706_ (.A(\cordic_inst.deg_handler_inst.theta_norm[11] ),
    .B(_1831_),
    .Y(_0010_));
 sky130_fd_sc_hd__or3_1 _3707_ (.A(\cordic_inst.deg_handler_inst.theta_norm[11] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[10] ),
    .C(_1829_),
    .X(_1832_));
 sky130_fd_sc_hd__nand2_1 _3708_ (.A(net253),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__xnor2_1 _3709_ (.A(\cordic_inst.deg_handler_inst.theta_norm[12] ),
    .B(_1833_),
    .Y(_0011_));
 sky130_fd_sc_hd__or2_1 _3710_ (.A(\cordic_inst.deg_handler_inst.theta_norm[12] ),
    .B(_1832_),
    .X(_1834_));
 sky130_fd_sc_hd__nand2_1 _3711_ (.A(net253),
    .B(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__xnor2_1 _3712_ (.A(\cordic_inst.deg_handler_inst.theta_norm[13] ),
    .B(_1835_),
    .Y(_0012_));
 sky130_fd_sc_hd__o21ai_1 _3713_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[13] ),
    .A2(_1834_),
    .B1(net253),
    .Y(_1836_));
 sky130_fd_sc_hd__xnor2_1 _3714_ (.A(\cordic_inst.deg_handler_inst.theta_norm[14] ),
    .B(_1836_),
    .Y(_0013_));
 sky130_fd_sc_hd__or3_1 _3715_ (.A(\cordic_inst.deg_handler_inst.theta_norm[14] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[13] ),
    .C(_1834_),
    .X(_1837_));
 sky130_fd_sc_hd__nand2_1 _3716_ (.A(net253),
    .B(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__xnor2_1 _3717_ (.A(\cordic_inst.deg_handler_inst.theta_norm[15] ),
    .B(_1838_),
    .Y(_0014_));
 sky130_fd_sc_hd__or2_1 _3718_ (.A(\cordic_inst.deg_handler_inst.theta_norm[15] ),
    .B(_1837_),
    .X(_1839_));
 sky130_fd_sc_hd__nand2_1 _3719_ (.A(net253),
    .B(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__xnor2_1 _3720_ (.A(\cordic_inst.deg_handler_inst.theta_norm[16] ),
    .B(_1840_),
    .Y(_0015_));
 sky130_fd_sc_hd__o21ai_1 _3721_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[16] ),
    .A2(_1839_),
    .B1(net253),
    .Y(_1841_));
 sky130_fd_sc_hd__xnor2_1 _3722_ (.A(\cordic_inst.deg_handler_inst.theta_norm[17] ),
    .B(_1841_),
    .Y(_0016_));
 sky130_fd_sc_hd__or3_1 _3723_ (.A(\cordic_inst.deg_handler_inst.theta_norm[17] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[16] ),
    .C(_1839_),
    .X(_1842_));
 sky130_fd_sc_hd__nand2_1 _3724_ (.A(net253),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__xnor2_1 _3725_ (.A(\cordic_inst.deg_handler_inst.theta_norm[18] ),
    .B(_1843_),
    .Y(_0017_));
 sky130_fd_sc_hd__or2_1 _3726_ (.A(\cordic_inst.deg_handler_inst.theta_norm[18] ),
    .B(_1842_),
    .X(_1844_));
 sky130_fd_sc_hd__nand2_1 _3727_ (.A(net253),
    .B(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__xnor2_1 _3728_ (.A(\cordic_inst.deg_handler_inst.theta_norm[19] ),
    .B(_1845_),
    .Y(_0018_));
 sky130_fd_sc_hd__o21ai_1 _3729_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[19] ),
    .A2(_1844_),
    .B1(net253),
    .Y(_1846_));
 sky130_fd_sc_hd__xnor2_1 _3730_ (.A(\cordic_inst.deg_handler_inst.theta_norm[20] ),
    .B(_1846_),
    .Y(_0020_));
 sky130_fd_sc_hd__or3_1 _3731_ (.A(\cordic_inst.deg_handler_inst.theta_norm[20] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[19] ),
    .C(_1844_),
    .X(_1847_));
 sky130_fd_sc_hd__nand2_1 _3732_ (.A(net254),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__xnor2_1 _3733_ (.A(\cordic_inst.deg_handler_inst.theta_norm[21] ),
    .B(_1848_),
    .Y(_0021_));
 sky130_fd_sc_hd__or2_1 _3734_ (.A(\cordic_inst.deg_handler_inst.theta_norm[21] ),
    .B(_1847_),
    .X(_1849_));
 sky130_fd_sc_hd__nand2_1 _3735_ (.A(net254),
    .B(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__xnor2_1 _3736_ (.A(\cordic_inst.deg_handler_inst.theta_norm[22] ),
    .B(_1850_),
    .Y(_0022_));
 sky130_fd_sc_hd__o21ai_1 _3737_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[22] ),
    .A2(_1849_),
    .B1(net254),
    .Y(_1851_));
 sky130_fd_sc_hd__xnor2_1 _3738_ (.A(\cordic_inst.deg_handler_inst.theta_norm[23] ),
    .B(_1851_),
    .Y(_0023_));
 sky130_fd_sc_hd__or3_1 _3739_ (.A(\cordic_inst.deg_handler_inst.theta_norm[23] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[22] ),
    .C(_1849_),
    .X(_1852_));
 sky130_fd_sc_hd__nand2_1 _3740_ (.A(net254),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__xnor2_1 _3741_ (.A(\cordic_inst.deg_handler_inst.theta_norm[24] ),
    .B(_1853_),
    .Y(_0024_));
 sky130_fd_sc_hd__or2_1 _3742_ (.A(\cordic_inst.deg_handler_inst.theta_norm[24] ),
    .B(_1852_),
    .X(_1854_));
 sky130_fd_sc_hd__nand2_1 _3743_ (.A(net255),
    .B(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__xnor2_1 _3744_ (.A(\cordic_inst.deg_handler_inst.theta_norm[25] ),
    .B(_1855_),
    .Y(_0025_));
 sky130_fd_sc_hd__o21ai_1 _3745_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[25] ),
    .A2(_1854_),
    .B1(net254),
    .Y(_1856_));
 sky130_fd_sc_hd__xnor2_1 _3746_ (.A(\cordic_inst.deg_handler_inst.theta_norm[26] ),
    .B(_1856_),
    .Y(_0026_));
 sky130_fd_sc_hd__or3_1 _3747_ (.A(\cordic_inst.deg_handler_inst.theta_norm[26] ),
    .B(\cordic_inst.deg_handler_inst.theta_norm[25] ),
    .C(_1854_),
    .X(_1857_));
 sky130_fd_sc_hd__nand2_1 _3748_ (.A(net254),
    .B(_1857_),
    .Y(_1858_));
 sky130_fd_sc_hd__xnor2_1 _3749_ (.A(\cordic_inst.deg_handler_inst.theta_norm[27] ),
    .B(_1858_),
    .Y(_0027_));
 sky130_fd_sc_hd__or2_1 _3750_ (.A(\cordic_inst.deg_handler_inst.theta_norm[27] ),
    .B(_1857_),
    .X(_1859_));
 sky130_fd_sc_hd__nand2_1 _3751_ (.A(net254),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__xnor2_1 _3752_ (.A(\cordic_inst.deg_handler_inst.theta_norm[28] ),
    .B(_1860_),
    .Y(_0028_));
 sky130_fd_sc_hd__nor2_1 _3753_ (.A(\cordic_inst.deg_handler_inst.theta_norm[28] ),
    .B(_1859_),
    .Y(_1861_));
 sky130_fd_sc_hd__o21ai_1 _3754_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[28] ),
    .A2(_1859_),
    .B1(net254),
    .Y(_1862_));
 sky130_fd_sc_hd__xnor2_1 _3755_ (.A(\cordic_inst.deg_handler_inst.theta_norm[29] ),
    .B(_1862_),
    .Y(_0029_));
 sky130_fd_sc_hd__o31a_1 _3756_ (.A1(\cordic_inst.deg_handler_inst.theta_norm[29] ),
    .A2(\cordic_inst.deg_handler_inst.theta_norm[28] ),
    .A3(_1859_),
    .B1(net254),
    .X(_1863_));
 sky130_fd_sc_hd__xor2_1 _3757_ (.A(\cordic_inst.deg_handler_inst.theta_norm[30] ),
    .B(_1863_),
    .X(_0031_));
 sky130_fd_sc_hd__and4bb_1 _3758_ (.A_N(\cordic_inst.deg_handler_inst.theta_norm[30] ),
    .B_N(\cordic_inst.deg_handler_inst.theta_norm[29] ),
    .C(_1861_),
    .D(net254),
    .X(_0032_));
 sky130_fd_sc_hd__or4_1 _3759_ (.A(\axi_controller.reg_input_data[11] ),
    .B(\axi_controller.reg_input_data[10] ),
    .C(\axi_controller.reg_input_data[9] ),
    .D(\axi_controller.reg_input_data[8] ),
    .X(_1864_));
 sky130_fd_sc_hd__or4_1 _3760_ (.A(\axi_controller.reg_input_data[15] ),
    .B(\axi_controller.reg_input_data[14] ),
    .C(\axi_controller.reg_input_data[13] ),
    .D(\axi_controller.reg_input_data[12] ),
    .X(_1865_));
 sky130_fd_sc_hd__or4_1 _3761_ (.A(\axi_controller.reg_input_data[3] ),
    .B(\axi_controller.reg_input_data[2] ),
    .C(\axi_controller.reg_input_data[1] ),
    .D(\axi_controller.reg_input_data[0] ),
    .X(_1866_));
 sky130_fd_sc_hd__or4_1 _3762_ (.A(\axi_controller.reg_input_data[7] ),
    .B(\axi_controller.reg_input_data[6] ),
    .C(\axi_controller.reg_input_data[5] ),
    .D(\axi_controller.reg_input_data[4] ),
    .X(_1867_));
 sky130_fd_sc_hd__or4_1 _3763_ (.A(_1864_),
    .B(_1865_),
    .C(_1866_),
    .D(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__o31a_1 _3764_ (.A1(\axi_controller.reg_input_data[17] ),
    .A2(\axi_controller.reg_input_data[16] ),
    .A3(_1868_),
    .B1(\axi_controller.reg_input_data[18] ),
    .X(_1869_));
 sky130_fd_sc_hd__o211a_1 _3765_ (.A1(\axi_controller.reg_input_data[19] ),
    .A2(_1869_),
    .B1(\axi_controller.reg_input_data[21] ),
    .C1(\axi_controller.reg_input_data[20] ),
    .X(_1870_));
 sky130_fd_sc_hd__o21a_1 _3766_ (.A1(\axi_controller.reg_input_data[22] ),
    .A2(_1870_),
    .B1(\axi_controller.reg_input_data[23] ),
    .X(_1871_));
 sky130_fd_sc_hd__or4_1 _3767_ (.A(\axi_controller.reg_input_data[30] ),
    .B(\axi_controller.reg_input_data[29] ),
    .C(\axi_controller.reg_input_data[28] ),
    .D(\axi_controller.reg_input_data[27] ),
    .X(_1872_));
 sky130_fd_sc_hd__or4_1 _3768_ (.A(\axi_controller.reg_input_data[26] ),
    .B(\axi_controller.reg_input_data[25] ),
    .C(_1871_),
    .D(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__o21bai_2 _3769_ (.A1(\axi_controller.reg_input_data[24] ),
    .A2(_1873_),
    .B1_N(\axi_controller.reg_input_data[31] ),
    .Y(_1874_));
 sky130_fd_sc_hd__a211o_1 _3770_ (.A1(\axi_controller.reg_input_data[19] ),
    .A2(\axi_controller.reg_input_data[18] ),
    .B1(\axi_controller.reg_input_data[21] ),
    .C1(\axi_controller.reg_input_data[20] ),
    .X(_1875_));
 sky130_fd_sc_hd__a21oi_1 _3771_ (.A1(\axi_controller.reg_input_data[22] ),
    .A2(_1875_),
    .B1(\axi_controller.reg_input_data[23] ),
    .Y(_1876_));
 sky130_fd_sc_hd__and4_1 _3772_ (.A(\axi_controller.reg_input_data[28] ),
    .B(\axi_controller.reg_input_data[27] ),
    .C(\axi_controller.reg_input_data[26] ),
    .D(\axi_controller.reg_input_data[25] ),
    .X(_1877_));
 sky130_fd_sc_hd__nand3_1 _3773_ (.A(\axi_controller.reg_input_data[30] ),
    .B(\axi_controller.reg_input_data[29] ),
    .C(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__or3b_1 _3774_ (.A(_1876_),
    .B(_1878_),
    .C_N(\axi_controller.reg_input_data[24] ),
    .X(_1879_));
 sky130_fd_sc_hd__nand2_2 _3775_ (.A(\axi_controller.reg_input_data[31] ),
    .B(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__nand2_1 _3776_ (.A(_1874_),
    .B(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hd__xor2_1 _3777_ (.A(\axi_controller.reg_input_data[19] ),
    .B(_1881_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(_1874_),
    .A1(_1880_),
    .S(\axi_controller.reg_input_data[19] ),
    .X(_1882_));
 sky130_fd_sc_hd__xnor2_1 _3779_ (.A(\axi_controller.reg_input_data[20] ),
    .B(_1882_),
    .Y(_0041_));
 sky130_fd_sc_hd__and2_1 _3780_ (.A(\axi_controller.reg_input_data[20] ),
    .B(\axi_controller.reg_input_data[19] ),
    .X(_1883_));
 sky130_fd_sc_hd__nor3_1 _3781_ (.A(\axi_controller.reg_input_data[21] ),
    .B(_1880_),
    .C(_1883_),
    .Y(_1884_));
 sky130_fd_sc_hd__o21a_1 _3782_ (.A1(_1880_),
    .A2(_1883_),
    .B1(\axi_controller.reg_input_data[21] ),
    .X(_1885_));
 sky130_fd_sc_hd__o21ba_1 _3783_ (.A1(\axi_controller.reg_input_data[20] ),
    .A2(\axi_controller.reg_input_data[19] ),
    .B1_N(_1874_),
    .X(_1886_));
 sky130_fd_sc_hd__nand2_1 _3784_ (.A(\axi_controller.reg_input_data[21] ),
    .B(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__or3_1 _3785_ (.A(_1884_),
    .B(_1885_),
    .C(_1886_),
    .X(_1888_));
 sky130_fd_sc_hd__and2_1 _3786_ (.A(_1887_),
    .B(_1888_),
    .X(_0042_));
 sky130_fd_sc_hd__o31a_1 _3787_ (.A1(\axi_controller.reg_input_data[21] ),
    .A2(_1880_),
    .A3(_1883_),
    .B1(_1887_),
    .X(_1889_));
 sky130_fd_sc_hd__xnor2_1 _3788_ (.A(\axi_controller.reg_input_data[22] ),
    .B(_1889_),
    .Y(_0043_));
 sky130_fd_sc_hd__o211a_1 _3789_ (.A1(\axi_controller.reg_input_data[20] ),
    .A2(\axi_controller.reg_input_data[19] ),
    .B1(\axi_controller.reg_input_data[22] ),
    .C1(\axi_controller.reg_input_data[21] ),
    .X(_1890_));
 sky130_fd_sc_hd__nor2_1 _3790_ (.A(_1874_),
    .B(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__or3_1 _3791_ (.A(\axi_controller.reg_input_data[22] ),
    .B(\axi_controller.reg_input_data[21] ),
    .C(_1883_),
    .X(_1892_));
 sky130_fd_sc_hd__a21oi_1 _3792_ (.A1(\axi_controller.reg_input_data[23] ),
    .A2(_1892_),
    .B1(_1880_),
    .Y(_1893_));
 sky130_fd_sc_hd__o21a_1 _3793_ (.A1(\axi_controller.reg_input_data[23] ),
    .A2(_1892_),
    .B1(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__a21oi_1 _3794_ (.A1(\axi_controller.reg_input_data[23] ),
    .A2(_1880_),
    .B1(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__xnor2_1 _3795_ (.A(_1891_),
    .B(_1895_),
    .Y(_0044_));
 sky130_fd_sc_hd__o21ba_1 _3796_ (.A1(\axi_controller.reg_input_data[23] ),
    .A2(_1890_),
    .B1_N(_1874_),
    .X(_1896_));
 sky130_fd_sc_hd__xnor2_1 _3797_ (.A(\axi_controller.reg_input_data[24] ),
    .B(_1893_),
    .Y(_1897_));
 sky130_fd_sc_hd__xnor2_1 _3798_ (.A(_1896_),
    .B(_1897_),
    .Y(_0045_));
 sky130_fd_sc_hd__a21oi_1 _3799_ (.A1(\axi_controller.reg_input_data[23] ),
    .A2(_1892_),
    .B1(\axi_controller.reg_input_data[24] ),
    .Y(_1898_));
 sky130_fd_sc_hd__or2_1 _3800_ (.A(_1880_),
    .B(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__inv_2 _3801_ (.A(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__xnor2_1 _3802_ (.A(\axi_controller.reg_input_data[25] ),
    .B(_1899_),
    .Y(_1901_));
 sky130_fd_sc_hd__o21a_1 _3803_ (.A1(\axi_controller.reg_input_data[23] ),
    .A2(_1890_),
    .B1(\axi_controller.reg_input_data[24] ),
    .X(_1902_));
 sky130_fd_sc_hd__or2_1 _3804_ (.A(_1874_),
    .B(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__xnor2_1 _3805_ (.A(_1901_),
    .B(_1903_),
    .Y(_0046_));
 sky130_fd_sc_hd__mux2_1 _3806_ (.A0(_1903_),
    .A1(_1899_),
    .S(\axi_controller.reg_input_data[25] ),
    .X(_1904_));
 sky130_fd_sc_hd__xnor2_1 _3807_ (.A(\axi_controller.reg_input_data[26] ),
    .B(_1904_),
    .Y(_0047_));
 sky130_fd_sc_hd__and3_1 _3808_ (.A(\axi_controller.reg_input_data[26] ),
    .B(\axi_controller.reg_input_data[25] ),
    .C(_1900_),
    .X(_1905_));
 sky130_fd_sc_hd__inv_2 _3809_ (.A(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__xor2_1 _3810_ (.A(\axi_controller.reg_input_data[27] ),
    .B(_1905_),
    .X(_1907_));
 sky130_fd_sc_hd__or3_1 _3811_ (.A(\axi_controller.reg_input_data[26] ),
    .B(\axi_controller.reg_input_data[25] ),
    .C(_1903_),
    .X(_1908_));
 sky130_fd_sc_hd__xnor2_1 _3812_ (.A(_1907_),
    .B(_1908_),
    .Y(_0048_));
 sky130_fd_sc_hd__mux2_1 _3813_ (.A0(_1908_),
    .A1(_1906_),
    .S(\axi_controller.reg_input_data[27] ),
    .X(_1909_));
 sky130_fd_sc_hd__xnor2_1 _3814_ (.A(\axi_controller.reg_input_data[28] ),
    .B(_1909_),
    .Y(_0049_));
 sky130_fd_sc_hd__and2_1 _3815_ (.A(_1877_),
    .B(_1900_),
    .X(_1910_));
 sky130_fd_sc_hd__xnor2_1 _3816_ (.A(\axi_controller.reg_input_data[29] ),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__nor3_1 _3817_ (.A(\axi_controller.reg_input_data[28] ),
    .B(\axi_controller.reg_input_data[27] ),
    .C(_1908_),
    .Y(_1912_));
 sky130_fd_sc_hd__xnor2_1 _3818_ (.A(_1911_),
    .B(_1912_),
    .Y(_0050_));
 sky130_fd_sc_hd__mux2_1 _3819_ (.A0(_1912_),
    .A1(_1910_),
    .S(\axi_controller.reg_input_data[29] ),
    .X(_1913_));
 sky130_fd_sc_hd__xor2_1 _3820_ (.A(\axi_controller.reg_input_data[30] ),
    .B(_1913_),
    .X(_0051_));
 sky130_fd_sc_hd__nor2_1 _3821_ (.A(_1878_),
    .B(_1898_),
    .Y(_1914_));
 sky130_fd_sc_hd__xnor2_1 _3822_ (.A(_1880_),
    .B(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__or4_1 _3823_ (.A(\axi_controller.reg_input_data[26] ),
    .B(\axi_controller.reg_input_data[25] ),
    .C(_1872_),
    .D(_1903_),
    .X(_1916_));
 sky130_fd_sc_hd__a21bo_1 _3824_ (.A1(_1874_),
    .A2(_1915_),
    .B1_N(_1916_),
    .X(_0052_));
 sky130_fd_sc_hd__o21ba_1 _3825_ (.A1(\cordic_inst.cordic_inst.start ),
    .A2(\cordic_inst.cordic_inst.state[1] ),
    .B1_N(\cordic_inst.cordic_inst.state[0] ),
    .X(_1917_));
 sky130_fd_sc_hd__o21a_1 _3826_ (.A1(net274),
    .A2(_0614_),
    .B1(_1917_),
    .X(\cordic_inst.cordic_inst.next_state[0] ));
 sky130_fd_sc_hd__nand2b_1 _3827_ (.A_N(\axi_controller.reg_done_flag ),
    .B(\axi_controller.start_pulse_reg ),
    .Y(_1918_));
 sky130_fd_sc_hd__nor2_1 _3828_ (.A(_0618_),
    .B(_1918_),
    .Y(_0000_));
 sky130_fd_sc_hd__and2b_1 _3829_ (.A_N(\cordic_inst.sign_handler_inst.done_d ),
    .B(\cordic_inst.cordic_inst.done ),
    .X(\cordic_inst.sign_handler_inst.done_pulse ));
 sky130_fd_sc_hd__nand2b_1 _3830_ (.A_N(\cordic_inst.done_d ),
    .B(\axi_controller.done ),
    .Y(_1919_));
 sky130_fd_sc_hd__a21o_1 _3831_ (.A1(\cordic_inst.state[1] ),
    .A2(_1919_),
    .B1(\cordic_inst.state[2] ),
    .X(_0007_));
 sky130_fd_sc_hd__a2bb2o_1 _3832_ (.A1_N(_0620_),
    .A2_N(_1919_),
    .B1(_1918_),
    .B2(\cordic_inst.state[0] ),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _3833_ (.A(net111),
    .B(net69),
    .Y(_1920_));
 sky130_fd_sc_hd__a31o_1 _3834_ (.A1(net111),
    .A2(\axi_controller.state[2] ),
    .A3(net69),
    .B1(_0621_),
    .X(_1921_));
 sky130_fd_sc_hd__or2_1 _3835_ (.A(_0610_),
    .B(net68),
    .X(_1922_));
 sky130_fd_sc_hd__nor2_1 _3836_ (.A(net68),
    .B(net35),
    .Y(_1923_));
 sky130_fd_sc_hd__nor2_1 _3837_ (.A(net35),
    .B(_1922_),
    .Y(_1924_));
 sky130_fd_sc_hd__a31o_1 _3838_ (.A1(net145),
    .A2(\axi_controller.state[1] ),
    .A3(net70),
    .B1(_1921_),
    .X(_1925_));
 sky130_fd_sc_hd__or2_1 _3839_ (.A(_1924_),
    .B(_1925_),
    .X(_0001_));
 sky130_fd_sc_hd__and4b_1 _3840_ (.A_N(net68),
    .B(net35),
    .C(\axi_controller.state[0] ),
    .D(net349),
    .X(_1926_));
 sky130_fd_sc_hd__nand2_1 _3841_ (.A(\axi_controller.state[1] ),
    .B(net349),
    .Y(_1927_));
 sky130_fd_sc_hd__a21oi_1 _3842_ (.A1(net145),
    .A2(net70),
    .B1(net194),
    .Y(_1928_));
 sky130_fd_sc_hd__or2_1 _3843_ (.A(net199),
    .B(_1928_),
    .X(_0002_));
 sky130_fd_sc_hd__and4_1 _3844_ (.A(\axi_controller.state[0] ),
    .B(net349),
    .C(net68),
    .D(_0622_),
    .X(_1929_));
 sky130_fd_sc_hd__a31o_1 _3845_ (.A1(net349),
    .A2(_0622_),
    .A3(\axi_controller.state[3] ),
    .B1(net188),
    .X(_0004_));
 sky130_fd_sc_hd__and3_1 _3846_ (.A(net349),
    .B(net107),
    .C(\axi_controller.state[3] ),
    .X(_1930_));
 sky130_fd_sc_hd__a32o_1 _3847_ (.A1(\axi_controller.state[0] ),
    .A2(net68),
    .A3(net107),
    .B1(_1920_),
    .B2(\axi_controller.state[2] ),
    .X(_1931_));
 sky130_fd_sc_hd__a21o_1 _3848_ (.A1(net349),
    .A2(_1931_),
    .B1(_1930_),
    .X(_0003_));
 sky130_fd_sc_hd__nand3b_1 _3849_ (.A_N(net63),
    .B(net62),
    .C(net61),
    .Y(_1932_));
 sky130_fd_sc_hd__or4_1 _3850_ (.A(net58),
    .B(net65),
    .C(net64),
    .D(net67),
    .X(_1933_));
 sky130_fd_sc_hd__or4_1 _3851_ (.A(net66),
    .B(net38),
    .C(net37),
    .D(net40),
    .X(_1934_));
 sky130_fd_sc_hd__or4_1 _3852_ (.A(net49),
    .B(net48),
    .C(net51),
    .D(net50),
    .X(_1935_));
 sky130_fd_sc_hd__or4_1 _3853_ (.A(net44),
    .B(net43),
    .C(net46),
    .D(net45),
    .X(_1936_));
 sky130_fd_sc_hd__or4_1 _3854_ (.A(net53),
    .B(net52),
    .C(net55),
    .D(net54),
    .X(_1937_));
 sky130_fd_sc_hd__and4_1 _3855_ (.A(net56),
    .B(net57),
    .C(net59),
    .D(net60),
    .X(_1938_));
 sky130_fd_sc_hd__or4b_1 _3856_ (.A(_1935_),
    .B(_1936_),
    .C(_1937_),
    .D_N(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__or4_1 _3857_ (.A(net39),
    .B(net42),
    .C(net41),
    .D(_1934_),
    .X(_1940_));
 sky130_fd_sc_hd__or4_1 _3858_ (.A(net47),
    .B(net36),
    .C(_1933_),
    .D(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__o311a_1 _3859_ (.A1(_1932_),
    .A2(_1939_),
    .A3(_1941_),
    .B1(net107),
    .C1(net68),
    .X(_1942_));
 sky130_fd_sc_hd__or2_1 _3860_ (.A(\axi_controller.state[0] ),
    .B(\axi_controller.state[3] ),
    .X(_1943_));
 sky130_fd_sc_hd__or4_1 _3861_ (.A(\axi_controller.write_addr_reg[20] ),
    .B(\axi_controller.write_addr_reg[23] ),
    .C(\axi_controller.write_addr_reg[22] ),
    .D(\axi_controller.write_addr_reg[25] ),
    .X(_1944_));
 sky130_fd_sc_hd__or4_1 _3862_ (.A(\axi_controller.write_addr_reg[16] ),
    .B(\axi_controller.write_addr_reg[19] ),
    .C(\axi_controller.write_addr_reg[18] ),
    .D(\axi_controller.write_addr_reg[21] ),
    .X(_1945_));
 sky130_fd_sc_hd__nand3_1 _3863_ (.A(\axi_controller.write_addr_reg[29] ),
    .B(\axi_controller.write_addr_reg[30] ),
    .C(\axi_controller.write_addr_reg[31] ),
    .Y(_1946_));
 sky130_fd_sc_hd__or4b_1 _3864_ (.A(\axi_controller.write_addr_reg[24] ),
    .B(\axi_controller.write_addr_reg[27] ),
    .C(\axi_controller.write_addr_reg[26] ),
    .D_N(\axi_controller.write_addr_reg[28] ),
    .X(_1947_));
 sky130_fd_sc_hd__or4_1 _3865_ (.A(_1944_),
    .B(_1945_),
    .C(_1946_),
    .D(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__or4_1 _3866_ (.A(\axi_controller.write_addr_reg[2] ),
    .B(\axi_controller.write_addr_reg[7] ),
    .C(\axi_controller.write_addr_reg[6] ),
    .D(\axi_controller.write_addr_reg[9] ),
    .X(_1949_));
 sky130_fd_sc_hd__or3_1 _3867_ (.A(\axi_controller.write_addr_reg[1] ),
    .B(\axi_controller.write_addr_reg[0] ),
    .C(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__or4_1 _3868_ (.A(\axi_controller.write_addr_reg[8] ),
    .B(\axi_controller.write_addr_reg[11] ),
    .C(\axi_controller.write_addr_reg[10] ),
    .D(\axi_controller.write_addr_reg[13] ),
    .X(_1951_));
 sky130_fd_sc_hd__or4_1 _3869_ (.A(\axi_controller.write_addr_reg[12] ),
    .B(\axi_controller.write_addr_reg[15] ),
    .C(\axi_controller.write_addr_reg[14] ),
    .D(\axi_controller.write_addr_reg[17] ),
    .X(_1952_));
 sky130_fd_sc_hd__or4_1 _3870_ (.A(_1948_),
    .B(_1950_),
    .C(_1951_),
    .D(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__or4_1 _3871_ (.A(\axi_controller.write_addr_reg[12] ),
    .B(\axi_controller.write_addr_reg[15] ),
    .C(\axi_controller.write_addr_reg[14] ),
    .D(_1951_),
    .X(_1954_));
 sky130_fd_sc_hd__or4_1 _3872_ (.A(\axi_controller.write_addr_reg[21] ),
    .B(\axi_controller.write_addr_reg[20] ),
    .C(\axi_controller.write_addr_reg[23] ),
    .D(\axi_controller.write_addr_reg[22] ),
    .X(_1955_));
 sky130_fd_sc_hd__nand4_1 _3873_ (.A(\axi_controller.write_addr_reg[28] ),
    .B(\axi_controller.write_addr_reg[29] ),
    .C(\axi_controller.write_addr_reg[30] ),
    .D(\axi_controller.write_addr_reg[31] ),
    .Y(_1956_));
 sky130_fd_sc_hd__or4_1 _3874_ (.A(\axi_controller.write_addr_reg[25] ),
    .B(\axi_controller.write_addr_reg[24] ),
    .C(\axi_controller.write_addr_reg[27] ),
    .D(\axi_controller.write_addr_reg[26] ),
    .X(_1957_));
 sky130_fd_sc_hd__or4_1 _3875_ (.A(\axi_controller.write_addr_reg[17] ),
    .B(\axi_controller.write_addr_reg[16] ),
    .C(\axi_controller.write_addr_reg[19] ),
    .D(\axi_controller.write_addr_reg[18] ),
    .X(_1958_));
 sky130_fd_sc_hd__or4_1 _3876_ (.A(_1955_),
    .B(_1956_),
    .C(_1957_),
    .D(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__or3b_1 _3877_ (.A(\axi_controller.write_addr_reg[5] ),
    .B(_1959_),
    .C_N(\axi_controller.write_addr_reg[3] ),
    .X(_1960_));
 sky130_fd_sc_hd__or4_1 _3878_ (.A(_0623_),
    .B(_1950_),
    .C(_1954_),
    .D(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__a32o_1 _3879_ (.A1(net107),
    .A2(\axi_controller.state[3] ),
    .A3(_1961_),
    .B1(_1942_),
    .B2(\axi_controller.state[0] ),
    .X(_1962_));
 sky130_fd_sc_hd__and4bb_4 _3880_ (.A_N(_0622_),
    .B_N(_1962_),
    .C(_1943_),
    .D(_1922_),
    .X(_1963_));
 sky130_fd_sc_hd__and2_1 _3881_ (.A(net104),
    .B(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__nand2_2 _3882_ (.A(net104),
    .B(_1963_),
    .Y(_1965_));
 sky130_fd_sc_hd__or2_1 _3883_ (.A(\axi_controller.reg_input_data[8] ),
    .B(_1964_),
    .X(_1966_));
 sky130_fd_sc_hd__o211a_1 _3884_ (.A1(net101),
    .A2(_1965_),
    .B1(_1966_),
    .C1(net346),
    .X(_0258_));
 sky130_fd_sc_hd__or2_1 _3885_ (.A(\axi_controller.reg_input_data[9] ),
    .B(_1964_),
    .X(_1967_));
 sky130_fd_sc_hd__o211a_1 _3886_ (.A1(net102),
    .A2(_1965_),
    .B1(_1967_),
    .C1(net347),
    .X(_0259_));
 sky130_fd_sc_hd__or2_1 _3887_ (.A(\axi_controller.reg_input_data[10] ),
    .B(_1964_),
    .X(_1968_));
 sky130_fd_sc_hd__o211a_1 _3888_ (.A1(net72),
    .A2(_1965_),
    .B1(_1968_),
    .C1(net346),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _3889_ (.A(\axi_controller.reg_input_data[11] ),
    .B(_1964_),
    .X(_1969_));
 sky130_fd_sc_hd__o211a_1 _3890_ (.A1(net73),
    .A2(_1965_),
    .B1(_1969_),
    .C1(net347),
    .X(_0261_));
 sky130_fd_sc_hd__or2_1 _3891_ (.A(\axi_controller.reg_input_data[12] ),
    .B(_1964_),
    .X(_1970_));
 sky130_fd_sc_hd__o211a_1 _3892_ (.A1(net74),
    .A2(_1965_),
    .B1(_1970_),
    .C1(net347),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _3893_ (.A(\axi_controller.reg_input_data[13] ),
    .B(_1964_),
    .X(_1971_));
 sky130_fd_sc_hd__o211a_1 _3894_ (.A1(net75),
    .A2(_1965_),
    .B1(_1971_),
    .C1(net346),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _3895_ (.A(\axi_controller.reg_input_data[14] ),
    .B(_1964_),
    .X(_1972_));
 sky130_fd_sc_hd__o211a_1 _3896_ (.A1(net76),
    .A2(_1965_),
    .B1(_1972_),
    .C1(net347),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _3897_ (.A(\axi_controller.reg_input_data[15] ),
    .B(_1964_),
    .X(_1973_));
 sky130_fd_sc_hd__o211a_1 _3898_ (.A1(net77),
    .A2(_1965_),
    .B1(_1973_),
    .C1(net347),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3899_ (.A0(\axi_controller.read_addr_reg[0] ),
    .A1(net2),
    .S(net197),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _3900_ (.A0(\axi_controller.read_addr_reg[1] ),
    .A1(net13),
    .S(net197),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3901_ (.A0(\axi_controller.read_addr_reg[2] ),
    .A1(net24),
    .S(net195),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3902_ (.A0(\axi_controller.read_addr_reg[3] ),
    .A1(net27),
    .S(net197),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3903_ (.A0(\axi_controller.read_addr_reg[4] ),
    .A1(net28),
    .S(net198),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _3904_ (.A0(\axi_controller.read_addr_reg[5] ),
    .A1(net29),
    .S(net198),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3905_ (.A0(\axi_controller.read_addr_reg[6] ),
    .A1(net30),
    .S(net198),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(\axi_controller.read_addr_reg[7] ),
    .A1(net31),
    .S(net198),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3907_ (.A0(\axi_controller.read_addr_reg[8] ),
    .A1(net32),
    .S(net195),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _3908_ (.A0(\axi_controller.read_addr_reg[9] ),
    .A1(net33),
    .S(net195),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3909_ (.A0(\axi_controller.read_addr_reg[10] ),
    .A1(net3),
    .S(net196),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _3910_ (.A0(\axi_controller.read_addr_reg[11] ),
    .A1(net4),
    .S(net195),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3911_ (.A0(\axi_controller.read_addr_reg[12] ),
    .A1(net5),
    .S(net198),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(\axi_controller.read_addr_reg[13] ),
    .A1(net6),
    .S(net195),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3913_ (.A0(\axi_controller.read_addr_reg[14] ),
    .A1(net7),
    .S(net196),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(\axi_controller.read_addr_reg[15] ),
    .A1(net8),
    .S(net196),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3915_ (.A0(\axi_controller.read_addr_reg[16] ),
    .A1(net9),
    .S(net197),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _3916_ (.A0(\axi_controller.read_addr_reg[17] ),
    .A1(net10),
    .S(net197),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(\axi_controller.read_addr_reg[18] ),
    .A1(net11),
    .S(net196),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3918_ (.A0(\axi_controller.read_addr_reg[19] ),
    .A1(net12),
    .S(net197),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3919_ (.A0(\axi_controller.read_addr_reg[20] ),
    .A1(net14),
    .S(net196),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(\axi_controller.read_addr_reg[21] ),
    .A1(net15),
    .S(net196),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3921_ (.A0(\axi_controller.read_addr_reg[22] ),
    .A1(net16),
    .S(net196),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _3922_ (.A0(\axi_controller.read_addr_reg[23] ),
    .A1(net17),
    .S(net197),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3923_ (.A0(\axi_controller.read_addr_reg[24] ),
    .A1(net18),
    .S(net195),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _3924_ (.A0(\axi_controller.read_addr_reg[25] ),
    .A1(net19),
    .S(net197),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _3925_ (.A0(\axi_controller.read_addr_reg[26] ),
    .A1(net20),
    .S(net197),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _3926_ (.A0(\axi_controller.read_addr_reg[27] ),
    .A1(net21),
    .S(net195),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3927_ (.A0(\axi_controller.read_addr_reg[28] ),
    .A1(net22),
    .S(net197),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _3928_ (.A0(\axi_controller.read_addr_reg[29] ),
    .A1(net23),
    .S(net195),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3929_ (.A0(\axi_controller.read_addr_reg[30] ),
    .A1(net25),
    .S(net195),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _3930_ (.A0(\axi_controller.read_addr_reg[31] ),
    .A1(net26),
    .S(net195),
    .X(_0297_));
 sky130_fd_sc_hd__or4_1 _3931_ (.A(\axi_controller.read_addr_reg[13] ),
    .B(\axi_controller.read_addr_reg[12] ),
    .C(\axi_controller.read_addr_reg[15] ),
    .D(\axi_controller.read_addr_reg[14] ),
    .X(_1974_));
 sky130_fd_sc_hd__or4_1 _3932_ (.A(\axi_controller.read_addr_reg[9] ),
    .B(\axi_controller.read_addr_reg[8] ),
    .C(\axi_controller.read_addr_reg[11] ),
    .D(\axi_controller.read_addr_reg[10] ),
    .X(_1975_));
 sky130_fd_sc_hd__nor2_1 _3933_ (.A(_1974_),
    .B(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__nor4_1 _3934_ (.A(\axi_controller.read_addr_reg[1] ),
    .B(\axi_controller.read_addr_reg[0] ),
    .C(\axi_controller.read_addr_reg[7] ),
    .D(\axi_controller.read_addr_reg[6] ),
    .Y(_1977_));
 sky130_fd_sc_hd__and4bb_1 _3935_ (.A_N(\axi_controller.read_addr_reg[3] ),
    .B_N(\axi_controller.read_addr_reg[4] ),
    .C(\axi_controller.read_addr_reg[5] ),
    .D(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__nand2_1 _3936_ (.A(_1976_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__or4_1 _3937_ (.A(\axi_controller.read_addr_reg[16] ),
    .B(\axi_controller.read_addr_reg[19] ),
    .C(\axi_controller.read_addr_reg[18] ),
    .D(\axi_controller.read_addr_reg[21] ),
    .X(_1980_));
 sky130_fd_sc_hd__or3b_1 _3938_ (.A(\axi_controller.read_addr_reg[17] ),
    .B(_1980_),
    .C_N(\axi_controller.read_addr_reg[2] ),
    .X(_1981_));
 sky130_fd_sc_hd__nand2_1 _3939_ (.A(\axi_controller.read_addr_reg[29] ),
    .B(\axi_controller.read_addr_reg[30] ),
    .Y(_1982_));
 sky130_fd_sc_hd__or2_1 _3940_ (.A(_0625_),
    .B(_1982_),
    .X(_1983_));
 sky130_fd_sc_hd__or4b_1 _3941_ (.A(\axi_controller.read_addr_reg[24] ),
    .B(\axi_controller.read_addr_reg[27] ),
    .C(\axi_controller.read_addr_reg[26] ),
    .D_N(\axi_controller.read_addr_reg[28] ),
    .X(_1984_));
 sky130_fd_sc_hd__or4_1 _3942_ (.A(\axi_controller.read_addr_reg[20] ),
    .B(\axi_controller.read_addr_reg[23] ),
    .C(\axi_controller.read_addr_reg[22] ),
    .D(\axi_controller.read_addr_reg[25] ),
    .X(_1985_));
 sky130_fd_sc_hd__or4_1 _3943_ (.A(\axi_controller.read_addr_reg[20] ),
    .B(\axi_controller.read_addr_reg[23] ),
    .C(\axi_controller.read_addr_reg[22] ),
    .D(_1984_),
    .X(_1986_));
 sky130_fd_sc_hd__nor4_1 _3944_ (.A(\axi_controller.read_addr_reg[25] ),
    .B(_1981_),
    .C(_1983_),
    .D(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__or4_1 _3945_ (.A(_0625_),
    .B(_1982_),
    .C(_1984_),
    .D(_1985_),
    .X(_1988_));
 sky130_fd_sc_hd__or4b_1 _3946_ (.A(\axi_controller.read_addr_reg[17] ),
    .B(_1980_),
    .C(_1988_),
    .D_N(\axi_controller.read_addr_reg[2] ),
    .X(_1989_));
 sky130_fd_sc_hd__nor2_1 _3947_ (.A(_1979_),
    .B(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__nand2_1 _3948_ (.A(net70),
    .B(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__o21a_1 _3949_ (.A1(_0619_),
    .A2(_1991_),
    .B1(\axi_controller.reg_done_flag ),
    .X(_1992_));
 sky130_fd_sc_hd__o2111a_1 _3950_ (.A1(\axi_controller.done ),
    .A2(_1992_),
    .B1(net349),
    .C1(_0085_),
    .D1(_1918_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _3951_ (.A0(\axi_controller.write_addr_reg[0] ),
    .A1(net36),
    .S(net187),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(\axi_controller.write_addr_reg[1] ),
    .A1(net47),
    .S(net187),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _3953_ (.A0(\axi_controller.write_addr_reg[2] ),
    .A1(net58),
    .S(net187),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3954_ (.A0(\axi_controller.write_addr_reg[3] ),
    .A1(net61),
    .S(net190),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _3955_ (.A0(\axi_controller.write_addr_reg[4] ),
    .A1(net62),
    .S(net188),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3956_ (.A0(\axi_controller.write_addr_reg[5] ),
    .A1(net63),
    .S(net188),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _3957_ (.A0(\axi_controller.write_addr_reg[6] ),
    .A1(net64),
    .S(net187),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(\axi_controller.write_addr_reg[7] ),
    .A1(net65),
    .S(net187),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _3959_ (.A0(\axi_controller.write_addr_reg[8] ),
    .A1(net66),
    .S(net187),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _3960_ (.A0(\axi_controller.write_addr_reg[9] ),
    .A1(net67),
    .S(net187),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _3961_ (.A0(\axi_controller.write_addr_reg[10] ),
    .A1(net37),
    .S(net187),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3962_ (.A0(\axi_controller.write_addr_reg[11] ),
    .A1(net38),
    .S(net187),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _3963_ (.A0(\axi_controller.write_addr_reg[12] ),
    .A1(net39),
    .S(net188),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(\axi_controller.write_addr_reg[13] ),
    .A1(net40),
    .S(net187),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _3965_ (.A0(\axi_controller.write_addr_reg[14] ),
    .A1(net41),
    .S(net188),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3966_ (.A0(\axi_controller.write_addr_reg[15] ),
    .A1(net42),
    .S(net188),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _3967_ (.A0(\axi_controller.write_addr_reg[16] ),
    .A1(net43),
    .S(net190),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(\axi_controller.write_addr_reg[17] ),
    .A1(net44),
    .S(net190),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _3969_ (.A0(\axi_controller.write_addr_reg[18] ),
    .A1(net45),
    .S(net190),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3970_ (.A0(\axi_controller.write_addr_reg[19] ),
    .A1(net46),
    .S(net190),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _3971_ (.A0(\axi_controller.write_addr_reg[20] ),
    .A1(net48),
    .S(net189),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3972_ (.A0(\axi_controller.write_addr_reg[21] ),
    .A1(net49),
    .S(net190),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3973_ (.A0(\axi_controller.write_addr_reg[22] ),
    .A1(net50),
    .S(net189),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(\axi_controller.write_addr_reg[23] ),
    .A1(net51),
    .S(net189),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _3975_ (.A0(\axi_controller.write_addr_reg[24] ),
    .A1(net52),
    .S(net190),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3976_ (.A0(\axi_controller.write_addr_reg[25] ),
    .A1(net53),
    .S(net189),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(\axi_controller.write_addr_reg[26] ),
    .A1(net54),
    .S(net189),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3978_ (.A0(\axi_controller.write_addr_reg[27] ),
    .A1(net55),
    .S(net189),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(\axi_controller.write_addr_reg[28] ),
    .A1(net56),
    .S(net189),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(\axi_controller.write_addr_reg[29] ),
    .A1(net57),
    .S(net189),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3981_ (.A0(\axi_controller.write_addr_reg[30] ),
    .A1(net59),
    .S(net189),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(\axi_controller.write_addr_reg[31] ),
    .A1(net60),
    .S(net189),
    .X(_0330_));
 sky130_fd_sc_hd__or4b_1 _3983_ (.A(\axi_controller.write_addr_reg[3] ),
    .B(\axi_controller.write_addr_reg[4] ),
    .C(_1953_),
    .D_N(\axi_controller.write_addr_reg[5] ),
    .X(_1993_));
 sky130_fd_sc_hd__inv_2 _3984_ (.A(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__nor2_1 _3985_ (.A(_0624_),
    .B(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__nand4_1 _3986_ (.A(net107),
    .B(net103),
    .C(_1922_),
    .D(_1943_),
    .Y(_1996_));
 sky130_fd_sc_hd__or3b_1 _3987_ (.A(net61),
    .B(net62),
    .C_N(net63),
    .X(_1997_));
 sky130_fd_sc_hd__or3_1 _3988_ (.A(_1939_),
    .B(_1941_),
    .C(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__a211o_1 _3989_ (.A1(\axi_controller.state[0] ),
    .A2(_1998_),
    .B1(_1996_),
    .C1(_1995_),
    .X(_1999_));
 sky130_fd_sc_hd__mux2_1 _3990_ (.A0(net71),
    .A1(net319),
    .S(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__and2_1 _3991_ (.A(net350),
    .B(_2000_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3992_ (.A0(net93),
    .A1(net313),
    .S(_1999_),
    .X(_2001_));
 sky130_fd_sc_hd__and2_1 _3993_ (.A(net350),
    .B(_2001_),
    .X(_0332_));
 sky130_fd_sc_hd__a41o_1 _3994_ (.A1(_0610_),
    .A2(net145),
    .A3(_0619_),
    .A4(net350),
    .B1(_1928_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _3995_ (.A1(net107),
    .A2(_0624_),
    .B1(_1943_),
    .Y(_2002_));
 sky130_fd_sc_hd__a31o_1 _3996_ (.A1(_0624_),
    .A2(_1942_),
    .A3(_1998_),
    .B1(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__a21oi_1 _3997_ (.A1(_1961_),
    .A2(_1995_),
    .B1(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__a211oi_1 _3998_ (.A1(_0611_),
    .A2(_2002_),
    .B1(_2004_),
    .C1(_0621_),
    .Y(_0334_));
 sky130_fd_sc_hd__a21oi_1 _3999_ (.A1(net108),
    .A2(_0610_),
    .B1(_1924_),
    .Y(_2005_));
 sky130_fd_sc_hd__nor2_1 _4000_ (.A(_0621_),
    .B(_2005_),
    .Y(_0335_));
 sky130_fd_sc_hd__a21oi_1 _4001_ (.A1(net111),
    .A2(_0610_),
    .B1(\axi_controller.state[2] ),
    .Y(_2006_));
 sky130_fd_sc_hd__nor2_1 _4002_ (.A(_1921_),
    .B(_2006_),
    .Y(_0336_));
 sky130_fd_sc_hd__a22o_1 _4003_ (.A1(net68),
    .A2(_0622_),
    .B1(_0624_),
    .B2(_1923_),
    .X(_2007_));
 sky130_fd_sc_hd__o221a_1 _4004_ (.A1(net146),
    .A2(_1943_),
    .B1(_2002_),
    .B2(_2007_),
    .C1(net350),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _4005_ (.A(net106),
    .B(_1963_),
    .X(_2008_));
 sky130_fd_sc_hd__nand2_2 _4006_ (.A(net106),
    .B(_1963_),
    .Y(_2009_));
 sky130_fd_sc_hd__or2_1 _4007_ (.A(\axi_controller.reg_input_data[24] ),
    .B(_2008_),
    .X(_2010_));
 sky130_fd_sc_hd__o211a_1 _4008_ (.A1(net87),
    .A2(_2009_),
    .B1(_2010_),
    .C1(net346),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _4009_ (.A(\axi_controller.reg_input_data[25] ),
    .B(_2008_),
    .X(_2011_));
 sky130_fd_sc_hd__o211a_1 _4010_ (.A1(net88),
    .A2(_2009_),
    .B1(_2011_),
    .C1(net347),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _4011_ (.A(\axi_controller.reg_input_data[26] ),
    .B(_2008_),
    .X(_2012_));
 sky130_fd_sc_hd__o211a_1 _4012_ (.A1(net89),
    .A2(_2009_),
    .B1(_2012_),
    .C1(net346),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _4013_ (.A(\axi_controller.reg_input_data[27] ),
    .B(_2008_),
    .X(_2013_));
 sky130_fd_sc_hd__o211a_1 _4014_ (.A1(net90),
    .A2(_2009_),
    .B1(_2013_),
    .C1(net348),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _4015_ (.A(\axi_controller.reg_input_data[28] ),
    .B(_2008_),
    .X(_2014_));
 sky130_fd_sc_hd__o211a_1 _4016_ (.A1(net91),
    .A2(_2009_),
    .B1(_2014_),
    .C1(net348),
    .X(_0342_));
 sky130_fd_sc_hd__or2_1 _4017_ (.A(\axi_controller.reg_input_data[29] ),
    .B(_2008_),
    .X(_2015_));
 sky130_fd_sc_hd__o211a_1 _4018_ (.A1(net92),
    .A2(_2009_),
    .B1(_2015_),
    .C1(net346),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _4019_ (.A(\axi_controller.reg_input_data[30] ),
    .B(_2008_),
    .X(_2016_));
 sky130_fd_sc_hd__o211a_1 _4020_ (.A1(net94),
    .A2(_2009_),
    .B1(_2016_),
    .C1(net347),
    .X(_0344_));
 sky130_fd_sc_hd__or2_1 _4021_ (.A(\axi_controller.reg_input_data[31] ),
    .B(_2008_),
    .X(_2017_));
 sky130_fd_sc_hd__o211a_1 _4022_ (.A1(net95),
    .A2(_2009_),
    .B1(_2017_),
    .C1(net346),
    .X(_0345_));
 sky130_fd_sc_hd__and2_1 _4023_ (.A(net103),
    .B(_1963_),
    .X(_2018_));
 sky130_fd_sc_hd__nand2_2 _4024_ (.A(net103),
    .B(_1963_),
    .Y(_2019_));
 sky130_fd_sc_hd__or2_1 _4025_ (.A(\axi_controller.reg_input_data[0] ),
    .B(_2018_),
    .X(_2020_));
 sky130_fd_sc_hd__o211a_1 _4026_ (.A1(net71),
    .A2(_2019_),
    .B1(_2020_),
    .C1(net349),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _4027_ (.A(\axi_controller.reg_input_data[1] ),
    .B(_2018_),
    .X(_2021_));
 sky130_fd_sc_hd__o211a_1 _4028_ (.A1(net82),
    .A2(_2019_),
    .B1(_2021_),
    .C1(net349),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _4029_ (.A(\axi_controller.reg_input_data[2] ),
    .B(_2018_),
    .X(_2022_));
 sky130_fd_sc_hd__o211a_1 _4030_ (.A1(net93),
    .A2(_2019_),
    .B1(_2022_),
    .C1(net350),
    .X(_0348_));
 sky130_fd_sc_hd__or2_1 _4031_ (.A(\axi_controller.reg_input_data[3] ),
    .B(_2018_),
    .X(_2023_));
 sky130_fd_sc_hd__o211a_1 _4032_ (.A1(net96),
    .A2(_2019_),
    .B1(_2023_),
    .C1(net350),
    .X(_0349_));
 sky130_fd_sc_hd__or2_1 _4033_ (.A(\axi_controller.reg_input_data[4] ),
    .B(_2018_),
    .X(_2024_));
 sky130_fd_sc_hd__o211a_1 _4034_ (.A1(net97),
    .A2(_2019_),
    .B1(_2024_),
    .C1(net350),
    .X(_0350_));
 sky130_fd_sc_hd__or2_1 _4035_ (.A(\axi_controller.reg_input_data[5] ),
    .B(_2018_),
    .X(_2025_));
 sky130_fd_sc_hd__o211a_1 _4036_ (.A1(net98),
    .A2(_2019_),
    .B1(_2025_),
    .C1(net350),
    .X(_0351_));
 sky130_fd_sc_hd__or2_1 _4037_ (.A(\axi_controller.reg_input_data[6] ),
    .B(_2018_),
    .X(_2026_));
 sky130_fd_sc_hd__o211a_1 _4038_ (.A1(net99),
    .A2(_2019_),
    .B1(_2026_),
    .C1(net350),
    .X(_0352_));
 sky130_fd_sc_hd__or2_1 _4039_ (.A(\axi_controller.reg_input_data[7] ),
    .B(_2018_),
    .X(_2027_));
 sky130_fd_sc_hd__o211a_1 _4040_ (.A1(net100),
    .A2(_2019_),
    .B1(_2027_),
    .C1(net350),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_2 _4041_ (.A0(\cordic_inst.cordic_inst.cos_out[0] ),
    .A1(\cordic_inst.cordic_inst.sin_out[0] ),
    .S(net316),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(\axi_controller.result_out[0] ),
    .A1(_2028_),
    .S(net200),
    .X(_0354_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(\cordic_inst.cordic_inst.sin_out[0] ),
    .B(net261),
    .Y(_2029_));
 sky130_fd_sc_hd__xnor2_1 _4044_ (.A(\cordic_inst.cordic_inst.sin_out[1] ),
    .B(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__nand2_1 _4045_ (.A(\cordic_inst.cordic_inst.cos_out[0] ),
    .B(net223),
    .Y(_2031_));
 sky130_fd_sc_hd__xnor2_1 _4046_ (.A(\cordic_inst.cordic_inst.cos_out[1] ),
    .B(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__mux2_1 _4047_ (.A0(_2030_),
    .A1(_2032_),
    .S(net230),
    .X(_2033_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(\axi_controller.result_out[1] ),
    .A1(_2033_),
    .S(net202),
    .X(_0355_));
 sky130_fd_sc_hd__o21ai_1 _4049_ (.A1(\cordic_inst.cordic_inst.sin_out[1] ),
    .A2(\cordic_inst.cordic_inst.sin_out[0] ),
    .B1(net261),
    .Y(_2034_));
 sky130_fd_sc_hd__xnor2_1 _4050_ (.A(\cordic_inst.cordic_inst.sin_out[2] ),
    .B(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__o21a_1 _4051_ (.A1(\cordic_inst.cordic_inst.cos_out[1] ),
    .A2(\cordic_inst.cordic_inst.cos_out[0] ),
    .B1(net224),
    .X(_2036_));
 sky130_fd_sc_hd__xor2_1 _4052_ (.A(\cordic_inst.cordic_inst.cos_out[2] ),
    .B(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__mux2_1 _4053_ (.A0(_2035_),
    .A1(_2037_),
    .S(net230),
    .X(_2038_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(\axi_controller.result_out[2] ),
    .A1(_2038_),
    .S(net203),
    .X(_0356_));
 sky130_fd_sc_hd__o31a_1 _4055_ (.A1(\cordic_inst.cordic_inst.sin_out[2] ),
    .A2(\cordic_inst.cordic_inst.sin_out[1] ),
    .A3(\cordic_inst.cordic_inst.sin_out[0] ),
    .B1(net261),
    .X(_2039_));
 sky130_fd_sc_hd__xor2_1 _4056_ (.A(\cordic_inst.cordic_inst.sin_out[3] ),
    .B(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__o31a_1 _4057_ (.A1(\cordic_inst.cordic_inst.cos_out[2] ),
    .A2(\cordic_inst.cordic_inst.cos_out[1] ),
    .A3(\cordic_inst.cordic_inst.cos_out[0] ),
    .B1(net223),
    .X(_2041_));
 sky130_fd_sc_hd__xor2_1 _4058_ (.A(\cordic_inst.cordic_inst.cos_out[3] ),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__mux2_1 _4059_ (.A0(_2040_),
    .A1(_2042_),
    .S(net230),
    .X(_2043_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(\axi_controller.result_out[3] ),
    .A1(_2043_),
    .S(net202),
    .X(_0357_));
 sky130_fd_sc_hd__nor2_1 _4061_ (.A(\axi_controller.result_out[4] ),
    .B(net202),
    .Y(_2044_));
 sky130_fd_sc_hd__or4_2 _4062_ (.A(\cordic_inst.cordic_inst.sin_out[3] ),
    .B(\cordic_inst.cordic_inst.sin_out[2] ),
    .C(\cordic_inst.cordic_inst.sin_out[1] ),
    .D(\cordic_inst.cordic_inst.sin_out[0] ),
    .X(_2045_));
 sky130_fd_sc_hd__and3_1 _4063_ (.A(\cordic_inst.cordic_inst.sin_out[4] ),
    .B(net259),
    .C(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__a21oi_1 _4064_ (.A1(net259),
    .A2(_2045_),
    .B1(\cordic_inst.cordic_inst.sin_out[4] ),
    .Y(_2047_));
 sky130_fd_sc_hd__or4_4 _4065_ (.A(\cordic_inst.cordic_inst.cos_out[3] ),
    .B(\cordic_inst.cordic_inst.cos_out[2] ),
    .C(\cordic_inst.cordic_inst.cos_out[1] ),
    .D(\cordic_inst.cordic_inst.cos_out[0] ),
    .X(_2048_));
 sky130_fd_sc_hd__a21oi_1 _4066_ (.A1(net226),
    .A2(_2048_),
    .B1(\cordic_inst.cordic_inst.cos_out[4] ),
    .Y(_2049_));
 sky130_fd_sc_hd__a31o_1 _4067_ (.A1(\cordic_inst.cordic_inst.cos_out[4] ),
    .A2(net226),
    .A3(_2048_),
    .B1(net314),
    .X(_2050_));
 sky130_fd_sc_hd__o32a_1 _4068_ (.A1(net228),
    .A2(_2046_),
    .A3(_2047_),
    .B1(_2049_),
    .B2(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__a21oi_1 _4069_ (.A1(net202),
    .A2(_2051_),
    .B1(_2044_),
    .Y(_0358_));
 sky130_fd_sc_hd__o21ai_1 _4070_ (.A1(\cordic_inst.cordic_inst.sin_out[4] ),
    .A2(_2045_),
    .B1(net259),
    .Y(_2052_));
 sky130_fd_sc_hd__xnor2_1 _4071_ (.A(\cordic_inst.cordic_inst.sin_out[5] ),
    .B(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__o21a_1 _4072_ (.A1(\cordic_inst.cordic_inst.cos_out[4] ),
    .A2(_2048_),
    .B1(net225),
    .X(_2054_));
 sky130_fd_sc_hd__or2_1 _4073_ (.A(\cordic_inst.cordic_inst.cos_out[5] ),
    .B(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__a21oi_1 _4074_ (.A1(\cordic_inst.cordic_inst.cos_out[5] ),
    .A2(_2054_),
    .B1(net314),
    .Y(_2056_));
 sky130_fd_sc_hd__a22o_1 _4075_ (.A1(net314),
    .A2(_2053_),
    .B1(_2055_),
    .B2(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(\axi_controller.result_out[5] ),
    .A1(_2057_),
    .S(net202),
    .X(_0359_));
 sky130_fd_sc_hd__o31a_1 _4077_ (.A1(\cordic_inst.cordic_inst.cos_out[5] ),
    .A2(\cordic_inst.cordic_inst.cos_out[4] ),
    .A3(_2048_),
    .B1(net225),
    .X(_2058_));
 sky130_fd_sc_hd__xor2_1 _4078_ (.A(\cordic_inst.cordic_inst.cos_out[6] ),
    .B(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__o31a_1 _4079_ (.A1(\cordic_inst.cordic_inst.sin_out[5] ),
    .A2(\cordic_inst.cordic_inst.sin_out[4] ),
    .A3(_2045_),
    .B1(net259),
    .X(_2060_));
 sky130_fd_sc_hd__or2_1 _4080_ (.A(\cordic_inst.cordic_inst.sin_out[6] ),
    .B(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__a21oi_1 _4081_ (.A1(\cordic_inst.cordic_inst.sin_out[6] ),
    .A2(_2060_),
    .B1(net228),
    .Y(_2062_));
 sky130_fd_sc_hd__a22o_1 _4082_ (.A1(net228),
    .A2(_2059_),
    .B1(_2061_),
    .B2(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(\axi_controller.result_out[6] ),
    .A1(_2063_),
    .S(net202),
    .X(_0360_));
 sky130_fd_sc_hd__nor2_1 _4084_ (.A(\axi_controller.result_out[7] ),
    .B(net202),
    .Y(_2064_));
 sky130_fd_sc_hd__or4_1 _4085_ (.A(\cordic_inst.cordic_inst.sin_out[6] ),
    .B(\cordic_inst.cordic_inst.sin_out[5] ),
    .C(\cordic_inst.cordic_inst.sin_out[4] ),
    .D(_2045_),
    .X(_2065_));
 sky130_fd_sc_hd__and3_1 _4086_ (.A(\cordic_inst.cordic_inst.sin_out[7] ),
    .B(net258),
    .C(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__a21oi_1 _4087_ (.A1(net258),
    .A2(_2065_),
    .B1(\cordic_inst.cordic_inst.sin_out[7] ),
    .Y(_2067_));
 sky130_fd_sc_hd__or4_2 _4088_ (.A(\cordic_inst.cordic_inst.cos_out[6] ),
    .B(\cordic_inst.cordic_inst.cos_out[5] ),
    .C(\cordic_inst.cordic_inst.cos_out[4] ),
    .D(_2048_),
    .X(_2068_));
 sky130_fd_sc_hd__a21oi_1 _4089_ (.A1(net225),
    .A2(_2068_),
    .B1(\cordic_inst.cordic_inst.cos_out[7] ),
    .Y(_2069_));
 sky130_fd_sc_hd__a31o_1 _4090_ (.A1(\cordic_inst.cordic_inst.cos_out[7] ),
    .A2(net225),
    .A3(_2068_),
    .B1(net314),
    .X(_2070_));
 sky130_fd_sc_hd__o32a_1 _4091_ (.A1(net229),
    .A2(_2066_),
    .A3(_2067_),
    .B1(_2069_),
    .B2(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__a21oi_1 _4092_ (.A1(net202),
    .A2(_2071_),
    .B1(_2064_),
    .Y(_0361_));
 sky130_fd_sc_hd__o21a_1 _4093_ (.A1(\cordic_inst.cordic_inst.cos_out[7] ),
    .A2(_2068_),
    .B1(net225),
    .X(_2072_));
 sky130_fd_sc_hd__o21ai_1 _4094_ (.A1(\cordic_inst.cordic_inst.cos_out[8] ),
    .A2(_2072_),
    .B1(net228),
    .Y(_2073_));
 sky130_fd_sc_hd__a21o_1 _4095_ (.A1(\cordic_inst.cordic_inst.cos_out[8] ),
    .A2(_2072_),
    .B1(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__or2_1 _4096_ (.A(\cordic_inst.cordic_inst.sin_out[7] ),
    .B(_2065_),
    .X(_2075_));
 sky130_fd_sc_hd__a21oi_1 _4097_ (.A1(net258),
    .A2(_2075_),
    .B1(\cordic_inst.cordic_inst.sin_out[8] ),
    .Y(_2076_));
 sky130_fd_sc_hd__a31o_1 _4098_ (.A1(\cordic_inst.cordic_inst.sin_out[8] ),
    .A2(net258),
    .A3(_2075_),
    .B1(net228),
    .X(_2077_));
 sky130_fd_sc_hd__o211a_1 _4099_ (.A1(_2076_),
    .A2(_2077_),
    .B1(net203),
    .C1(_2074_),
    .X(_2078_));
 sky130_fd_sc_hd__o21ba_1 _4100_ (.A1(\axi_controller.result_out[8] ),
    .A2(net202),
    .B1_N(_2078_),
    .X(_0362_));
 sky130_fd_sc_hd__o31a_1 _4101_ (.A1(\cordic_inst.cordic_inst.cos_out[8] ),
    .A2(\cordic_inst.cordic_inst.cos_out[7] ),
    .A3(_2068_),
    .B1(net225),
    .X(_2079_));
 sky130_fd_sc_hd__xor2_1 _4102_ (.A(\cordic_inst.cordic_inst.cos_out[9] ),
    .B(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__or2_1 _4103_ (.A(\cordic_inst.cordic_inst.sin_out[8] ),
    .B(_2075_),
    .X(_2081_));
 sky130_fd_sc_hd__a21oi_1 _4104_ (.A1(net258),
    .A2(_2081_),
    .B1(\cordic_inst.cordic_inst.sin_out[9] ),
    .Y(_2082_));
 sky130_fd_sc_hd__a31o_1 _4105_ (.A1(\cordic_inst.cordic_inst.sin_out[9] ),
    .A2(net258),
    .A3(_2081_),
    .B1(net228),
    .X(_2083_));
 sky130_fd_sc_hd__a2bb2o_1 _4106_ (.A1_N(_2083_),
    .A2_N(_2082_),
    .B1(_2080_),
    .B2(net228),
    .X(_2084_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(\axi_controller.result_out[9] ),
    .A1(_2084_),
    .S(net202),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_1 _4108_ (.A(\axi_controller.result_out[10] ),
    .B(net203),
    .Y(_2085_));
 sky130_fd_sc_hd__or4_1 _4109_ (.A(\cordic_inst.cordic_inst.sin_out[9] ),
    .B(\cordic_inst.cordic_inst.sin_out[8] ),
    .C(\cordic_inst.cordic_inst.sin_out[7] ),
    .D(_2065_),
    .X(_2086_));
 sky130_fd_sc_hd__and3_1 _4110_ (.A(\cordic_inst.cordic_inst.sin_out[10] ),
    .B(net258),
    .C(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__a21oi_1 _4111_ (.A1(net259),
    .A2(_2086_),
    .B1(\cordic_inst.cordic_inst.sin_out[10] ),
    .Y(_2088_));
 sky130_fd_sc_hd__or4_2 _4112_ (.A(\cordic_inst.cordic_inst.cos_out[9] ),
    .B(\cordic_inst.cordic_inst.cos_out[8] ),
    .C(\cordic_inst.cordic_inst.cos_out[7] ),
    .D(_2068_),
    .X(_2089_));
 sky130_fd_sc_hd__a21oi_1 _4113_ (.A1(net226),
    .A2(_2089_),
    .B1(\cordic_inst.cordic_inst.cos_out[10] ),
    .Y(_2090_));
 sky130_fd_sc_hd__a31o_1 _4114_ (.A1(\cordic_inst.cordic_inst.cos_out[10] ),
    .A2(net225),
    .A3(_2089_),
    .B1(net314),
    .X(_2091_));
 sky130_fd_sc_hd__o32a_1 _4115_ (.A1(net228),
    .A2(_2087_),
    .A3(_2088_),
    .B1(_2090_),
    .B2(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__a21oi_1 _4116_ (.A1(net203),
    .A2(_2092_),
    .B1(_2085_),
    .Y(_0364_));
 sky130_fd_sc_hd__or2_1 _4117_ (.A(\cordic_inst.cordic_inst.sin_out[10] ),
    .B(_2086_),
    .X(_2093_));
 sky130_fd_sc_hd__a21oi_1 _4118_ (.A1(net258),
    .A2(_2093_),
    .B1(\cordic_inst.cordic_inst.sin_out[11] ),
    .Y(_2094_));
 sky130_fd_sc_hd__a31o_1 _4119_ (.A1(\cordic_inst.cordic_inst.sin_out[11] ),
    .A2(net258),
    .A3(_2093_),
    .B1(net228),
    .X(_2095_));
 sky130_fd_sc_hd__o21a_1 _4120_ (.A1(\cordic_inst.cordic_inst.cos_out[10] ),
    .A2(_2089_),
    .B1(net225),
    .X(_2096_));
 sky130_fd_sc_hd__xnor2_1 _4121_ (.A(\cordic_inst.cordic_inst.cos_out[11] ),
    .B(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__o22ai_1 _4122_ (.A1(_2094_),
    .A2(_2095_),
    .B1(_2097_),
    .B2(net314),
    .Y(_2098_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(\axi_controller.result_out[11] ),
    .A1(_2098_),
    .S(net203),
    .X(_0365_));
 sky130_fd_sc_hd__or3_1 _4124_ (.A(\cordic_inst.cordic_inst.sin_out[11] ),
    .B(\cordic_inst.cordic_inst.sin_out[10] ),
    .C(_2086_),
    .X(_2099_));
 sky130_fd_sc_hd__and3_1 _4125_ (.A(\cordic_inst.cordic_inst.sin_out[12] ),
    .B(net258),
    .C(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__a21oi_1 _4126_ (.A1(net259),
    .A2(_2099_),
    .B1(\cordic_inst.cordic_inst.sin_out[12] ),
    .Y(_2101_));
 sky130_fd_sc_hd__or3_1 _4127_ (.A(net228),
    .B(_2100_),
    .C(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__or3_1 _4128_ (.A(\cordic_inst.cordic_inst.cos_out[11] ),
    .B(\cordic_inst.cordic_inst.cos_out[10] ),
    .C(_2089_),
    .X(_2103_));
 sky130_fd_sc_hd__a21oi_1 _4129_ (.A1(net225),
    .A2(_2103_),
    .B1(\cordic_inst.cordic_inst.cos_out[12] ),
    .Y(_2104_));
 sky130_fd_sc_hd__a31o_1 _4130_ (.A1(\cordic_inst.cordic_inst.cos_out[12] ),
    .A2(net225),
    .A3(_2103_),
    .B1(net314),
    .X(_2105_));
 sky130_fd_sc_hd__o21a_1 _4131_ (.A1(_2104_),
    .A2(_2105_),
    .B1(net203),
    .X(_2106_));
 sky130_fd_sc_hd__o2bb2a_1 _4132_ (.A1_N(_2102_),
    .A2_N(_2106_),
    .B1(\axi_controller.result_out[12] ),
    .B2(net203),
    .X(_0366_));
 sky130_fd_sc_hd__or2_1 _4133_ (.A(\cordic_inst.cordic_inst.sin_out[12] ),
    .B(_2099_),
    .X(_2107_));
 sky130_fd_sc_hd__a21oi_1 _4134_ (.A1(net260),
    .A2(_2107_),
    .B1(\cordic_inst.cordic_inst.sin_out[13] ),
    .Y(_2108_));
 sky130_fd_sc_hd__a31o_1 _4135_ (.A1(\cordic_inst.cordic_inst.sin_out[13] ),
    .A2(net260),
    .A3(_2107_),
    .B1(net229),
    .X(_2109_));
 sky130_fd_sc_hd__or2_1 _4136_ (.A(_2108_),
    .B(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__or4_2 _4137_ (.A(\cordic_inst.cordic_inst.cos_out[12] ),
    .B(\cordic_inst.cordic_inst.cos_out[11] ),
    .C(\cordic_inst.cordic_inst.cos_out[10] ),
    .D(_2089_),
    .X(_2111_));
 sky130_fd_sc_hd__a21oi_1 _4138_ (.A1(net227),
    .A2(_2111_),
    .B1(\cordic_inst.cordic_inst.cos_out[13] ),
    .Y(_2112_));
 sky130_fd_sc_hd__a31o_1 _4139_ (.A1(\cordic_inst.cordic_inst.cos_out[13] ),
    .A2(net227),
    .A3(_2111_),
    .B1(net315),
    .X(_2113_));
 sky130_fd_sc_hd__o21ai_1 _4140_ (.A1(_2112_),
    .A2(_2113_),
    .B1(_2110_),
    .Y(_2114_));
 sky130_fd_sc_hd__mux2_1 _4141_ (.A0(\axi_controller.result_out[13] ),
    .A1(_2114_),
    .S(net204),
    .X(_0367_));
 sky130_fd_sc_hd__o21a_1 _4142_ (.A1(\cordic_inst.cordic_inst.sin_out[13] ),
    .A2(_2107_),
    .B1(net261),
    .X(_2115_));
 sky130_fd_sc_hd__xor2_1 _4143_ (.A(\cordic_inst.cordic_inst.sin_out[14] ),
    .B(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__o21a_1 _4144_ (.A1(\cordic_inst.cordic_inst.cos_out[13] ),
    .A2(_2111_),
    .B1(net227),
    .X(_2117_));
 sky130_fd_sc_hd__xor2_1 _4145_ (.A(\cordic_inst.cordic_inst.cos_out[14] ),
    .B(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(_2116_),
    .A1(_2118_),
    .S(net229),
    .X(_2119_));
 sky130_fd_sc_hd__mux2_1 _4147_ (.A0(\axi_controller.result_out[14] ),
    .A1(_2119_),
    .S(net204),
    .X(_0368_));
 sky130_fd_sc_hd__or3_1 _4148_ (.A(\cordic_inst.cordic_inst.cos_out[14] ),
    .B(\cordic_inst.cordic_inst.cos_out[13] ),
    .C(_2111_),
    .X(_2120_));
 sky130_fd_sc_hd__a21oi_1 _4149_ (.A1(net227),
    .A2(_2120_),
    .B1(\cordic_inst.cordic_inst.cos_out[15] ),
    .Y(_2121_));
 sky130_fd_sc_hd__a31o_1 _4150_ (.A1(\cordic_inst.cordic_inst.cos_out[15] ),
    .A2(net226),
    .A3(_2120_),
    .B1(net315),
    .X(_2122_));
 sky130_fd_sc_hd__or3_1 _4151_ (.A(\cordic_inst.cordic_inst.sin_out[14] ),
    .B(\cordic_inst.cordic_inst.sin_out[13] ),
    .C(_2107_),
    .X(_2123_));
 sky130_fd_sc_hd__a21oi_1 _4152_ (.A1(net260),
    .A2(_2123_),
    .B1(\cordic_inst.cordic_inst.sin_out[15] ),
    .Y(_2124_));
 sky130_fd_sc_hd__a31o_1 _4153_ (.A1(\cordic_inst.cordic_inst.sin_out[15] ),
    .A2(net260),
    .A3(_2123_),
    .B1(net229),
    .X(_2125_));
 sky130_fd_sc_hd__or2_1 _4154_ (.A(_2124_),
    .B(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__o211a_1 _4155_ (.A1(_2121_),
    .A2(_2122_),
    .B1(_2126_),
    .C1(net204),
    .X(_2127_));
 sky130_fd_sc_hd__o21ba_1 _4156_ (.A1(\axi_controller.result_out[15] ),
    .A2(net204),
    .B1_N(_2127_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _4157_ (.A(\cordic_inst.cordic_inst.sin_out[15] ),
    .B(_2123_),
    .X(_2128_));
 sky130_fd_sc_hd__a21o_1 _4158_ (.A1(net260),
    .A2(_2128_),
    .B1(\cordic_inst.cordic_inst.sin_out[16] ),
    .X(_2129_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(net315),
    .B(_2129_),
    .Y(_2130_));
 sky130_fd_sc_hd__a31o_1 _4160_ (.A1(\cordic_inst.cordic_inst.sin_out[16] ),
    .A2(net260),
    .A3(_2128_),
    .B1(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__or4_2 _4161_ (.A(\cordic_inst.cordic_inst.cos_out[15] ),
    .B(\cordic_inst.cordic_inst.cos_out[14] ),
    .C(\cordic_inst.cordic_inst.cos_out[13] ),
    .D(_2111_),
    .X(_2132_));
 sky130_fd_sc_hd__a21oi_1 _4162_ (.A1(net226),
    .A2(_2132_),
    .B1(\cordic_inst.cordic_inst.cos_out[16] ),
    .Y(_2133_));
 sky130_fd_sc_hd__a31o_1 _4163_ (.A1(\cordic_inst.cordic_inst.cos_out[16] ),
    .A2(net226),
    .A3(_2132_),
    .B1(net315),
    .X(_2134_));
 sky130_fd_sc_hd__o21ai_1 _4164_ (.A1(_2133_),
    .A2(_2134_),
    .B1(_2131_),
    .Y(_2135_));
 sky130_fd_sc_hd__mux2_1 _4165_ (.A0(\axi_controller.result_out[16] ),
    .A1(_2135_),
    .S(net204),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _4166_ (.A(\cordic_inst.cordic_inst.sin_out[16] ),
    .B(_2128_),
    .X(_2136_));
 sky130_fd_sc_hd__a21oi_1 _4167_ (.A1(net260),
    .A2(_2136_),
    .B1(\cordic_inst.cordic_inst.sin_out[17] ),
    .Y(_2137_));
 sky130_fd_sc_hd__a31o_1 _4168_ (.A1(\cordic_inst.cordic_inst.sin_out[17] ),
    .A2(net260),
    .A3(_2136_),
    .B1(net229),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _4169_ (.A(_2137_),
    .B(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__o21a_1 _4170_ (.A1(\cordic_inst.cordic_inst.cos_out[16] ),
    .A2(_2132_),
    .B1(net226),
    .X(_2140_));
 sky130_fd_sc_hd__xnor2_1 _4171_ (.A(\cordic_inst.cordic_inst.cos_out[17] ),
    .B(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__o21a_1 _4172_ (.A1(net314),
    .A2(_2141_),
    .B1(net204),
    .X(_2142_));
 sky130_fd_sc_hd__o2bb2a_1 _4173_ (.A1_N(_2139_),
    .A2_N(_2142_),
    .B1(\axi_controller.result_out[17] ),
    .B2(net204),
    .X(_0371_));
 sky130_fd_sc_hd__or3_1 _4174_ (.A(\cordic_inst.cordic_inst.sin_out[17] ),
    .B(\cordic_inst.cordic_inst.sin_out[16] ),
    .C(_2128_),
    .X(_2143_));
 sky130_fd_sc_hd__a21o_1 _4175_ (.A1(net260),
    .A2(_2143_),
    .B1(\cordic_inst.cordic_inst.sin_out[18] ),
    .X(_2144_));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(net315),
    .B(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__a31o_1 _4177_ (.A1(\cordic_inst.cordic_inst.sin_out[18] ),
    .A2(net260),
    .A3(_2143_),
    .B1(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__or3_1 _4178_ (.A(\cordic_inst.cordic_inst.cos_out[17] ),
    .B(\cordic_inst.cordic_inst.cos_out[16] ),
    .C(_2132_),
    .X(_2147_));
 sky130_fd_sc_hd__a21oi_1 _4179_ (.A1(net226),
    .A2(_2147_),
    .B1(\cordic_inst.cordic_inst.cos_out[18] ),
    .Y(_2148_));
 sky130_fd_sc_hd__a31o_1 _4180_ (.A1(\cordic_inst.cordic_inst.cos_out[18] ),
    .A2(net226),
    .A3(_2147_),
    .B1(net315),
    .X(_2149_));
 sky130_fd_sc_hd__o21a_1 _4181_ (.A1(_2148_),
    .A2(_2149_),
    .B1(net204),
    .X(_2150_));
 sky130_fd_sc_hd__o2bb2a_1 _4182_ (.A1_N(_2146_),
    .A2_N(_2150_),
    .B1(\axi_controller.result_out[18] ),
    .B2(net204),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _4183_ (.A(\cordic_inst.cordic_inst.sin_out[18] ),
    .B(_2143_),
    .X(_2151_));
 sky130_fd_sc_hd__and3_1 _4184_ (.A(\cordic_inst.cordic_inst.sin_out[19] ),
    .B(net261),
    .C(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__a21oi_1 _4185_ (.A1(net261),
    .A2(_2151_),
    .B1(\cordic_inst.cordic_inst.sin_out[19] ),
    .Y(_2153_));
 sky130_fd_sc_hd__or3_1 _4186_ (.A(net230),
    .B(_2152_),
    .C(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__or2_1 _4187_ (.A(\cordic_inst.cordic_inst.cos_out[18] ),
    .B(_2147_),
    .X(_2155_));
 sky130_fd_sc_hd__a21oi_1 _4188_ (.A1(net227),
    .A2(_2155_),
    .B1(\cordic_inst.cordic_inst.cos_out[19] ),
    .Y(_2156_));
 sky130_fd_sc_hd__a31o_1 _4189_ (.A1(\cordic_inst.cordic_inst.cos_out[19] ),
    .A2(net227),
    .A3(_2155_),
    .B1(net314),
    .X(_2157_));
 sky130_fd_sc_hd__o21a_1 _4190_ (.A1(_2156_),
    .A2(_2157_),
    .B1(net205),
    .X(_2158_));
 sky130_fd_sc_hd__o2bb2a_1 _4191_ (.A1_N(_2154_),
    .A2_N(_2158_),
    .B1(\axi_controller.result_out[19] ),
    .B2(net205),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _4192_ (.A(\cordic_inst.cordic_inst.sin_out[19] ),
    .B(_2151_),
    .X(_2159_));
 sky130_fd_sc_hd__a21o_1 _4193_ (.A1(net261),
    .A2(_2159_),
    .B1(\cordic_inst.cordic_inst.sin_out[20] ),
    .X(_2160_));
 sky130_fd_sc_hd__nand2_1 _4194_ (.A(net316),
    .B(_2160_),
    .Y(_2161_));
 sky130_fd_sc_hd__a31o_1 _4195_ (.A1(\cordic_inst.cordic_inst.sin_out[20] ),
    .A2(net261),
    .A3(_2159_),
    .B1(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__o21a_1 _4196_ (.A1(\cordic_inst.cordic_inst.cos_out[19] ),
    .A2(_2155_),
    .B1(net227),
    .X(_2163_));
 sky130_fd_sc_hd__xnor2_1 _4197_ (.A(\cordic_inst.cordic_inst.cos_out[20] ),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__o21a_1 _4198_ (.A1(net314),
    .A2(_2164_),
    .B1(net205),
    .X(_2165_));
 sky130_fd_sc_hd__o2bb2a_1 _4199_ (.A1_N(_2162_),
    .A2_N(_2165_),
    .B1(\axi_controller.result_out[20] ),
    .B2(net205),
    .X(_0374_));
 sky130_fd_sc_hd__or3_1 _4200_ (.A(\cordic_inst.cordic_inst.cos_out[20] ),
    .B(\cordic_inst.cordic_inst.cos_out[19] ),
    .C(_2155_),
    .X(_2166_));
 sky130_fd_sc_hd__a21o_1 _4201_ (.A1(net227),
    .A2(_2166_),
    .B1(\cordic_inst.cordic_inst.cos_out[21] ),
    .X(_2167_));
 sky130_fd_sc_hd__a31oi_1 _4202_ (.A1(\cordic_inst.cordic_inst.cos_out[21] ),
    .A2(net227),
    .A3(_2166_),
    .B1(net316),
    .Y(_2168_));
 sky130_fd_sc_hd__or3_1 _4203_ (.A(\cordic_inst.cordic_inst.sin_out[20] ),
    .B(\cordic_inst.cordic_inst.sin_out[19] ),
    .C(_2151_),
    .X(_2169_));
 sky130_fd_sc_hd__a21o_1 _4204_ (.A1(net261),
    .A2(_2169_),
    .B1(\cordic_inst.cordic_inst.sin_out[21] ),
    .X(_2170_));
 sky130_fd_sc_hd__nand3_1 _4205_ (.A(\cordic_inst.cordic_inst.sin_out[21] ),
    .B(net261),
    .C(_2169_),
    .Y(_2171_));
 sky130_fd_sc_hd__a32o_1 _4206_ (.A1(net316),
    .A2(_2170_),
    .A3(_2171_),
    .B1(_2167_),
    .B2(_2168_),
    .X(_2172_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(\axi_controller.result_out[21] ),
    .A1(_2172_),
    .S(net205),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _4208_ (.A(\cordic_inst.cordic_inst.cos_out[21] ),
    .B(_2166_),
    .X(_2173_));
 sky130_fd_sc_hd__a21o_1 _4209_ (.A1(net224),
    .A2(_2173_),
    .B1(\cordic_inst.cordic_inst.cos_out[22] ),
    .X(_2174_));
 sky130_fd_sc_hd__a31oi_1 _4210_ (.A1(\cordic_inst.cordic_inst.cos_out[22] ),
    .A2(net224),
    .A3(_2173_),
    .B1(net316),
    .Y(_2175_));
 sky130_fd_sc_hd__or2_1 _4211_ (.A(\cordic_inst.cordic_inst.sin_out[21] ),
    .B(_2169_),
    .X(_2176_));
 sky130_fd_sc_hd__a21o_1 _4212_ (.A1(net257),
    .A2(_2176_),
    .B1(\cordic_inst.cordic_inst.sin_out[22] ),
    .X(_2177_));
 sky130_fd_sc_hd__nand3_1 _4213_ (.A(\cordic_inst.cordic_inst.sin_out[22] ),
    .B(net257),
    .C(_2176_),
    .Y(_2178_));
 sky130_fd_sc_hd__a32o_1 _4214_ (.A1(net316),
    .A2(_2177_),
    .A3(_2178_),
    .B1(_2174_),
    .B2(_2175_),
    .X(_2179_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(\axi_controller.result_out[22] ),
    .A1(_2179_),
    .S(net201),
    .X(_0376_));
 sky130_fd_sc_hd__or2_1 _4216_ (.A(\cordic_inst.cordic_inst.sin_out[22] ),
    .B(_2176_),
    .X(_2180_));
 sky130_fd_sc_hd__a21o_1 _4217_ (.A1(net257),
    .A2(_2180_),
    .B1(\cordic_inst.cordic_inst.sin_out[23] ),
    .X(_2181_));
 sky130_fd_sc_hd__nand2_1 _4218_ (.A(net316),
    .B(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__a31o_1 _4219_ (.A1(\cordic_inst.cordic_inst.sin_out[23] ),
    .A2(net257),
    .A3(_2180_),
    .B1(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__o21a_1 _4220_ (.A1(\cordic_inst.cordic_inst.cos_out[22] ),
    .A2(_2173_),
    .B1(net224),
    .X(_2184_));
 sky130_fd_sc_hd__xnor2_1 _4221_ (.A(\cordic_inst.cordic_inst.cos_out[23] ),
    .B(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__o21a_1 _4222_ (.A1(net316),
    .A2(_2185_),
    .B1(net201),
    .X(_2186_));
 sky130_fd_sc_hd__o2bb2a_1 _4223_ (.A1_N(_2183_),
    .A2_N(_2186_),
    .B1(\axi_controller.result_out[23] ),
    .B2(net201),
    .X(_0377_));
 sky130_fd_sc_hd__nor2_1 _4224_ (.A(\axi_controller.result_out[24] ),
    .B(net201),
    .Y(_2187_));
 sky130_fd_sc_hd__or3_1 _4225_ (.A(\cordic_inst.cordic_inst.cos_out[23] ),
    .B(\cordic_inst.cordic_inst.cos_out[22] ),
    .C(_2173_),
    .X(_2188_));
 sky130_fd_sc_hd__a21oi_1 _4226_ (.A1(net224),
    .A2(_2188_),
    .B1(\cordic_inst.cordic_inst.cos_out[24] ),
    .Y(_2189_));
 sky130_fd_sc_hd__a31o_1 _4227_ (.A1(\cordic_inst.cordic_inst.cos_out[24] ),
    .A2(net223),
    .A3(_2188_),
    .B1(net316),
    .X(_2190_));
 sky130_fd_sc_hd__or3_1 _4228_ (.A(\cordic_inst.cordic_inst.sin_out[23] ),
    .B(\cordic_inst.cordic_inst.sin_out[22] ),
    .C(_2176_),
    .X(_2191_));
 sky130_fd_sc_hd__a21oi_1 _4229_ (.A1(net257),
    .A2(_2191_),
    .B1(\cordic_inst.cordic_inst.sin_out[24] ),
    .Y(_2192_));
 sky130_fd_sc_hd__and3_1 _4230_ (.A(\cordic_inst.cordic_inst.sin_out[24] ),
    .B(net257),
    .C(_2191_),
    .X(_2193_));
 sky130_fd_sc_hd__or2_1 _4231_ (.A(_2192_),
    .B(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__o22a_1 _4232_ (.A1(_2189_),
    .A2(_2190_),
    .B1(_2194_),
    .B2(net231),
    .X(_2195_));
 sky130_fd_sc_hd__a21oi_1 _4233_ (.A1(net201),
    .A2(_2195_),
    .B1(_2187_),
    .Y(_0378_));
 sky130_fd_sc_hd__or2_1 _4234_ (.A(\cordic_inst.cordic_inst.cos_out[24] ),
    .B(_2188_),
    .X(_2196_));
 sky130_fd_sc_hd__and3_1 _4235_ (.A(\cordic_inst.cordic_inst.cos_out[25] ),
    .B(net223),
    .C(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__a21oi_1 _4236_ (.A1(net223),
    .A2(_2196_),
    .B1(\cordic_inst.cordic_inst.cos_out[25] ),
    .Y(_2198_));
 sky130_fd_sc_hd__or2_1 _4237_ (.A(\cordic_inst.cordic_inst.sin_out[24] ),
    .B(_2191_),
    .X(_2199_));
 sky130_fd_sc_hd__a21oi_1 _4238_ (.A1(net257),
    .A2(_2199_),
    .B1(\cordic_inst.cordic_inst.sin_out[25] ),
    .Y(_2200_));
 sky130_fd_sc_hd__a31o_1 _4239_ (.A1(\cordic_inst.cordic_inst.sin_out[25] ),
    .A2(net257),
    .A3(_2199_),
    .B1(net231),
    .X(_2201_));
 sky130_fd_sc_hd__o32ai_1 _4240_ (.A1(\axi_controller.mode ),
    .A2(_2197_),
    .A3(_2198_),
    .B1(_2200_),
    .B2(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__mux2_1 _4241_ (.A0(\axi_controller.result_out[25] ),
    .A1(_2202_),
    .S(net201),
    .X(_0379_));
 sky130_fd_sc_hd__nor2_1 _4242_ (.A(\cordic_inst.cordic_inst.cos_out[25] ),
    .B(_2196_),
    .Y(_2203_));
 sky130_fd_sc_hd__o21a_1 _4243_ (.A1(\cordic_inst.deg_handler_inst.kuadran[0] ),
    .A2(_2203_),
    .B1(_0605_),
    .X(_2204_));
 sky130_fd_sc_hd__nor2_1 _4244_ (.A(net313),
    .B(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__o31a_1 _4245_ (.A1(_0605_),
    .A2(\cordic_inst.deg_handler_inst.kuadran[0] ),
    .A3(_2203_),
    .B1(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__o21ai_1 _4246_ (.A1(\cordic_inst.cordic_inst.sin_out[25] ),
    .A2(_2199_),
    .B1(net256),
    .Y(_2207_));
 sky130_fd_sc_hd__xnor2_1 _4247_ (.A(\cordic_inst.cordic_inst.sin_out[26] ),
    .B(_2207_),
    .Y(_2208_));
 sky130_fd_sc_hd__a21o_1 _4248_ (.A1(net313),
    .A2(_2208_),
    .B1(_2206_),
    .X(_2209_));
 sky130_fd_sc_hd__mux2_1 _4249_ (.A0(\axi_controller.result_out[26] ),
    .A1(_2209_),
    .S(net201),
    .X(_0380_));
 sky130_fd_sc_hd__nor2_1 _4250_ (.A(\cordic_inst.deg_handler_inst.kuadran[0] ),
    .B(_2204_),
    .Y(_2210_));
 sky130_fd_sc_hd__nor2_1 _4251_ (.A(\cordic_inst.cordic_inst.cos_out[27] ),
    .B(_2210_),
    .Y(_2211_));
 sky130_fd_sc_hd__a21o_1 _4252_ (.A1(\cordic_inst.cordic_inst.cos_out[27] ),
    .A2(_2210_),
    .B1(net313),
    .X(_2212_));
 sky130_fd_sc_hd__or3_1 _4253_ (.A(\cordic_inst.cordic_inst.sin_out[26] ),
    .B(\cordic_inst.cordic_inst.sin_out[25] ),
    .C(_2199_),
    .X(_2213_));
 sky130_fd_sc_hd__a21o_1 _4254_ (.A1(net256),
    .A2(_2213_),
    .B1(\cordic_inst.cordic_inst.sin_out[27] ),
    .X(_2214_));
 sky130_fd_sc_hd__nand3_1 _4255_ (.A(\cordic_inst.cordic_inst.sin_out[27] ),
    .B(net256),
    .C(_2213_),
    .Y(_2215_));
 sky130_fd_sc_hd__and3_1 _4256_ (.A(net313),
    .B(_2214_),
    .C(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__o21ai_1 _4257_ (.A1(_2211_),
    .A2(_2212_),
    .B1(net200),
    .Y(_2217_));
 sky130_fd_sc_hd__o22a_1 _4258_ (.A1(\axi_controller.result_out[27] ),
    .A2(net200),
    .B1(_2216_),
    .B2(_2217_),
    .X(_0381_));
 sky130_fd_sc_hd__nor2_1 _4259_ (.A(\cordic_inst.deg_handler_inst.kuadran[0] ),
    .B(_2211_),
    .Y(_2218_));
 sky130_fd_sc_hd__xnor2_1 _4260_ (.A(\cordic_inst.cordic_inst.cos_out[28] ),
    .B(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__and3_1 _4261_ (.A(\cordic_inst.cordic_inst.sin_out[28] ),
    .B(net256),
    .C(_2214_),
    .X(_2220_));
 sky130_fd_sc_hd__a21o_1 _4262_ (.A1(net256),
    .A2(_2214_),
    .B1(\cordic_inst.cordic_inst.sin_out[28] ),
    .X(_2221_));
 sky130_fd_sc_hd__or3b_1 _4263_ (.A(net231),
    .B(_2220_),
    .C_N(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__o21ai_1 _4264_ (.A1(net313),
    .A2(_2219_),
    .B1(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(\axi_controller.result_out[28] ),
    .A1(_2223_),
    .S(net200),
    .X(_0382_));
 sky130_fd_sc_hd__a21o_1 _4266_ (.A1(net256),
    .A2(_2221_),
    .B1(\cordic_inst.cordic_inst.sin_out[29] ),
    .X(_2224_));
 sky130_fd_sc_hd__nand3_1 _4267_ (.A(\cordic_inst.cordic_inst.sin_out[29] ),
    .B(net256),
    .C(_2221_),
    .Y(_2225_));
 sky130_fd_sc_hd__o311a_1 _4268_ (.A1(\cordic_inst.cordic_inst.cos_out[28] ),
    .A2(\cordic_inst.cordic_inst.cos_out[27] ),
    .A3(_2210_),
    .B1(net223),
    .C1(\cordic_inst.cordic_inst.cos_out[29] ),
    .X(_2226_));
 sky130_fd_sc_hd__a211o_1 _4269_ (.A1(\cordic_inst.cordic_inst.cos_out[28] ),
    .A2(net223),
    .B1(_2218_),
    .C1(\cordic_inst.cordic_inst.cos_out[29] ),
    .X(_2227_));
 sky130_fd_sc_hd__nor3b_1 _4270_ (.A(net313),
    .B(_2226_),
    .C_N(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__a31o_1 _4271_ (.A1(net313),
    .A2(_2224_),
    .A3(_2225_),
    .B1(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(\axi_controller.result_out[29] ),
    .A1(_2229_),
    .S(net200),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_1 _4273_ (.A(\axi_controller.result_out[30] ),
    .B(net200),
    .Y(_2230_));
 sky130_fd_sc_hd__and3_1 _4274_ (.A(\cordic_inst.cordic_inst.cos_out[30] ),
    .B(net223),
    .C(_2227_),
    .X(_2231_));
 sky130_fd_sc_hd__a21oi_1 _4275_ (.A1(net223),
    .A2(_2227_),
    .B1(\cordic_inst.cordic_inst.cos_out[30] ),
    .Y(_2232_));
 sky130_fd_sc_hd__a21oi_1 _4276_ (.A1(net256),
    .A2(_2224_),
    .B1(\cordic_inst.cordic_inst.sin_out[30] ),
    .Y(_2233_));
 sky130_fd_sc_hd__a31o_1 _4277_ (.A1(\cordic_inst.cordic_inst.sin_out[30] ),
    .A2(net256),
    .A3(_2224_),
    .B1(net231),
    .X(_2234_));
 sky130_fd_sc_hd__o32a_1 _4278_ (.A1(net313),
    .A2(_2231_),
    .A3(_2232_),
    .B1(_2233_),
    .B2(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__a21oi_1 _4279_ (.A1(net200),
    .A2(_2235_),
    .B1(_2230_),
    .Y(_0384_));
 sky130_fd_sc_hd__o21ba_1 _4280_ (.A1(\cordic_inst.deg_handler_inst.kuadran[0] ),
    .A2(_2232_),
    .B1_N(\cordic_inst.cordic_inst.cos_out[31] ),
    .X(_2236_));
 sky130_fd_sc_hd__o211a_1 _4281_ (.A1(\cordic_inst.cordic_inst.cos_out[30] ),
    .A2(_2227_),
    .B1(net223),
    .C1(\cordic_inst.cordic_inst.cos_out[31] ),
    .X(_2237_));
 sky130_fd_sc_hd__o21a_1 _4282_ (.A1(\cordic_inst.cordic_inst.sin_out[30] ),
    .A2(_2224_),
    .B1(net256),
    .X(_2238_));
 sky130_fd_sc_hd__a21oi_1 _4283_ (.A1(\cordic_inst.cordic_inst.sin_out[31] ),
    .A2(_2238_),
    .B1(net231),
    .Y(_2239_));
 sky130_fd_sc_hd__o21ai_1 _4284_ (.A1(\cordic_inst.cordic_inst.sin_out[31] ),
    .A2(_2238_),
    .B1(_2239_),
    .Y(_2240_));
 sky130_fd_sc_hd__o31a_1 _4285_ (.A1(net313),
    .A2(_2236_),
    .A3(_2237_),
    .B1(net200),
    .X(_2241_));
 sky130_fd_sc_hd__o2bb2a_1 _4286_ (.A1_N(_2240_),
    .A2_N(_2241_),
    .B1(\axi_controller.result_out[31] ),
    .B2(net200),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _4287_ (.A(net105),
    .B(_1963_),
    .X(_2242_));
 sky130_fd_sc_hd__nand2_2 _4288_ (.A(net105),
    .B(_1963_),
    .Y(_2243_));
 sky130_fd_sc_hd__or2_1 _4289_ (.A(\axi_controller.reg_input_data[16] ),
    .B(_2242_),
    .X(_2244_));
 sky130_fd_sc_hd__o211a_1 _4290_ (.A1(net78),
    .A2(_2243_),
    .B1(_2244_),
    .C1(net347),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _4291_ (.A(\axi_controller.reg_input_data[17] ),
    .B(_2242_),
    .X(_2245_));
 sky130_fd_sc_hd__o211a_1 _4292_ (.A1(net79),
    .A2(_2243_),
    .B1(_2245_),
    .C1(net346),
    .X(_0392_));
 sky130_fd_sc_hd__or2_1 _4293_ (.A(\axi_controller.reg_input_data[18] ),
    .B(_2242_),
    .X(_2246_));
 sky130_fd_sc_hd__o211a_1 _4294_ (.A1(net80),
    .A2(_2243_),
    .B1(_2246_),
    .C1(net347),
    .X(_0393_));
 sky130_fd_sc_hd__or2_1 _4295_ (.A(\axi_controller.reg_input_data[19] ),
    .B(_2242_),
    .X(_2247_));
 sky130_fd_sc_hd__o211a_1 _4296_ (.A1(net81),
    .A2(_2243_),
    .B1(_2247_),
    .C1(net347),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _4297_ (.A(\axi_controller.reg_input_data[20] ),
    .B(_2242_),
    .X(_2248_));
 sky130_fd_sc_hd__o211a_1 _4298_ (.A1(net83),
    .A2(_2243_),
    .B1(_2248_),
    .C1(net346),
    .X(_0395_));
 sky130_fd_sc_hd__or2_1 _4299_ (.A(\axi_controller.reg_input_data[21] ),
    .B(_2242_),
    .X(_2249_));
 sky130_fd_sc_hd__o211a_1 _4300_ (.A1(net84),
    .A2(_2243_),
    .B1(_2249_),
    .C1(net348),
    .X(_0396_));
 sky130_fd_sc_hd__or2_1 _4301_ (.A(\axi_controller.reg_input_data[22] ),
    .B(_2242_),
    .X(_2250_));
 sky130_fd_sc_hd__o211a_1 _4302_ (.A1(net85),
    .A2(_2243_),
    .B1(_2250_),
    .C1(net348),
    .X(_0397_));
 sky130_fd_sc_hd__or2_1 _4303_ (.A(\axi_controller.reg_input_data[23] ),
    .B(_2242_),
    .X(_2251_));
 sky130_fd_sc_hd__o211a_1 _4304_ (.A1(net86),
    .A2(_2243_),
    .B1(_2251_),
    .C1(net346),
    .X(_0398_));
 sky130_fd_sc_hd__and4b_1 _4305_ (.A_N(\axi_controller.read_addr_reg[5] ),
    .B(_1977_),
    .C(\axi_controller.read_addr_reg[3] ),
    .D(\axi_controller.read_addr_reg[4] ),
    .X(_2252_));
 sky130_fd_sc_hd__nand2_1 _4306_ (.A(_1976_),
    .B(_2252_),
    .Y(_2253_));
 sky130_fd_sc_hd__nor2_1 _4307_ (.A(_1989_),
    .B(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__or4b_1 _4308_ (.A(\axi_controller.state[0] ),
    .B(\axi_controller.state[1] ),
    .C(_0621_),
    .D_N(net144),
    .X(_2255_));
 sky130_fd_sc_hd__o31ai_1 _4309_ (.A1(net194),
    .A2(_1990_),
    .A3(_2254_),
    .B1(_2255_),
    .Y(_0399_));
 sky130_fd_sc_hd__and4_1 _4310_ (.A(net82),
    .B(net103),
    .C(_1930_),
    .D(_1994_),
    .X(_0562_));
 sky130_fd_sc_hd__and4b_4 _4311_ (.A_N(net194),
    .B(_1976_),
    .C(_1987_),
    .D(_2252_),
    .X(_2256_));
 sky130_fd_sc_hd__a22o_1 _4312_ (.A1(net136),
    .A2(net194),
    .B1(net157),
    .B2(\axi_controller.result_out[31] ),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _4313_ (.A1(net135),
    .A2(net194),
    .B1(net157),
    .B2(\axi_controller.result_out[30] ),
    .X(_0564_));
 sky130_fd_sc_hd__a22o_1 _4314_ (.A1(net133),
    .A2(net194),
    .B1(net157),
    .B2(\axi_controller.result_out[29] ),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_1 _4315_ (.A1(net132),
    .A2(net194),
    .B1(net157),
    .B2(\axi_controller.result_out[28] ),
    .X(_0566_));
 sky130_fd_sc_hd__a22o_1 _4316_ (.A1(net131),
    .A2(net194),
    .B1(net157),
    .B2(\axi_controller.result_out[27] ),
    .X(_0567_));
 sky130_fd_sc_hd__a22o_1 _4317_ (.A1(net130),
    .A2(net194),
    .B1(net157),
    .B2(\axi_controller.result_out[26] ),
    .X(_0568_));
 sky130_fd_sc_hd__a22o_1 _4318_ (.A1(net129),
    .A2(net193),
    .B1(net157),
    .B2(\axi_controller.result_out[25] ),
    .X(_0569_));
 sky130_fd_sc_hd__a22o_1 _4319_ (.A1(net128),
    .A2(net193),
    .B1(net157),
    .B2(\axi_controller.result_out[24] ),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _4320_ (.A1(net127),
    .A2(net193),
    .B1(net157),
    .B2(\axi_controller.result_out[23] ),
    .X(_0571_));
 sky130_fd_sc_hd__a22o_1 _4321_ (.A1(net126),
    .A2(net193),
    .B1(net157),
    .B2(\axi_controller.result_out[22] ),
    .X(_0572_));
 sky130_fd_sc_hd__a22o_1 _4322_ (.A1(net125),
    .A2(net193),
    .B1(_2256_),
    .B2(\axi_controller.result_out[21] ),
    .X(_0573_));
 sky130_fd_sc_hd__a22o_1 _4323_ (.A1(net124),
    .A2(net193),
    .B1(_2256_),
    .B2(\axi_controller.result_out[20] ),
    .X(_0574_));
 sky130_fd_sc_hd__a22o_1 _4324_ (.A1(net122),
    .A2(net192),
    .B1(_2256_),
    .B2(\axi_controller.result_out[19] ),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _4325_ (.A1(net121),
    .A2(net192),
    .B1(net156),
    .B2(\axi_controller.result_out[18] ),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _4326_ (.A1(net120),
    .A2(net192),
    .B1(net156),
    .B2(\axi_controller.result_out[17] ),
    .X(_0577_));
 sky130_fd_sc_hd__a22o_1 _4327_ (.A1(net119),
    .A2(net192),
    .B1(net156),
    .B2(\axi_controller.result_out[16] ),
    .X(_0578_));
 sky130_fd_sc_hd__a22o_1 _4328_ (.A1(net118),
    .A2(net192),
    .B1(net156),
    .B2(\axi_controller.result_out[15] ),
    .X(_0579_));
 sky130_fd_sc_hd__a22o_1 _4329_ (.A1(net117),
    .A2(net192),
    .B1(net156),
    .B2(\axi_controller.result_out[14] ),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _4330_ (.A1(net116),
    .A2(net192),
    .B1(net156),
    .B2(\axi_controller.result_out[13] ),
    .X(_0581_));
 sky130_fd_sc_hd__a22o_1 _4331_ (.A1(net115),
    .A2(net192),
    .B1(net156),
    .B2(\axi_controller.result_out[12] ),
    .X(_0582_));
 sky130_fd_sc_hd__a22o_1 _4332_ (.A1(net114),
    .A2(net191),
    .B1(net156),
    .B2(\axi_controller.result_out[11] ),
    .X(_0583_));
 sky130_fd_sc_hd__a22o_1 _4333_ (.A1(net113),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[10] ),
    .X(_0584_));
 sky130_fd_sc_hd__a22o_1 _4334_ (.A1(net143),
    .A2(net192),
    .B1(net155),
    .B2(\axi_controller.result_out[9] ),
    .X(_0585_));
 sky130_fd_sc_hd__a22o_1 _4335_ (.A1(net142),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[8] ),
    .X(_0586_));
 sky130_fd_sc_hd__a22o_1 _4336_ (.A1(net141),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[7] ),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _4337_ (.A1(net140),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[6] ),
    .X(_0588_));
 sky130_fd_sc_hd__a22o_1 _4338_ (.A1(net139),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[5] ),
    .X(_0589_));
 sky130_fd_sc_hd__a22o_1 _4339_ (.A1(net138),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[4] ),
    .X(_0590_));
 sky130_fd_sc_hd__a22o_1 _4340_ (.A1(net137),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[3] ),
    .X(_0591_));
 sky130_fd_sc_hd__a22o_1 _4341_ (.A1(net134),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[2] ),
    .X(_0592_));
 sky130_fd_sc_hd__a22o_1 _4342_ (.A1(net123),
    .A2(net191),
    .B1(net155),
    .B2(\axi_controller.result_out[1] ),
    .X(_0593_));
 sky130_fd_sc_hd__a22o_1 _4343_ (.A1(\axi_controller.reg_done_flag ),
    .A2(_1990_),
    .B1(_2254_),
    .B2(\axi_controller.result_out[0] ),
    .X(_2257_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(_2257_),
    .A1(net112),
    .S(net194),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_1 _4345_ (.A(\cordic_inst.deg_handler_inst.theta_abs[31] ),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_1 _4346_ (.A(net255),
    .X(_0008_));
 sky130_fd_sc_hd__inv_2 _4347_ (.A(net318),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _4348_ (.A(net318),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _4349_ (.A(net321),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _4350_ (.A(net321),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _4351_ (.A(net321),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _4352_ (.A(net323),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _4353_ (.A(net323),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _4354_ (.A(net322),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _4355_ (.A(net323),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _4356_ (.A(net318),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _4357_ (.A(net322),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _4358_ (.A(net329),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _4359_ (.A(net329),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _4360_ (.A(net329),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _4361_ (.A(net329),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _4362_ (.A(net335),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _4363_ (.A(net334),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _4364_ (.A(net334),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _4365_ (.A(net336),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _4366_ (.A(net336),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _4367_ (.A(net334),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _4368_ (.A(net338),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _4369_ (.A(net337),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _4370_ (.A(net337),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _4371_ (.A(net341),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _4372_ (.A(net341),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _4373_ (.A(net342),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _4374_ (.A(net341),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _4375_ (.A(net341),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _4376_ (.A(net340),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _4377_ (.A(net340),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _4378_ (.A(net340),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _4379_ (.A(net332),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _4380_ (.A(net331),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _4381_ (.A(net331),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _4382_ (.A(net326),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(net326),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _4384_ (.A(net324),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _4385_ (.A(net324),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _4386_ (.A(net324),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _4387_ (.A(net324),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _4388_ (.A(net324),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _4389_ (.A(net324),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _4390_ (.A(net317),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _4391_ (.A(net317),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _4392_ (.A(net317),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _4393_ (.A(net317),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _4394_ (.A(net317),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _4395_ (.A(net319),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _4396_ (.A(net319),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _4397_ (.A(net319),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _4398_ (.A(net320),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _4399_ (.A(net317),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _4400_ (.A(net320),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _4401_ (.A(net320),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _4402_ (.A(net320),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _4403_ (.A(net320),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _4404_ (.A(net320),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _4405_ (.A(net320),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _4406_ (.A(net320),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _4407_ (.A(net320),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _4408_ (.A(net320),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _4409_ (.A(net321),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _4410_ (.A(net328),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _4411_ (.A(net328),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _4412_ (.A(net321),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _4413_ (.A(net321),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _4414_ (.A(net321),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _4415_ (.A(net321),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _4416_ (.A(net321),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _4417_ (.A(net322),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _4418_ (.A(net322),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _4419_ (.A(net323),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _4420_ (.A(net322),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _4421_ (.A(net322),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _4422_ (.A(net329),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _4423_ (.A(net330),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _4424_ (.A(net330),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _4425_ (.A(net329),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _4426_ (.A(net334),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _4427_ (.A(net334),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _4428_ (.A(net334),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _4429_ (.A(net336),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _4430_ (.A(net336),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _4431_ (.A(net337),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _4432_ (.A(net337),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _4433_ (.A(net337),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _4434_ (.A(net337),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _4435_ (.A(net338),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _4436_ (.A(net341),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _4437_ (.A(net341),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _4438_ (.A(net343),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _4439_ (.A(net343),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _4440_ (.A(net340),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _4441_ (.A(net333),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _4442_ (.A(net333),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _4443_ (.A(net333),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _4444_ (.A(net331),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _4445_ (.A(net331),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _4446_ (.A(net327),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _4447_ (.A(net326),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _4448_ (.A(net326),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _4449_ (.A(net325),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _4450_ (.A(net325),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _4451_ (.A(net326),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _4452_ (.A(net325),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _4453_ (.A(net324),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _4454_ (.A(net323),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _4455_ (.A(net322),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _4456_ (.A(net323),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _4457_ (.A(net322),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _4458_ (.A(net329),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _4459_ (.A(net329),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _4460_ (.A(net329),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _4461_ (.A(net334),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _4462_ (.A(net334),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _4463_ (.A(net335),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _4464_ (.A(net335),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _4465_ (.A(net337),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _4466_ (.A(net337),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _4467_ (.A(net337),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _4468_ (.A(net335),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _4469_ (.A(net338),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _4470_ (.A(net340),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _4471_ (.A(net340),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _4472_ (.A(net344),
    .Y(_0211_));
 sky130_fd_sc_hd__inv_2 _4473_ (.A(net344),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _4474_ (.A(net332),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _4475_ (.A(net332),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _4476_ (.A(net331),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _4477_ (.A(net331),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _4478_ (.A(net327),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_2 _4479_ (.A(net327),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _4480_ (.A(net325),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _4481_ (.A(net324),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _4482_ (.A(net324),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _4483_ (.A(net317),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _4484_ (.A(net324),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _4485_ (.A(net321),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _4486_ (.A(net322),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _4487_ (.A(net329),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _4488_ (.A(net330),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _4489_ (.A(net330),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _4490_ (.A(net330),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_2 _4491_ (.A(net334),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_2 _4492_ (.A(net334),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_2 _4493_ (.A(net335),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _4494_ (.A(net338),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _4495_ (.A(net338),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _4496_ (.A(net337),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _4497_ (.A(net341),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _4498_ (.A(net341),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _4499_ (.A(net341),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _4500_ (.A(net342),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_2 _4501_ (.A(net341),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _4502_ (.A(net340),
    .Y(_0241_));
 sky130_fd_sc_hd__inv_2 _4503_ (.A(net340),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _4504_ (.A(net345),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_2 _4505_ (.A(net333),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _4506_ (.A(net333),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _4507_ (.A(net333),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _4508_ (.A(net332),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_2 _4509_ (.A(net332),
    .Y(_0248_));
 sky130_fd_sc_hd__inv_2 _4510_ (.A(net331),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_2 _4511_ (.A(net331),
    .Y(_0250_));
 sky130_fd_sc_hd__inv_2 _4512_ (.A(net327),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _4513_ (.A(net327),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _4514_ (.A(net326),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _4515_ (.A(net326),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _4516_ (.A(net328),
    .Y(_0255_));
 sky130_fd_sc_hd__inv_2 _4517_ (.A(net325),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _4518_ (.A(net318),
    .Y(_0257_));
 sky130_fd_sc_hd__dfstp_1 _4519_ (.CLK(net380),
    .D(_0006_),
    .SET_B(_0085_),
    .Q(\cordic_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4520_ (.CLK(net380),
    .D(_0007_),
    .RESET_B(_0086_),
    .Q(\cordic_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4521_ (.CLK(net380),
    .D(_0000_),
    .RESET_B(_0087_),
    .Q(\cordic_inst.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(net370),
    .D(_0001_),
    .Q(\axi_controller.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(net370),
    .D(_0002_),
    .Q(\axi_controller.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(net368),
    .D(_0003_),
    .Q(\axi_controller.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(net368),
    .D(_0004_),
    .Q(\axi_controller.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(net352),
    .D(_0258_),
    .Q(\axi_controller.reg_input_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(net352),
    .D(_0259_),
    .Q(\axi_controller.reg_input_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(net353),
    .D(_0260_),
    .Q(\axi_controller.reg_input_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(net353),
    .D(_0261_),
    .Q(\axi_controller.reg_input_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(net353),
    .D(_0262_),
    .Q(\axi_controller.reg_input_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(net353),
    .D(_0263_),
    .Q(\axi_controller.reg_input_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(net353),
    .D(_0264_),
    .Q(\axi_controller.reg_input_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(net357),
    .D(_0265_),
    .Q(\axi_controller.reg_input_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(net362),
    .D(_0266_),
    .Q(\axi_controller.read_addr_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(net362),
    .D(_0267_),
    .Q(\axi_controller.read_addr_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(net351),
    .D(_0268_),
    .Q(\axi_controller.read_addr_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(net362),
    .D(_0269_),
    .Q(\axi_controller.read_addr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(net362),
    .D(_0270_),
    .Q(\axi_controller.read_addr_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(net362),
    .D(_0271_),
    .Q(\axi_controller.read_addr_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(net364),
    .D(_0272_),
    .Q(\axi_controller.read_addr_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(net364),
    .D(_0273_),
    .Q(\axi_controller.read_addr_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(net351),
    .D(_0274_),
    .Q(\axi_controller.read_addr_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(net351),
    .D(_0275_),
    .Q(\axi_controller.read_addr_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(net355),
    .D(_0276_),
    .Q(\axi_controller.read_addr_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(net354),
    .D(_0277_),
    .Q(\axi_controller.read_addr_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(net362),
    .D(_0278_),
    .Q(\axi_controller.read_addr_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(net351),
    .D(_0279_),
    .Q(\axi_controller.read_addr_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(net355),
    .D(_0280_),
    .Q(\axi_controller.read_addr_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(net355),
    .D(_0281_),
    .Q(\axi_controller.read_addr_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(net362),
    .D(_0282_),
    .Q(\axi_controller.read_addr_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(net362),
    .D(_0283_),
    .Q(\axi_controller.read_addr_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(net355),
    .D(_0284_),
    .Q(\axi_controller.read_addr_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(net364),
    .D(_0285_),
    .Q(\axi_controller.read_addr_reg[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(net355),
    .D(_0286_),
    .Q(\axi_controller.read_addr_reg[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(net355),
    .D(_0287_),
    .Q(\axi_controller.read_addr_reg[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(net355),
    .D(_0288_),
    .Q(\axi_controller.read_addr_reg[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(net362),
    .D(_0289_),
    .Q(\axi_controller.read_addr_reg[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(net354),
    .D(_0290_),
    .Q(\axi_controller.read_addr_reg[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(net355),
    .D(_0291_),
    .Q(\axi_controller.read_addr_reg[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(net355),
    .D(_0292_),
    .Q(\axi_controller.read_addr_reg[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(net354),
    .D(_0293_),
    .Q(\axi_controller.read_addr_reg[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(net362),
    .D(_0294_),
    .Q(\axi_controller.read_addr_reg[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(net351),
    .D(_0295_),
    .Q(\axi_controller.read_addr_reg[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(net351),
    .D(_0296_),
    .Q(\axi_controller.read_addr_reg[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(net355),
    .D(_0297_),
    .Q(\axi_controller.read_addr_reg[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(net370),
    .D(_0298_),
    .Q(\axi_controller.reg_done_flag ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(net364),
    .D(_0299_),
    .Q(\axi_controller.write_addr_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(net364),
    .D(_0300_),
    .Q(\axi_controller.write_addr_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(net364),
    .D(_0301_),
    .Q(\axi_controller.write_addr_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(net370),
    .D(_0302_),
    .Q(\axi_controller.write_addr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(net369),
    .D(_0303_),
    .Q(\axi_controller.write_addr_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(net369),
    .D(_0304_),
    .Q(\axi_controller.write_addr_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(net364),
    .D(_0305_),
    .Q(\axi_controller.write_addr_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(net364),
    .D(_0306_),
    .Q(\axi_controller.write_addr_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(net363),
    .D(_0307_),
    .Q(\axi_controller.write_addr_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(net364),
    .D(_0308_),
    .Q(\axi_controller.write_addr_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(net363),
    .D(_0309_),
    .Q(\axi_controller.write_addr_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(net363),
    .D(_0310_),
    .Q(\axi_controller.write_addr_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(net369),
    .D(_0311_),
    .Q(\axi_controller.write_addr_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(net363),
    .D(_0312_),
    .Q(\axi_controller.write_addr_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(net363),
    .D(_0313_),
    .Q(\axi_controller.write_addr_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(net369),
    .D(_0314_),
    .Q(\axi_controller.write_addr_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(net380),
    .D(_0315_),
    .Q(\axi_controller.write_addr_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(net370),
    .D(_0316_),
    .Q(\axi_controller.write_addr_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(net380),
    .D(_0317_),
    .Q(\axi_controller.write_addr_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(net380),
    .D(_0318_),
    .Q(\axi_controller.write_addr_reg[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(net380),
    .D(_0319_),
    .Q(\axi_controller.write_addr_reg[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(net380),
    .D(_0320_),
    .Q(\axi_controller.write_addr_reg[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(net382),
    .D(_0321_),
    .Q(\axi_controller.write_addr_reg[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(net382),
    .D(_0322_),
    .Q(\axi_controller.write_addr_reg[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(net385),
    .D(_0323_),
    .Q(\axi_controller.write_addr_reg[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(net381),
    .D(_0324_),
    .Q(\axi_controller.write_addr_reg[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(net381),
    .D(_0325_),
    .Q(\axi_controller.write_addr_reg[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(net385),
    .D(_0326_),
    .Q(\axi_controller.write_addr_reg[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(net381),
    .D(_0327_),
    .Q(\axi_controller.write_addr_reg[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(net381),
    .D(_0328_),
    .Q(\axi_controller.write_addr_reg[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(net382),
    .D(_0329_),
    .Q(\axi_controller.write_addr_reg[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(net385),
    .D(_0330_),
    .Q(\axi_controller.write_addr_reg[31] ));
 sky130_fd_sc_hd__dfxtp_2 _4599_ (.CLK(net369),
    .D(_0331_),
    .Q(\axi_controller.rst ));
 sky130_fd_sc_hd__dfxtp_2 _4600_ (.CLK(net365),
    .D(_0332_),
    .Q(\axi_controller.mode ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(net370),
    .D(_0333_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(net370),
    .D(_0334_),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_1 _4603_ (.CLK(net382),
    .D(_0335_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(net370),
    .D(_0336_),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(net371),
    .D(_0337_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(net352),
    .D(_0338_),
    .Q(\axi_controller.reg_input_data[24] ));
 sky130_fd_sc_hd__dfxtp_2 _4607_ (.CLK(net352),
    .D(_0339_),
    .Q(\axi_controller.reg_input_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(net351),
    .D(_0340_),
    .Q(\axi_controller.reg_input_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(net357),
    .D(_0341_),
    .Q(\axi_controller.reg_input_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(net357),
    .D(_0342_),
    .Q(\axi_controller.reg_input_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(net352),
    .D(_0343_),
    .Q(\axi_controller.reg_input_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(net352),
    .D(_0344_),
    .Q(\axi_controller.reg_input_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(net351),
    .D(_0345_),
    .Q(\axi_controller.reg_input_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(net381),
    .D(_0005_),
    .Q(\cordic_inst.deg_handler_inst.kuadran[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(net368),
    .D(_0346_),
    .Q(\axi_controller.reg_input_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(net368),
    .D(_0347_),
    .Q(\axi_controller.reg_input_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(net368),
    .D(_0348_),
    .Q(\axi_controller.reg_input_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(net363),
    .D(_0349_),
    .Q(\axi_controller.reg_input_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4619_ (.CLK(net363),
    .D(_0350_),
    .Q(\axi_controller.reg_input_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4620_ (.CLK(net363),
    .D(_0351_),
    .Q(\axi_controller.reg_input_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(net363),
    .D(_0352_),
    .Q(\axi_controller.reg_input_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(net363),
    .D(_0353_),
    .Q(\axi_controller.reg_input_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4623_ (.CLK(net381),
    .D(_0354_),
    .RESET_B(net317),
    .Q(\axi_controller.result_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4624_ (.CLK(net399),
    .D(_0355_),
    .RESET_B(net336),
    .Q(\axi_controller.result_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4625_ (.CLK(net398),
    .D(_0356_),
    .RESET_B(net339),
    .Q(\axi_controller.result_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4626_ (.CLK(net398),
    .D(_0357_),
    .RESET_B(net339),
    .Q(\axi_controller.result_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4627_ (.CLK(net399),
    .D(_0358_),
    .RESET_B(net336),
    .Q(\axi_controller.result_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4628_ (.CLK(net398),
    .D(_0359_),
    .RESET_B(net336),
    .Q(\axi_controller.result_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4629_ (.CLK(net398),
    .D(_0360_),
    .RESET_B(net336),
    .Q(\axi_controller.result_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4630_ (.CLK(net398),
    .D(_0361_),
    .RESET_B(net336),
    .Q(\axi_controller.result_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4631_ (.CLK(net398),
    .D(_0362_),
    .RESET_B(net336),
    .Q(\axi_controller.result_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4632_ (.CLK(net401),
    .D(_0363_),
    .RESET_B(net338),
    .Q(\axi_controller.result_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4633_ (.CLK(net401),
    .D(_0364_),
    .RESET_B(net338),
    .Q(\axi_controller.result_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4634_ (.CLK(net401),
    .D(_0365_),
    .RESET_B(net338),
    .Q(\axi_controller.result_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4635_ (.CLK(net401),
    .D(_0366_),
    .RESET_B(net338),
    .Q(\axi_controller.result_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4636_ (.CLK(net406),
    .D(_0367_),
    .RESET_B(net342),
    .Q(\axi_controller.result_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4637_ (.CLK(net406),
    .D(_0368_),
    .RESET_B(net342),
    .Q(\axi_controller.result_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4638_ (.CLK(net406),
    .D(_0369_),
    .RESET_B(net342),
    .Q(\axi_controller.result_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4639_ (.CLK(net407),
    .D(_0370_),
    .RESET_B(net343),
    .Q(\axi_controller.result_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4640_ (.CLK(net407),
    .D(_0371_),
    .RESET_B(net343),
    .Q(\axi_controller.result_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4641_ (.CLK(net403),
    .D(_0372_),
    .RESET_B(net340),
    .Q(\axi_controller.result_out[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4642_ (.CLK(net403),
    .D(_0373_),
    .RESET_B(net340),
    .Q(\axi_controller.result_out[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4643_ (.CLK(net394),
    .D(_0374_),
    .RESET_B(net333),
    .Q(\axi_controller.result_out[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4644_ (.CLK(net394),
    .D(_0375_),
    .RESET_B(net333),
    .Q(\axi_controller.result_out[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4645_ (.CLK(net394),
    .D(_0376_),
    .RESET_B(net331),
    .Q(\axi_controller.result_out[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4646_ (.CLK(net392),
    .D(_0377_),
    .RESET_B(net331),
    .Q(\axi_controller.result_out[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4647_ (.CLK(net393),
    .D(_0378_),
    .RESET_B(net326),
    .Q(\axi_controller.result_out[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4648_ (.CLK(net393),
    .D(_0379_),
    .RESET_B(net326),
    .Q(\axi_controller.result_out[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4649_ (.CLK(net384),
    .D(_0380_),
    .RESET_B(net326),
    .Q(\axi_controller.result_out[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4650_ (.CLK(net384),
    .D(_0381_),
    .RESET_B(net325),
    .Q(\axi_controller.result_out[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4651_ (.CLK(net385),
    .D(_0382_),
    .RESET_B(net325),
    .Q(\axi_controller.result_out[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4652_ (.CLK(net385),
    .D(_0383_),
    .RESET_B(net325),
    .Q(\axi_controller.result_out[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4653_ (.CLK(net381),
    .D(_0384_),
    .RESET_B(net317),
    .Q(\axi_controller.result_out[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4654_ (.CLK(net382),
    .D(_0385_),
    .RESET_B(net325),
    .Q(\axi_controller.result_out[31] ));
 sky130_fd_sc_hd__dfrtp_1 _4655_ (.CLK(net381),
    .D(net200),
    .RESET_B(net317),
    .Q(\axi_controller.done ));
 sky130_fd_sc_hd__dfrtp_1 _4656_ (.CLK(net377),
    .D(_0386_),
    .RESET_B(_0088_),
    .Q(\cordic_inst.cordic_inst.i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4657_ (.CLK(net377),
    .D(_0387_),
    .RESET_B(_0089_),
    .Q(\cordic_inst.cordic_inst.i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4658_ (.CLK(net377),
    .D(_0388_),
    .RESET_B(_0090_),
    .Q(\cordic_inst.cordic_inst.i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4659_ (.CLK(net377),
    .D(_0389_),
    .RESET_B(_0091_),
    .Q(\cordic_inst.cordic_inst.i[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4660_ (.CLK(net377),
    .D(_0390_),
    .RESET_B(_0092_),
    .Q(\cordic_inst.cordic_inst.i[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4661_ (.CLK(net389),
    .D(\cordic_inst.cordic_inst.done ),
    .RESET_B(net322),
    .Q(\cordic_inst.sign_handler_inst.done_d ));
 sky130_fd_sc_hd__dfxtp_1 _4662_ (.CLK(net352),
    .D(_0391_),
    .Q(\axi_controller.reg_input_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(net352),
    .D(_0392_),
    .Q(\axi_controller.reg_input_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4664_ (.CLK(net352),
    .D(_0393_),
    .Q(\axi_controller.reg_input_data[18] ));
 sky130_fd_sc_hd__dfxtp_2 _4665_ (.CLK(net352),
    .D(_0394_),
    .Q(\axi_controller.reg_input_data[19] ));
 sky130_fd_sc_hd__dfxtp_2 _4666_ (.CLK(net351),
    .D(_0395_),
    .Q(\axi_controller.reg_input_data[20] ));
 sky130_fd_sc_hd__dfxtp_2 _4667_ (.CLK(net357),
    .D(_0396_),
    .Q(\axi_controller.reg_input_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4668_ (.CLK(net357),
    .D(_0397_),
    .Q(\axi_controller.reg_input_data[22] ));
 sky130_fd_sc_hd__dfxtp_2 _4669_ (.CLK(net351),
    .D(_0398_),
    .Q(\axi_controller.reg_input_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4670_ (.CLK(net371),
    .D(_0399_),
    .Q(net144));
 sky130_fd_sc_hd__dfrtp_1 _4671_ (.CLK(net375),
    .D(\cordic_inst.cordic_inst.next_state[0] ),
    .RESET_B(_0093_),
    .Q(\cordic_inst.cordic_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4672_ (.CLK(net377),
    .D(net158),
    .RESET_B(_0094_),
    .Q(\cordic_inst.cordic_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4673_ (.CLK(net381),
    .D(_0400_),
    .RESET_B(_0095_),
    .Q(\cordic_inst.cordic_inst.start ));
 sky130_fd_sc_hd__dfrtp_1 _4674_ (.CLK(net375),
    .D(_0401_),
    .RESET_B(_0096_),
    .Q(\cordic_inst.cordic_inst.done ));
 sky130_fd_sc_hd__dfrtp_1 _4675_ (.CLK(net389),
    .D(_0402_),
    .RESET_B(_0097_),
    .Q(\cordic_inst.cordic_inst.cos_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4676_ (.CLK(net391),
    .D(_0403_),
    .RESET_B(_0098_),
    .Q(\cordic_inst.cordic_inst.cos_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4677_ (.CLK(net389),
    .D(_0404_),
    .RESET_B(_0099_),
    .Q(\cordic_inst.cordic_inst.cos_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4678_ (.CLK(net389),
    .D(_0405_),
    .RESET_B(_0100_),
    .Q(\cordic_inst.cordic_inst.cos_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4679_ (.CLK(net396),
    .D(_0406_),
    .RESET_B(_0101_),
    .Q(\cordic_inst.cordic_inst.cos_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4680_ (.CLK(net396),
    .D(_0407_),
    .RESET_B(_0102_),
    .Q(\cordic_inst.cordic_inst.cos_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4681_ (.CLK(net399),
    .D(_0408_),
    .RESET_B(_0103_),
    .Q(\cordic_inst.cordic_inst.cos_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4682_ (.CLK(net399),
    .D(_0409_),
    .RESET_B(_0104_),
    .Q(\cordic_inst.cordic_inst.cos_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4683_ (.CLK(net399),
    .D(_0410_),
    .RESET_B(_0105_),
    .Q(\cordic_inst.cordic_inst.cos_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4684_ (.CLK(net396),
    .D(_0411_),
    .RESET_B(_0106_),
    .Q(\cordic_inst.cordic_inst.cos_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4685_ (.CLK(net401),
    .D(_0412_),
    .RESET_B(_0107_),
    .Q(\cordic_inst.cordic_inst.cos_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4686_ (.CLK(net400),
    .D(_0413_),
    .RESET_B(_0108_),
    .Q(\cordic_inst.cordic_inst.cos_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4687_ (.CLK(net400),
    .D(_0414_),
    .RESET_B(_0109_),
    .Q(\cordic_inst.cordic_inst.cos_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4688_ (.CLK(net405),
    .D(_0415_),
    .RESET_B(_0110_),
    .Q(\cordic_inst.cordic_inst.cos_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4689_ (.CLK(net405),
    .D(_0416_),
    .RESET_B(_0111_),
    .Q(\cordic_inst.cordic_inst.cos_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4690_ (.CLK(net405),
    .D(_0417_),
    .RESET_B(_0112_),
    .Q(\cordic_inst.cordic_inst.cos_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4691_ (.CLK(net405),
    .D(_0418_),
    .RESET_B(_0113_),
    .Q(\cordic_inst.cordic_inst.cos_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4692_ (.CLK(net405),
    .D(_0419_),
    .RESET_B(_0114_),
    .Q(\cordic_inst.cordic_inst.cos_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4693_ (.CLK(net404),
    .D(_0420_),
    .RESET_B(_0115_),
    .Q(\cordic_inst.cordic_inst.cos_out[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4694_ (.CLK(net403),
    .D(_0421_),
    .RESET_B(_0116_),
    .Q(\cordic_inst.cordic_inst.cos_out[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4695_ (.CLK(net403),
    .D(_0422_),
    .RESET_B(_0117_),
    .Q(\cordic_inst.cordic_inst.cos_out[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4696_ (.CLK(net394),
    .D(_0423_),
    .RESET_B(_0118_),
    .Q(\cordic_inst.cordic_inst.cos_out[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4697_ (.CLK(net392),
    .D(_0424_),
    .RESET_B(_0119_),
    .Q(\cordic_inst.cordic_inst.cos_out[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4698_ (.CLK(net392),
    .D(_0425_),
    .RESET_B(_0120_),
    .Q(\cordic_inst.cordic_inst.cos_out[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4699_ (.CLK(net393),
    .D(_0426_),
    .RESET_B(_0121_),
    .Q(\cordic_inst.cordic_inst.cos_out[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4700_ (.CLK(net384),
    .D(_0427_),
    .RESET_B(_0122_),
    .Q(\cordic_inst.cordic_inst.cos_out[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4701_ (.CLK(net386),
    .D(_0428_),
    .RESET_B(_0123_),
    .Q(\cordic_inst.cordic_inst.cos_out[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4702_ (.CLK(net386),
    .D(_0429_),
    .RESET_B(_0124_),
    .Q(\cordic_inst.cordic_inst.cos_out[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4703_ (.CLK(net386),
    .D(_0430_),
    .RESET_B(_0125_),
    .Q(\cordic_inst.cordic_inst.cos_out[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4704_ (.CLK(net386),
    .D(_0431_),
    .RESET_B(_0126_),
    .Q(\cordic_inst.cordic_inst.cos_out[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4705_ (.CLK(net379),
    .D(_0432_),
    .RESET_B(_0127_),
    .Q(\cordic_inst.cordic_inst.cos_out[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4706_ (.CLK(net379),
    .D(_0433_),
    .RESET_B(_0128_),
    .Q(\cordic_inst.cordic_inst.cos_out[31] ));
 sky130_fd_sc_hd__dfrtp_1 _4707_ (.CLK(net379),
    .D(_0434_),
    .RESET_B(_0129_),
    .Q(\cordic_inst.cordic_inst.z[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4708_ (.CLK(net379),
    .D(_0435_),
    .RESET_B(_0130_),
    .Q(\cordic_inst.cordic_inst.z[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4709_ (.CLK(net379),
    .D(_0436_),
    .RESET_B(_0131_),
    .Q(\cordic_inst.cordic_inst.z[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4710_ (.CLK(net379),
    .D(_0437_),
    .RESET_B(_0132_),
    .Q(\cordic_inst.cordic_inst.z[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4711_ (.CLK(net379),
    .D(_0438_),
    .RESET_B(_0133_),
    .Q(\cordic_inst.cordic_inst.z[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4712_ (.CLK(net367),
    .D(_0439_),
    .RESET_B(_0134_),
    .Q(\cordic_inst.cordic_inst.z[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4713_ (.CLK(net367),
    .D(_0440_),
    .RESET_B(_0135_),
    .Q(\cordic_inst.cordic_inst.z[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4714_ (.CLK(net366),
    .D(_0441_),
    .RESET_B(_0136_),
    .Q(\cordic_inst.cordic_inst.z[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4715_ (.CLK(net367),
    .D(_0442_),
    .RESET_B(_0137_),
    .Q(\cordic_inst.cordic_inst.z[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4716_ (.CLK(net367),
    .D(_0443_),
    .RESET_B(_0138_),
    .Q(\cordic_inst.cordic_inst.z[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4717_ (.CLK(net359),
    .D(_0444_),
    .RESET_B(_0139_),
    .Q(\cordic_inst.cordic_inst.z[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4718_ (.CLK(net360),
    .D(_0445_),
    .RESET_B(_0140_),
    .Q(\cordic_inst.cordic_inst.z[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4719_ (.CLK(net360),
    .D(_0446_),
    .RESET_B(_0141_),
    .Q(\cordic_inst.cordic_inst.z[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4720_ (.CLK(net360),
    .D(_0447_),
    .RESET_B(_0142_),
    .Q(\cordic_inst.cordic_inst.z[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4721_ (.CLK(net360),
    .D(_0448_),
    .RESET_B(_0143_),
    .Q(\cordic_inst.cordic_inst.z[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4722_ (.CLK(net360),
    .D(_0449_),
    .RESET_B(_0144_),
    .Q(\cordic_inst.cordic_inst.z[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4723_ (.CLK(net374),
    .D(_0450_),
    .RESET_B(_0145_),
    .Q(\cordic_inst.cordic_inst.z[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4724_ (.CLK(net374),
    .D(_0451_),
    .RESET_B(_0146_),
    .Q(\cordic_inst.cordic_inst.z[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4725_ (.CLK(net374),
    .D(_0452_),
    .RESET_B(_0147_),
    .Q(\cordic_inst.cordic_inst.z[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4726_ (.CLK(net377),
    .D(_0453_),
    .RESET_B(_0148_),
    .Q(\cordic_inst.cordic_inst.z[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4727_ (.CLK(net377),
    .D(_0454_),
    .RESET_B(_0149_),
    .Q(\cordic_inst.cordic_inst.z[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4728_ (.CLK(net378),
    .D(_0455_),
    .RESET_B(_0150_),
    .Q(\cordic_inst.cordic_inst.z[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4729_ (.CLK(net375),
    .D(_0456_),
    .RESET_B(_0151_),
    .Q(\cordic_inst.cordic_inst.z[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4730_ (.CLK(net376),
    .D(_0457_),
    .RESET_B(_0152_),
    .Q(\cordic_inst.cordic_inst.z[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4731_ (.CLK(net372),
    .D(_0458_),
    .RESET_B(_0153_),
    .Q(\cordic_inst.cordic_inst.z[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4732_ (.CLK(net375),
    .D(_0459_),
    .RESET_B(_0154_),
    .Q(\cordic_inst.cordic_inst.z[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4733_ (.CLK(net375),
    .D(_0460_),
    .RESET_B(_0155_),
    .Q(\cordic_inst.cordic_inst.z[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4734_ (.CLK(net376),
    .D(_0461_),
    .RESET_B(_0156_),
    .Q(\cordic_inst.cordic_inst.z[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4735_ (.CLK(net376),
    .D(_0462_),
    .RESET_B(_0157_),
    .Q(\cordic_inst.cordic_inst.z[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4736_ (.CLK(net389),
    .D(_0463_),
    .RESET_B(_0158_),
    .Q(\cordic_inst.cordic_inst.z[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4737_ (.CLK(net376),
    .D(_0464_),
    .RESET_B(_0159_),
    .Q(\cordic_inst.cordic_inst.z[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4738_ (.CLK(net389),
    .D(_0465_),
    .RESET_B(_0160_),
    .Q(\cordic_inst.cordic_inst.z[31] ));
 sky130_fd_sc_hd__dfrtp_2 _4739_ (.CLK(net390),
    .D(_0466_),
    .RESET_B(_0161_),
    .Q(\cordic_inst.cordic_inst.sin_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _4740_ (.CLK(net391),
    .D(_0467_),
    .RESET_B(_0162_),
    .Q(\cordic_inst.cordic_inst.sin_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _4741_ (.CLK(net391),
    .D(_0468_),
    .RESET_B(_0163_),
    .Q(\cordic_inst.cordic_inst.sin_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4742_ (.CLK(net391),
    .D(_0469_),
    .RESET_B(_0164_),
    .Q(\cordic_inst.cordic_inst.sin_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _4743_ (.CLK(net396),
    .D(_0470_),
    .RESET_B(_0165_),
    .Q(\cordic_inst.cordic_inst.sin_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _4744_ (.CLK(net396),
    .D(_0471_),
    .RESET_B(_0166_),
    .Q(\cordic_inst.cordic_inst.sin_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _4745_ (.CLK(net396),
    .D(_0472_),
    .RESET_B(_0167_),
    .Q(\cordic_inst.cordic_inst.sin_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _4746_ (.CLK(net399),
    .D(_0473_),
    .RESET_B(_0168_),
    .Q(\cordic_inst.cordic_inst.sin_out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _4747_ (.CLK(net400),
    .D(_0474_),
    .RESET_B(_0169_),
    .Q(\cordic_inst.cordic_inst.sin_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _4748_ (.CLK(net400),
    .D(_0475_),
    .RESET_B(_0170_),
    .Q(\cordic_inst.cordic_inst.sin_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _4749_ (.CLK(net400),
    .D(_0476_),
    .RESET_B(_0171_),
    .Q(\cordic_inst.cordic_inst.sin_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _4750_ (.CLK(net400),
    .D(_0477_),
    .RESET_B(_0172_),
    .Q(\cordic_inst.cordic_inst.sin_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _4751_ (.CLK(net400),
    .D(_0478_),
    .RESET_B(_0173_),
    .Q(\cordic_inst.cordic_inst.sin_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _4752_ (.CLK(net406),
    .D(_0479_),
    .RESET_B(_0174_),
    .Q(\cordic_inst.cordic_inst.sin_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _4753_ (.CLK(net405),
    .D(_0480_),
    .RESET_B(_0175_),
    .Q(\cordic_inst.cordic_inst.sin_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _4754_ (.CLK(net406),
    .D(_0481_),
    .RESET_B(_0176_),
    .Q(\cordic_inst.cordic_inst.sin_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _4755_ (.CLK(net407),
    .D(_0482_),
    .RESET_B(_0177_),
    .Q(\cordic_inst.cordic_inst.sin_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _4756_ (.CLK(net407),
    .D(_0483_),
    .RESET_B(_0178_),
    .Q(\cordic_inst.cordic_inst.sin_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _4757_ (.CLK(net404),
    .D(_0484_),
    .RESET_B(_0179_),
    .Q(\cordic_inst.cordic_inst.sin_out[18] ));
 sky130_fd_sc_hd__dfrtp_1 _4758_ (.CLK(net403),
    .D(_0485_),
    .RESET_B(_0180_),
    .Q(\cordic_inst.cordic_inst.sin_out[19] ));
 sky130_fd_sc_hd__dfrtp_1 _4759_ (.CLK(net394),
    .D(_0486_),
    .RESET_B(_0181_),
    .Q(\cordic_inst.cordic_inst.sin_out[20] ));
 sky130_fd_sc_hd__dfrtp_1 _4760_ (.CLK(net395),
    .D(_0487_),
    .RESET_B(_0182_),
    .Q(\cordic_inst.cordic_inst.sin_out[21] ));
 sky130_fd_sc_hd__dfrtp_1 _4761_ (.CLK(net394),
    .D(_0488_),
    .RESET_B(_0183_),
    .Q(\cordic_inst.cordic_inst.sin_out[22] ));
 sky130_fd_sc_hd__dfrtp_1 _4762_ (.CLK(net392),
    .D(_0489_),
    .RESET_B(_0184_),
    .Q(\cordic_inst.cordic_inst.sin_out[23] ));
 sky130_fd_sc_hd__dfrtp_1 _4763_ (.CLK(net393),
    .D(_0490_),
    .RESET_B(_0185_),
    .Q(\cordic_inst.cordic_inst.sin_out[24] ));
 sky130_fd_sc_hd__dfrtp_1 _4764_ (.CLK(net393),
    .D(_0491_),
    .RESET_B(_0186_),
    .Q(\cordic_inst.cordic_inst.sin_out[25] ));
 sky130_fd_sc_hd__dfrtp_1 _4765_ (.CLK(net384),
    .D(_0492_),
    .RESET_B(_0187_),
    .Q(\cordic_inst.cordic_inst.sin_out[26] ));
 sky130_fd_sc_hd__dfrtp_1 _4766_ (.CLK(net385),
    .D(_0493_),
    .RESET_B(_0188_),
    .Q(\cordic_inst.cordic_inst.sin_out[27] ));
 sky130_fd_sc_hd__dfrtp_1 _4767_ (.CLK(net385),
    .D(_0494_),
    .RESET_B(_0189_),
    .Q(\cordic_inst.cordic_inst.sin_out[28] ));
 sky130_fd_sc_hd__dfrtp_1 _4768_ (.CLK(net384),
    .D(_0495_),
    .RESET_B(_0190_),
    .Q(\cordic_inst.cordic_inst.sin_out[29] ));
 sky130_fd_sc_hd__dfrtp_1 _4769_ (.CLK(net384),
    .D(_0496_),
    .RESET_B(_0191_),
    .Q(\cordic_inst.cordic_inst.sin_out[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4770_ (.CLK(net381),
    .D(_0497_),
    .RESET_B(_0192_),
    .Q(\cordic_inst.cordic_inst.sin_out[31] ));
 sky130_fd_sc_hd__dfrtp_1 _4771_ (.CLK(net390),
    .D(_0498_),
    .RESET_B(_0193_),
    .Q(\cordic_inst.cordic_inst.x[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4772_ (.CLK(net390),
    .D(_0499_),
    .RESET_B(_0194_),
    .Q(\cordic_inst.cordic_inst.x[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4773_ (.CLK(net389),
    .D(_0500_),
    .RESET_B(_0195_),
    .Q(\cordic_inst.cordic_inst.x[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4774_ (.CLK(net389),
    .D(_0501_),
    .RESET_B(_0196_),
    .Q(\cordic_inst.cordic_inst.x[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4775_ (.CLK(net390),
    .D(_0502_),
    .RESET_B(_0197_),
    .Q(\cordic_inst.cordic_inst.x[4] ));
 sky130_fd_sc_hd__dfrtp_4 _4776_ (.CLK(net390),
    .D(_0503_),
    .RESET_B(_0198_),
    .Q(\cordic_inst.cordic_inst.x[5] ));
 sky130_fd_sc_hd__dfrtp_4 _4777_ (.CLK(net391),
    .D(_0504_),
    .RESET_B(_0199_),
    .Q(\cordic_inst.cordic_inst.x[6] ));
 sky130_fd_sc_hd__dfrtp_2 _4778_ (.CLK(net396),
    .D(_0505_),
    .RESET_B(_0200_),
    .Q(\cordic_inst.cordic_inst.x[7] ));
 sky130_fd_sc_hd__dfrtp_2 _4779_ (.CLK(net397),
    .D(_0506_),
    .RESET_B(_0201_),
    .Q(\cordic_inst.cordic_inst.x[8] ));
 sky130_fd_sc_hd__dfrtp_2 _4780_ (.CLK(net397),
    .D(_0507_),
    .RESET_B(_0202_),
    .Q(\cordic_inst.cordic_inst.x[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4781_ (.CLK(net400),
    .D(_0508_),
    .RESET_B(_0203_),
    .Q(\cordic_inst.cordic_inst.x[10] ));
 sky130_fd_sc_hd__dfrtp_2 _4782_ (.CLK(net400),
    .D(_0509_),
    .RESET_B(_0204_),
    .Q(\cordic_inst.cordic_inst.x[11] ));
 sky130_fd_sc_hd__dfrtp_4 _4783_ (.CLK(net400),
    .D(_0510_),
    .RESET_B(_0205_),
    .Q(\cordic_inst.cordic_inst.x[12] ));
 sky130_fd_sc_hd__dfrtp_4 _4784_ (.CLK(net401),
    .D(_0511_),
    .RESET_B(_0206_),
    .Q(\cordic_inst.cordic_inst.x[13] ));
 sky130_fd_sc_hd__dfrtp_4 _4785_ (.CLK(net397),
    .D(_0512_),
    .RESET_B(_0207_),
    .Q(\cordic_inst.cordic_inst.x[14] ));
 sky130_fd_sc_hd__dfrtp_4 _4786_ (.CLK(net401),
    .D(_0513_),
    .RESET_B(_0208_),
    .Q(\cordic_inst.cordic_inst.x[15] ));
 sky130_fd_sc_hd__dfrtp_4 _4787_ (.CLK(net404),
    .D(_0514_),
    .RESET_B(_0209_),
    .Q(\cordic_inst.cordic_inst.x[16] ));
 sky130_fd_sc_hd__dfrtp_2 _4788_ (.CLK(net404),
    .D(_0515_),
    .RESET_B(_0210_),
    .Q(\cordic_inst.cordic_inst.x[17] ));
 sky130_fd_sc_hd__dfrtp_4 _4789_ (.CLK(net404),
    .D(_0516_),
    .RESET_B(_0211_),
    .Q(\cordic_inst.cordic_inst.x[18] ));
 sky130_fd_sc_hd__dfrtp_2 _4790_ (.CLK(net403),
    .D(_0517_),
    .RESET_B(_0212_),
    .Q(\cordic_inst.cordic_inst.x[19] ));
 sky130_fd_sc_hd__dfrtp_4 _4791_ (.CLK(net394),
    .D(_0518_),
    .RESET_B(_0213_),
    .Q(\cordic_inst.cordic_inst.x[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4792_ (.CLK(net392),
    .D(_0519_),
    .RESET_B(_0214_),
    .Q(\cordic_inst.cordic_inst.x[21] ));
 sky130_fd_sc_hd__dfrtp_2 _4793_ (.CLK(net392),
    .D(_0520_),
    .RESET_B(_0215_),
    .Q(\cordic_inst.cordic_inst.x[22] ));
 sky130_fd_sc_hd__dfrtp_4 _4794_ (.CLK(net392),
    .D(_0521_),
    .RESET_B(_0216_),
    .Q(\cordic_inst.cordic_inst.x[23] ));
 sky130_fd_sc_hd__dfrtp_2 _4795_ (.CLK(net386),
    .D(_0522_),
    .RESET_B(_0217_),
    .Q(\cordic_inst.cordic_inst.x[24] ));
 sky130_fd_sc_hd__dfrtp_2 _4796_ (.CLK(net386),
    .D(_0523_),
    .RESET_B(_0218_),
    .Q(\cordic_inst.cordic_inst.x[25] ));
 sky130_fd_sc_hd__dfrtp_2 _4797_ (.CLK(net386),
    .D(_0524_),
    .RESET_B(_0219_),
    .Q(\cordic_inst.cordic_inst.x[26] ));
 sky130_fd_sc_hd__dfrtp_4 _4798_ (.CLK(net386),
    .D(_0525_),
    .RESET_B(_0220_),
    .Q(\cordic_inst.cordic_inst.x[27] ));
 sky130_fd_sc_hd__dfrtp_2 _4799_ (.CLK(net386),
    .D(_0526_),
    .RESET_B(_0221_),
    .Q(\cordic_inst.cordic_inst.x[28] ));
 sky130_fd_sc_hd__dfrtp_4 _4800_ (.CLK(net383),
    .D(_0527_),
    .RESET_B(_0222_),
    .Q(\cordic_inst.cordic_inst.x[29] ));
 sky130_fd_sc_hd__dfrtp_4 _4801_ (.CLK(net383),
    .D(_0528_),
    .RESET_B(_0223_),
    .Q(\cordic_inst.cordic_inst.x[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4802_ (.CLK(net383),
    .D(_0529_),
    .RESET_B(_0224_),
    .Q(\cordic_inst.cordic_inst.x[31] ));
 sky130_fd_sc_hd__dfrtp_1 _4803_ (.CLK(net389),
    .D(_0530_),
    .RESET_B(_0225_),
    .Q(\cordic_inst.cordic_inst.y[0] ));
 sky130_fd_sc_hd__dfrtp_2 _4804_ (.CLK(net391),
    .D(_0531_),
    .RESET_B(_0226_),
    .Q(\cordic_inst.cordic_inst.y[1] ));
 sky130_fd_sc_hd__dfrtp_2 _4805_ (.CLK(net391),
    .D(_0532_),
    .RESET_B(_0227_),
    .Q(\cordic_inst.cordic_inst.y[2] ));
 sky130_fd_sc_hd__dfrtp_1 _4806_ (.CLK(net391),
    .D(_0533_),
    .RESET_B(_0228_),
    .Q(\cordic_inst.cordic_inst.y[3] ));
 sky130_fd_sc_hd__dfrtp_4 _4807_ (.CLK(net396),
    .D(_0534_),
    .RESET_B(_0229_),
    .Q(\cordic_inst.cordic_inst.y[4] ));
 sky130_fd_sc_hd__dfrtp_2 _4808_ (.CLK(net396),
    .D(_0535_),
    .RESET_B(_0230_),
    .Q(\cordic_inst.cordic_inst.y[5] ));
 sky130_fd_sc_hd__dfrtp_2 _4809_ (.CLK(net396),
    .D(_0536_),
    .RESET_B(_0231_),
    .Q(\cordic_inst.cordic_inst.y[6] ));
 sky130_fd_sc_hd__dfrtp_4 _4810_ (.CLK(net397),
    .D(_0537_),
    .RESET_B(_0232_),
    .Q(\cordic_inst.cordic_inst.y[7] ));
 sky130_fd_sc_hd__dfrtp_4 _4811_ (.CLK(net401),
    .D(_0538_),
    .RESET_B(_0233_),
    .Q(\cordic_inst.cordic_inst.y[8] ));
 sky130_fd_sc_hd__dfrtp_4 _4812_ (.CLK(net401),
    .D(_0539_),
    .RESET_B(_0234_),
    .Q(\cordic_inst.cordic_inst.y[9] ));
 sky130_fd_sc_hd__dfrtp_2 _4813_ (.CLK(net405),
    .D(_0540_),
    .RESET_B(_0235_),
    .Q(\cordic_inst.cordic_inst.y[10] ));
 sky130_fd_sc_hd__dfrtp_2 _4814_ (.CLK(net405),
    .D(_0541_),
    .RESET_B(_0236_),
    .Q(\cordic_inst.cordic_inst.y[11] ));
 sky130_fd_sc_hd__dfrtp_2 _4815_ (.CLK(net405),
    .D(_0542_),
    .RESET_B(_0237_),
    .Q(\cordic_inst.cordic_inst.y[12] ));
 sky130_fd_sc_hd__dfrtp_4 _4816_ (.CLK(net405),
    .D(_0543_),
    .RESET_B(_0238_),
    .Q(\cordic_inst.cordic_inst.y[13] ));
 sky130_fd_sc_hd__dfrtp_4 _4817_ (.CLK(net406),
    .D(_0544_),
    .RESET_B(_0239_),
    .Q(\cordic_inst.cordic_inst.y[14] ));
 sky130_fd_sc_hd__dfrtp_4 _4818_ (.CLK(net406),
    .D(_0545_),
    .RESET_B(_0240_),
    .Q(\cordic_inst.cordic_inst.y[15] ));
 sky130_fd_sc_hd__dfrtp_2 _4819_ (.CLK(net403),
    .D(_0546_),
    .RESET_B(_0241_),
    .Q(\cordic_inst.cordic_inst.y[16] ));
 sky130_fd_sc_hd__dfrtp_4 _4820_ (.CLK(net404),
    .D(_0547_),
    .RESET_B(_0242_),
    .Q(\cordic_inst.cordic_inst.y[17] ));
 sky130_fd_sc_hd__dfrtp_4 _4821_ (.CLK(net403),
    .D(_0548_),
    .RESET_B(_0243_),
    .Q(\cordic_inst.cordic_inst.y[18] ));
 sky130_fd_sc_hd__dfrtp_4 _4822_ (.CLK(net395),
    .D(_0549_),
    .RESET_B(_0244_),
    .Q(\cordic_inst.cordic_inst.y[19] ));
 sky130_fd_sc_hd__dfrtp_4 _4823_ (.CLK(net395),
    .D(_0550_),
    .RESET_B(_0245_),
    .Q(\cordic_inst.cordic_inst.y[20] ));
 sky130_fd_sc_hd__dfrtp_2 _4824_ (.CLK(net395),
    .D(_0551_),
    .RESET_B(_0246_),
    .Q(\cordic_inst.cordic_inst.y[21] ));
 sky130_fd_sc_hd__dfrtp_2 _4825_ (.CLK(net394),
    .D(_0552_),
    .RESET_B(_0247_),
    .Q(\cordic_inst.cordic_inst.y[22] ));
 sky130_fd_sc_hd__dfrtp_4 _4826_ (.CLK(net394),
    .D(_0553_),
    .RESET_B(_0248_),
    .Q(\cordic_inst.cordic_inst.y[23] ));
 sky130_fd_sc_hd__dfrtp_4 _4827_ (.CLK(net392),
    .D(_0554_),
    .RESET_B(_0249_),
    .Q(\cordic_inst.cordic_inst.y[24] ));
 sky130_fd_sc_hd__dfrtp_4 _4828_ (.CLK(net392),
    .D(_0555_),
    .RESET_B(_0250_),
    .Q(\cordic_inst.cordic_inst.y[25] ));
 sky130_fd_sc_hd__dfrtp_4 _4829_ (.CLK(net393),
    .D(_0556_),
    .RESET_B(_0251_),
    .Q(\cordic_inst.cordic_inst.y[26] ));
 sky130_fd_sc_hd__dfrtp_4 _4830_ (.CLK(net393),
    .D(_0557_),
    .RESET_B(_0252_),
    .Q(\cordic_inst.cordic_inst.y[27] ));
 sky130_fd_sc_hd__dfrtp_4 _4831_ (.CLK(net384),
    .D(_0558_),
    .RESET_B(_0253_),
    .Q(\cordic_inst.cordic_inst.y[28] ));
 sky130_fd_sc_hd__dfrtp_4 _4832_ (.CLK(net384),
    .D(_0559_),
    .RESET_B(_0254_),
    .Q(\cordic_inst.cordic_inst.y[29] ));
 sky130_fd_sc_hd__dfrtp_2 _4833_ (.CLK(net384),
    .D(_0560_),
    .RESET_B(_0255_),
    .Q(\cordic_inst.cordic_inst.y[30] ));
 sky130_fd_sc_hd__dfrtp_1 _4834_ (.CLK(net386),
    .D(_0561_),
    .RESET_B(_0256_),
    .Q(\cordic_inst.cordic_inst.y[31] ));
 sky130_fd_sc_hd__dfxtp_2 _4835_ (.CLK(net383),
    .D(_0008_),
    .Q(\cordic_inst.deg_handler_inst.isNegative ));
 sky130_fd_sc_hd__dfxtp_1 _4836_ (.CLK(net379),
    .D(_0053_),
    .Q(\cordic_inst.cordic_inst.angle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4837_ (.CLK(net379),
    .D(_0064_),
    .Q(\cordic_inst.cordic_inst.angle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4838_ (.CLK(net379),
    .D(_0075_),
    .Q(\cordic_inst.cordic_inst.angle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4839_ (.CLK(net367),
    .D(_0078_),
    .Q(\cordic_inst.cordic_inst.angle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4840_ (.CLK(net367),
    .D(_0079_),
    .Q(\cordic_inst.cordic_inst.angle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4841_ (.CLK(net366),
    .D(_0080_),
    .Q(\cordic_inst.cordic_inst.angle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4842_ (.CLK(net366),
    .D(_0081_),
    .Q(\cordic_inst.cordic_inst.angle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4843_ (.CLK(net366),
    .D(_0082_),
    .Q(\cordic_inst.cordic_inst.angle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4844_ (.CLK(net366),
    .D(_0083_),
    .Q(\cordic_inst.cordic_inst.angle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4845_ (.CLK(net366),
    .D(_0084_),
    .Q(\cordic_inst.cordic_inst.angle[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4846_ (.CLK(net359),
    .D(_0054_),
    .Q(\cordic_inst.cordic_inst.angle[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4847_ (.CLK(net359),
    .D(_0055_),
    .Q(\cordic_inst.cordic_inst.angle[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4848_ (.CLK(net359),
    .D(_0056_),
    .Q(\cordic_inst.cordic_inst.angle[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4849_ (.CLK(net359),
    .D(_0057_),
    .Q(\cordic_inst.cordic_inst.angle[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4850_ (.CLK(net359),
    .D(_0058_),
    .Q(\cordic_inst.cordic_inst.angle[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4851_ (.CLK(net360),
    .D(_0059_),
    .Q(\cordic_inst.cordic_inst.angle[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4852_ (.CLK(net374),
    .D(_0060_),
    .Q(\cordic_inst.cordic_inst.angle[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4853_ (.CLK(net374),
    .D(_0061_),
    .Q(\cordic_inst.cordic_inst.angle[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4854_ (.CLK(net374),
    .D(_0062_),
    .Q(\cordic_inst.cordic_inst.angle[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4855_ (.CLK(net374),
    .D(_0063_),
    .Q(\cordic_inst.cordic_inst.angle[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4856_ (.CLK(net378),
    .D(_0065_),
    .Q(\cordic_inst.cordic_inst.angle[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4857_ (.CLK(net378),
    .D(_0066_),
    .Q(\cordic_inst.cordic_inst.angle[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4858_ (.CLK(net372),
    .D(_0067_),
    .Q(\cordic_inst.cordic_inst.angle[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4859_ (.CLK(net372),
    .D(_0068_),
    .Q(\cordic_inst.cordic_inst.angle[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4860_ (.CLK(net372),
    .D(_0069_),
    .Q(\cordic_inst.cordic_inst.angle[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4861_ (.CLK(net374),
    .D(_0070_),
    .Q(\cordic_inst.cordic_inst.angle[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4862_ (.CLK(net375),
    .D(_0071_),
    .Q(\cordic_inst.cordic_inst.angle[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4863_ (.CLK(net375),
    .D(_0072_),
    .Q(\cordic_inst.cordic_inst.angle[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4864_ (.CLK(net376),
    .D(_0073_),
    .Q(\cordic_inst.cordic_inst.angle[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4865_ (.CLK(net389),
    .D(_0074_),
    .Q(\cordic_inst.cordic_inst.angle[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4866_ (.CLK(net376),
    .D(_0076_),
    .Q(\cordic_inst.cordic_inst.angle[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4867_ (.CLK(net376),
    .D(_0077_),
    .Q(\cordic_inst.cordic_inst.angle[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4868_ (.CLK(net368),
    .D(\axi_controller.reg_input_data[0] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4869_ (.CLK(net368),
    .D(\axi_controller.reg_input_data[1] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4870_ (.CLK(net368),
    .D(\axi_controller.reg_input_data[2] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4871_ (.CLK(net368),
    .D(\axi_controller.reg_input_data[3] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4872_ (.CLK(net365),
    .D(\axi_controller.reg_input_data[4] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4873_ (.CLK(net365),
    .D(\axi_controller.reg_input_data[5] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4874_ (.CLK(net365),
    .D(\axi_controller.reg_input_data[6] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4875_ (.CLK(net365),
    .D(\axi_controller.reg_input_data[7] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4876_ (.CLK(net356),
    .D(\axi_controller.reg_input_data[8] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4877_ (.CLK(net356),
    .D(\axi_controller.reg_input_data[9] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4878_ (.CLK(net356),
    .D(\axi_controller.reg_input_data[10] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4879_ (.CLK(net356),
    .D(\axi_controller.reg_input_data[11] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4880_ (.CLK(net356),
    .D(\axi_controller.reg_input_data[12] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4881_ (.CLK(net356),
    .D(\axi_controller.reg_input_data[13] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4882_ (.CLK(net356),
    .D(\axi_controller.reg_input_data[14] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4883_ (.CLK(net357),
    .D(\axi_controller.reg_input_data[15] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4884_ (.CLK(net357),
    .D(\axi_controller.reg_input_data[16] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4885_ (.CLK(net357),
    .D(\axi_controller.reg_input_data[17] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4886_ (.CLK(net357),
    .D(\axi_controller.reg_input_data[18] ),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4887_ (.CLK(net358),
    .D(_0040_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4888_ (.CLK(net358),
    .D(_0041_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4889_ (.CLK(net358),
    .D(_0042_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4890_ (.CLK(net358),
    .D(_0043_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4891_ (.CLK(net358),
    .D(_0044_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4892_ (.CLK(net373),
    .D(_0045_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4893_ (.CLK(net373),
    .D(_0046_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4894_ (.CLK(net373),
    .D(_0047_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4895_ (.CLK(net373),
    .D(_0048_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4896_ (.CLK(net372),
    .D(_0049_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4897_ (.CLK(net372),
    .D(_0050_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4898_ (.CLK(net373),
    .D(_0051_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4899_ (.CLK(net358),
    .D(_0052_),
    .Q(\cordic_inst.deg_handler_inst.theta_norm[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4900_ (.CLK(net367),
    .D(\cordic_inst.deg_handler_inst.theta_norm[0] ),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4901_ (.CLK(net367),
    .D(_0019_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4902_ (.CLK(net371),
    .D(_0030_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4903_ (.CLK(net371),
    .D(_0033_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4904_ (.CLK(net366),
    .D(_0034_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4905_ (.CLK(net366),
    .D(_0035_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4906_ (.CLK(net367),
    .D(_0036_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4907_ (.CLK(net366),
    .D(_0037_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4908_ (.CLK(net366),
    .D(_0038_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4909_ (.CLK(net360),
    .D(_0039_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4910_ (.CLK(net360),
    .D(_0009_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4911_ (.CLK(net360),
    .D(_0010_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4912_ (.CLK(net359),
    .D(_0011_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4913_ (.CLK(net359),
    .D(_0012_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4914_ (.CLK(net359),
    .D(_0013_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4915_ (.CLK(net359),
    .D(_0014_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4916_ (.CLK(net358),
    .D(_0015_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4917_ (.CLK(net357),
    .D(_0016_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[17] ));
 sky130_fd_sc_hd__dfxtp_2 _4918_ (.CLK(net358),
    .D(_0017_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4919_ (.CLK(net358),
    .D(_0018_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4920_ (.CLK(net373),
    .D(_0020_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4921_ (.CLK(net373),
    .D(_0021_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4922_ (.CLK(net373),
    .D(_0022_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4923_ (.CLK(net373),
    .D(_0023_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4924_ (.CLK(net374),
    .D(_0024_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4925_ (.CLK(net372),
    .D(_0025_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4926_ (.CLK(net372),
    .D(_0026_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4927_ (.CLK(net372),
    .D(_0027_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4928_ (.CLK(net375),
    .D(_0028_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4929_ (.CLK(net375),
    .D(_0029_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4930_ (.CLK(net375),
    .D(_0031_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4931_ (.CLK(net372),
    .D(_0032_),
    .Q(\cordic_inst.deg_handler_inst.theta_abs[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4932_ (.CLK(net368),
    .D(_0562_),
    .Q(\axi_controller.start_pulse_reg ));
 sky130_fd_sc_hd__dfrtp_1 _4933_ (.CLK(net380),
    .D(\axi_controller.done ),
    .RESET_B(_0257_),
    .Q(\cordic_inst.done_d ));
 sky130_fd_sc_hd__dfxtp_1 _4934_ (.CLK(net385),
    .D(_0563_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _4935_ (.CLK(net382),
    .D(_0564_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _4936_ (.CLK(net385),
    .D(_0565_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _4937_ (.CLK(net385),
    .D(_0566_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _4938_ (.CLK(net384),
    .D(_0567_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _4939_ (.CLK(net387),
    .D(_0568_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _4940_ (.CLK(net393),
    .D(_0569_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _4941_ (.CLK(net392),
    .D(_0570_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _4942_ (.CLK(net393),
    .D(_0571_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _4943_ (.CLK(net394),
    .D(_0572_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _4944_ (.CLK(net395),
    .D(_0573_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _4945_ (.CLK(net403),
    .D(_0574_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _4946_ (.CLK(net403),
    .D(_0575_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _4947_ (.CLK(net407),
    .D(_0576_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _4948_ (.CLK(net407),
    .D(_0577_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _4949_ (.CLK(net407),
    .D(_0578_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _4950_ (.CLK(net406),
    .D(_0579_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _4951_ (.CLK(net406),
    .D(_0580_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _4952_ (.CLK(net407),
    .D(_0581_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _4953_ (.CLK(net402),
    .D(_0582_),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _4954_ (.CLK(net402),
    .D(_0583_),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_1 _4955_ (.CLK(net402),
    .D(_0584_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_1 _4956_ (.CLK(net402),
    .D(_0585_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _4957_ (.CLK(net402),
    .D(_0586_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _4958_ (.CLK(net399),
    .D(_0587_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _4959_ (.CLK(net398),
    .D(_0588_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 _4960_ (.CLK(net399),
    .D(_0589_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _4961_ (.CLK(net398),
    .D(_0590_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _4962_ (.CLK(net398),
    .D(_0591_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 _4963_ (.CLK(net398),
    .D(_0592_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _4964_ (.CLK(net399),
    .D(_0593_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _4965_ (.CLK(net380),
    .D(_0594_),
    .Q(net112));
 sky130_fd_sc_hd__conb_1 cordic_system_410 (.LO(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_2028_));
 sky130_fd_sc_hd__clkbuf_1 _4968_ (.A(net108),
    .X(net109));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_828 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(aclk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(araddr[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(araddr[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(araddr[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(araddr[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(araddr[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(araddr[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(araddr[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(araddr[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(araddr[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(araddr[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(araddr[19]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(araddr[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(araddr[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(araddr[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(araddr[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(araddr[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(araddr[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(araddr[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(araddr[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(araddr[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(araddr[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(araddr[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(araddr[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(araddr[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(araddr[31]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(araddr[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(araddr[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(araddr[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(araddr[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(araddr[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(araddr[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(araddr[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(aresetn),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(arvalid),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(awaddr[0]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(awaddr[10]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(awaddr[11]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(awaddr[12]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(awaddr[13]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(awaddr[14]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(awaddr[15]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(awaddr[16]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(awaddr[17]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(awaddr[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(awaddr[19]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(awaddr[1]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(awaddr[20]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(awaddr[21]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(awaddr[22]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(awaddr[23]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(awaddr[24]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(awaddr[25]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(awaddr[26]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(awaddr[27]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(awaddr[28]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(awaddr[29]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(awaddr[2]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(awaddr[30]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(awaddr[31]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(awaddr[3]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(awaddr[4]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(awaddr[5]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(awaddr[6]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(awaddr[7]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(awaddr[8]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(awaddr[9]),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(awvalid),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(bready),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(rready),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(wdata[0]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(wdata[10]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(wdata[11]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(wdata[12]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(wdata[13]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(wdata[14]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(wdata[15]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(wdata[16]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(wdata[17]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(wdata[18]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(wdata[19]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(wdata[1]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(wdata[20]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(wdata[21]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(wdata[22]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(wdata[23]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(wdata[24]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(wdata[25]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(wdata[26]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(wdata[27]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(wdata[28]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(wdata[29]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(wdata[2]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(wdata[30]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(wdata[31]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(wdata[3]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(wdata[4]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(wdata[5]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(wdata[6]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(wdata[7]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(wdata[8]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(wdata[9]),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input103 (.A(wstrb[0]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(wstrb[1]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(wstrb[2]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(wstrb[3]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(wvalid),
    .X(net107));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(arready));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(awready));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(bresp[1]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(bvalid));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(rdata[0]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(rdata[10]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(rdata[11]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(rdata[12]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(rdata[13]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(rdata[14]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(rdata[15]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(rdata[16]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(rdata[17]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(rdata[18]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(rdata[19]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(rdata[1]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(rdata[20]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(rdata[21]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(rdata[22]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(rdata[23]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(rdata[24]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(rdata[25]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(rdata[26]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(rdata[27]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(rdata[28]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(rdata[29]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(rdata[2]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(rdata[30]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(rdata[31]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(rdata[3]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(rdata[4]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(rdata[5]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(rdata[6]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(rdata[7]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(rdata[8]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(rdata[9]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(rresp[1]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(rvalid));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(wready));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net149),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(_1790_),
    .X(net149));
 sky130_fd_sc_hd__buf_2 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net153),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(_1781_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 max_cap154 (.A(_0743_),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(_2256_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(_2256_),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(\cordic_inst.cordic_inst.next_state[1] ),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(_0629_),
    .X(net159));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(_0629_),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__buf_2 fanout162 (.A(net164),
    .X(net162));
 sky130_fd_sc_hd__buf_2 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 fanout164 (.A(_0629_),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net169),
    .X(net165));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(_0629_),
    .X(net169));
 sky130_fd_sc_hd__buf_2 fanout170 (.A(_0630_),
    .X(net170));
 sky130_fd_sc_hd__buf_2 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(_0628_),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(_0628_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 fanout174 (.A(_0628_),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_2 fanout178 (.A(_0627_),
    .X(net178));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(net182),
    .X(net179));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(_0626_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net186),
    .X(net183));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(net186),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(_0626_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(_1929_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 fanout188 (.A(_1929_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_2 fanout190 (.A(_1929_),
    .X(net190));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(_1927_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(_1927_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net199),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(net199),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net199),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 fanout199 (.A(_1926_),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_2 fanout201 (.A(\cordic_inst.sign_handler_inst.done_pulse ),
    .X(net201));
 sky130_fd_sc_hd__buf_2 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_2 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_2 fanout205 (.A(\cordic_inst.sign_handler_inst.done_pulse ),
    .X(net205));
 sky130_fd_sc_hd__buf_1 max_cap206 (.A(_1502_),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(net209),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_2 fanout209 (.A(_1472_),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(net213),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_2 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(_1472_),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 fanout215 (.A(_1068_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 max_cap216 (.A(_0709_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 max_cap217 (.A(_0708_),
    .X(net217));
 sky130_fd_sc_hd__buf_2 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 fanout220 (.A(_0680_),
    .X(net220));
 sky130_fd_sc_hd__buf_2 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__buf_2 fanout222 (.A(_0678_),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 fanout223 (.A(_0613_),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 fanout224 (.A(_0613_),
    .X(net224));
 sky130_fd_sc_hd__buf_2 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(_0613_),
    .X(net227));
 sky130_fd_sc_hd__buf_2 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__buf_2 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_2 fanout231 (.A(_0612_),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(_0609_),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(net236),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_2 fanout237 (.A(_0608_),
    .X(net237));
 sky130_fd_sc_hd__buf_2 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(_0607_),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_4 fanout240 (.A(_0607_),
    .X(net240));
 sky130_fd_sc_hd__buf_2 fanout241 (.A(_0607_),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 fanout242 (.A(_0606_),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net247),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net246),
    .X(net244));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(_0606_),
    .X(net247));
 sky130_fd_sc_hd__buf_2 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_2 fanout249 (.A(_0604_),
    .X(net249));
 sky130_fd_sc_hd__buf_2 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_2 fanout251 (.A(_0604_),
    .X(net251));
 sky130_fd_sc_hd__buf_2 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__buf_2 fanout253 (.A(net255),
    .X(net253));
 sky130_fd_sc_hd__buf_2 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 fanout255 (.A(\cordic_inst.deg_handler_inst.theta_norm[31] ),
    .X(net255));
 sky130_fd_sc_hd__buf_2 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_2 fanout257 (.A(\cordic_inst.deg_handler_inst.isNegative ),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_2 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 fanout259 (.A(\cordic_inst.deg_handler_inst.isNegative ),
    .X(net259));
 sky130_fd_sc_hd__buf_2 fanout260 (.A(\cordic_inst.deg_handler_inst.isNegative ),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(\cordic_inst.deg_handler_inst.isNegative ),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 fanout262 (.A(\cordic_inst.cordic_inst.y[31] ),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_4 fanout263 (.A(\cordic_inst.cordic_inst.y[31] ),
    .X(net263));
 sky130_fd_sc_hd__buf_2 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(\cordic_inst.cordic_inst.x[31] ),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__buf_2 fanout267 (.A(\cordic_inst.cordic_inst.z[31] ),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(\cordic_inst.cordic_inst.z[31] ),
    .X(net268));
 sky130_fd_sc_hd__buf_2 fanout269 (.A(\cordic_inst.cordic_inst.z[31] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net273),
    .X(net270));
 sky130_fd_sc_hd__buf_2 fanout271 (.A(net273),
    .X(net271));
 sky130_fd_sc_hd__buf_2 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(\cordic_inst.cordic_inst.z[31] ),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net279),
    .X(net274));
 sky130_fd_sc_hd__buf_2 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 fanout276 (.A(net279),
    .X(net276));
 sky130_fd_sc_hd__buf_2 fanout277 (.A(net279),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_2 fanout279 (.A(\cordic_inst.cordic_inst.i[4] ),
    .X(net279));
 sky130_fd_sc_hd__buf_2 fanout280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__buf_1 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_2 fanout282 (.A(net287),
    .X(net282));
 sky130_fd_sc_hd__buf_2 fanout283 (.A(net287),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 fanout284 (.A(net287),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 fanout285 (.A(net287),
    .X(net285));
 sky130_fd_sc_hd__buf_2 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 fanout287 (.A(\cordic_inst.cordic_inst.i[3] ),
    .X(net287));
 sky130_fd_sc_hd__buf_2 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout289 (.A(net293),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_4 fanout290 (.A(net292),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net293),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_2 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(\cordic_inst.cordic_inst.i[2] ),
    .X(net293));
 sky130_fd_sc_hd__buf_2 fanout294 (.A(net296),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_2 fanout296 (.A(\cordic_inst.cordic_inst.i[1] ),
    .X(net296));
 sky130_fd_sc_hd__buf_2 fanout297 (.A(net300),
    .X(net297));
 sky130_fd_sc_hd__buf_1 fanout298 (.A(net300),
    .X(net298));
 sky130_fd_sc_hd__buf_2 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__buf_2 fanout300 (.A(\cordic_inst.cordic_inst.i[1] ),
    .X(net300));
 sky130_fd_sc_hd__buf_2 fanout301 (.A(\cordic_inst.cordic_inst.i[1] ),
    .X(net301));
 sky130_fd_sc_hd__buf_2 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_2 fanout303 (.A(\cordic_inst.cordic_inst.i[0] ),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__buf_2 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout306 (.A(\cordic_inst.cordic_inst.i[0] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 fanout307 (.A(net312),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(net311),
    .X(net308));
 sky130_fd_sc_hd__buf_2 fanout309 (.A(net312),
    .X(net309));
 sky130_fd_sc_hd__buf_4 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_4 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_2 fanout312 (.A(\cordic_inst.cordic_inst.i[0] ),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 fanout313 (.A(\axi_controller.mode ),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(\axi_controller.mode ),
    .X(net314));
 sky130_fd_sc_hd__buf_2 fanout315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_4 fanout316 (.A(\axi_controller.mode ),
    .X(net316));
 sky130_fd_sc_hd__buf_4 fanout317 (.A(net319),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__buf_2 fanout319 (.A(\axi_controller.rst ),
    .X(net319));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(\axi_controller.rst ),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(net328),
    .X(net321));
 sky130_fd_sc_hd__buf_4 fanout322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(net328),
    .X(net323));
 sky130_fd_sc_hd__buf_4 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 fanout325 (.A(net328),
    .X(net325));
 sky130_fd_sc_hd__buf_4 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__buf_2 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_4 fanout328 (.A(\axi_controller.rst ),
    .X(net328));
 sky130_fd_sc_hd__buf_4 fanout329 (.A(net345),
    .X(net329));
 sky130_fd_sc_hd__buf_2 fanout330 (.A(net345),
    .X(net330));
 sky130_fd_sc_hd__buf_4 fanout331 (.A(net333),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(net345),
    .X(net333));
 sky130_fd_sc_hd__buf_4 fanout334 (.A(net335),
    .X(net334));
 sky130_fd_sc_hd__buf_2 fanout335 (.A(net339),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_4 fanout336 (.A(net339),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_4 fanout338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 fanout339 (.A(net344),
    .X(net339));
 sky130_fd_sc_hd__buf_4 fanout340 (.A(net344),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_2 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__buf_2 fanout345 (.A(\axi_controller.rst ),
    .X(net345));
 sky130_fd_sc_hd__buf_2 fanout346 (.A(net348),
    .X(net346));
 sky130_fd_sc_hd__buf_2 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_2 fanout348 (.A(net34),
    .X(net348));
 sky130_fd_sc_hd__buf_2 fanout349 (.A(net34),
    .X(net349));
 sky130_fd_sc_hd__buf_2 fanout350 (.A(net34),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 fanout351 (.A(net354),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 fanout352 (.A(net354),
    .X(net352));
 sky130_fd_sc_hd__buf_1 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 fanout354 (.A(net361),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 fanout355 (.A(net361),
    .X(net355));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout356 (.A(net361),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 fanout357 (.A(net361),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 fanout358 (.A(net361),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_2 fanout361 (.A(net388),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 fanout362 (.A(net365),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_2 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 fanout365 (.A(net388),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__buf_2 fanout367 (.A(net371),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_2 fanout368 (.A(net370),
    .X(net368));
 sky130_fd_sc_hd__buf_1 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_2 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 fanout371 (.A(net388),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 fanout372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_2 fanout374 (.A(net378),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 fanout375 (.A(net377),
    .X(net375));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_2 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 fanout378 (.A(net388),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(net383),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 fanout380 (.A(net382),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_2 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 fanout382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_2 fanout383 (.A(net387),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 fanout384 (.A(net387),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_2 fanout385 (.A(net387),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_2 fanout388 (.A(net1),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__buf_2 fanout391 (.A(net408),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_2 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(net408),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_2 fanout394 (.A(net408),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 fanout395 (.A(net408),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout397 (.A(net408),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 fanout399 (.A(net402),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__buf_2 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 fanout402 (.A(net408),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 fanout404 (.A(net408),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_2 fanout406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_4 fanout408 (.A(net1),
    .X(net408));
 sky130_fd_sc_hd__conb_1 cordic_system_409 (.LO(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net361));
 sky130_fd_sc_hd__fill_2 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_841 ();
 assign bresp[0] = net409;
 assign rresp[0] = net410;
endmodule
