// `include "picorv32.v"
// `include "axi4_master_riscv.v"
// `include "axi4_interconnect.v"
// `include "dram_controller.v"
// `include "cordic_system.v"

module top (
    input wire clk,
    input wire reset_n,
    
    // DRAM Interface (simplified)
    output wire                    dram_ck,
    output wire                    dram_cs,
    output wire                    dram_we,
    output wire                    dram_ras,
    output wire                    dram_cas,
    output wire [13:0]             dram_addr,
    output wire [2:0]              dram_ba,
    inout  wire [31:0]             dram_dq,
    output wire [3:0]              dram_dm,
    output wire                    dram_dqs,
    
    // External debug/control signals
    output wire trap
);

    // System Parameters
    parameter ADDR_WIDTH = 32;
    parameter DATA_WIDTH = 32;
    parameter AXI4_ID_WIDTH = 4;
    parameter LPDDR4_CAPACITY_GB = 4;

    // Clock and reset for all components
    wire clk_sys = clk;
    wire reset_sys_n = reset_n;
    
    // ========== PicoRV32 to AXI4 Master Connection ==========
    // PicoRV32 Memory Interface
    wire        mem_valid;
    wire        mem_instr;
    wire        mem_ready;
    wire [31:0] mem_addr;
    wire [31:0] mem_wdata;
    wire [3:0]  mem_wstrb;
    wire [31:0] mem_rdata;
    
    // ========== AXI4 Master Interface Signals (from PicoRV32) ==========
    // Write Address Channel
    wire [AXI4_ID_WIDTH-1:0]   cpu_m_axi_awid;
    wire [ADDR_WIDTH-1:0]      cpu_m_axi_awaddr;
    wire [7:0]                 cpu_m_axi_awlen;
    wire [2:0]                 cpu_m_axi_awsize;
    wire [1:0]                 cpu_m_axi_awburst;
    wire                       cpu_m_axi_awvalid;
    wire                       cpu_m_axi_awready;
    
    // Write Data Channel
    wire [DATA_WIDTH-1:0]      cpu_m_axi_wdata;
    wire [(DATA_WIDTH/8)-1:0]  cpu_m_axi_wstrb;
    wire                       cpu_m_axi_wlast;
    wire                       cpu_m_axi_wvalid;
    wire                       cpu_m_axi_wready;
    
    // Write Response Channel
    wire [AXI4_ID_WIDTH-1:0]   cpu_m_axi_bid;
    wire [1:0]                 cpu_m_axi_bresp;
    wire                       cpu_m_axi_bvalid;
    wire                       cpu_m_axi_bready;
    
    // Read Address Channel
    wire [AXI4_ID_WIDTH-1:0]   cpu_m_axi_arid;
    wire [ADDR_WIDTH-1:0]      cpu_m_axi_araddr;
    wire [7:0]                 cpu_m_axi_arlen;
    wire [2:0]                 cpu_m_axi_arsize;
    wire [1:0]                 cpu_m_axi_arburst;
    wire                       cpu_m_axi_arvalid;
    wire                       cpu_m_axi_arready;
    
    // Read Data Channel
    wire [AXI4_ID_WIDTH-1:0]   cpu_m_axi_rid;
    wire [DATA_WIDTH-1:0]      cpu_m_axi_rdata;
    wire [1:0]                 cpu_m_axi_rresp;
    wire                       cpu_m_axi_rlast;
    wire                       cpu_m_axi_rvalid;
    wire                       cpu_m_axi_rready;
    
    // ========== AXI4 Master Interface for SA (Placeholder) ==========
    // Write Address Channel
    wire [AXI4_ID_WIDTH-1:0]   sa_m_axi_awid;
    wire [ADDR_WIDTH-1:0]      sa_m_axi_awaddr;
    wire [7:0]                 sa_m_axi_awlen;
    wire [2:0]                 sa_m_axi_awsize;
    wire [1:0]                 sa_m_axi_awburst;
    wire                       sa_m_axi_awvalid;
    wire                       sa_m_axi_awready;
    
    // Write Data Channel
    wire [DATA_WIDTH-1:0]      sa_m_axi_wdata;
    wire [(DATA_WIDTH/8)-1:0]  sa_m_axi_wstrb;
    wire                       sa_m_axi_wlast;
    wire                       sa_m_axi_wvalid;
    wire                       sa_m_axi_wready;
    
    // Write Response Channel
    wire [AXI4_ID_WIDTH-1:0]   sa_m_axi_bid;
    wire [1:0]                 sa_m_axi_bresp;
    wire                       sa_m_axi_bvalid;
    wire                       sa_m_axi_bready;
    
    // Read Address Channel
    wire [AXI4_ID_WIDTH-1:0]   sa_m_axi_arid;
    wire [ADDR_WIDTH-1:0]      sa_m_axi_araddr;
    wire [7:0]                 sa_m_axi_arlen;
    wire [2:0]                 sa_m_axi_arsize;
    wire [1:0]                 sa_m_axi_arburst;
    wire                       sa_m_axi_arvalid;
    wire                       sa_m_axi_arready;
    
    // Read Data Channel
    wire [AXI4_ID_WIDTH-1:0]   sa_m_axi_rid;
    wire [DATA_WIDTH-1:0]      sa_m_axi_rdata;
    wire [1:0]                 sa_m_axi_rresp;
    wire                       sa_m_axi_rlast;
    wire                       sa_m_axi_rvalid;
    wire                       sa_m_axi_rready;

    // ========== AXI4-Lite Interface for Cordic (Placeholder) ==========
    wire [ADDR_WIDTH-1:0]      cordic_axil_awaddr;
    wire [2:0]                 cordic_axil_awprot;
    wire                       cordic_axil_awvalid;
    wire                       cordic_axil_awready;
    wire [DATA_WIDTH-1:0]      cordic_axil_wdata;
    wire [(DATA_WIDTH/8)-1:0]  cordic_axil_wstrb;
    wire                       cordic_axil_wvalid;
    wire                       cordic_axil_wready;
    wire [1:0]                 cordic_axil_bresp;
    wire                       cordic_axil_bvalid;
    wire                       cordic_axil_bready;
    wire [ADDR_WIDTH-1:0]      cordic_axil_araddr;
    wire [2:0]                 cordic_axil_arprot;
    wire                       cordic_axil_arvalid;
    wire                       cordic_axil_arready;
    wire [DATA_WIDTH-1:0]      cordic_axil_rdata;
    wire [1:0]                 cordic_axil_rresp;
    wire                       cordic_axil_rvalid;
    wire                       cordic_axil_rready;

    // ========== AXI4-Lite Interface for SA Control (Placeholder) ==========
    wire [ADDR_WIDTH-1:0]      sa_axil_awaddr;
    wire [2:0]                 sa_axil_awprot;
    wire                       sa_axil_awvalid;
    wire                       sa_axil_awready;
    wire [DATA_WIDTH-1:0]      sa_axil_wdata;
    wire [(DATA_WIDTH/8)-1:0]  sa_axil_wstrb;
    wire                       sa_axil_wvalid;
    wire                       sa_axil_wready;
    wire [1:0]                 sa_axil_bresp;
    wire                       sa_axil_bvalid;
    wire                       sa_axil_bready;
    wire [ADDR_WIDTH-1:0]      sa_axil_araddr;
    wire [2:0]                 sa_axil_arprot;
    wire                       sa_axil_arvalid;
    wire                       sa_axil_arready;
    wire [DATA_WIDTH-1:0]      sa_axil_rdata;
    wire [1:0]                 sa_axil_rresp;
    wire                       sa_axil_rvalid;
    wire                       sa_axil_rready;
    
    // ========== DRAM Controller AXI4 Interface ==========
    // Write Address Channel
    wire [AXI4_ID_WIDTH-1:0]   dram_s_axi_awid;
    wire [ADDR_WIDTH-1:0]      dram_s_axi_awaddr;
    wire [7:0]                 dram_s_axi_awlen;
    wire [2:0]                 dram_s_axi_awsize;
    wire [1:0]                 dram_s_axi_awburst;
    wire                       dram_s_axi_awvalid;
    wire                       dram_s_axi_awready;
    
    // Write Data Channel
    wire [DATA_WIDTH-1:0]      dram_s_axi_wdata;
    wire [(DATA_WIDTH/8)-1:0]  dram_s_axi_wstrb;
    wire                       dram_s_axi_wlast;
    wire                       dram_s_axi_wvalid;
    wire                       dram_s_axi_wready;
    
    // Write Response Channel
    wire [AXI4_ID_WIDTH-1:0]   dram_s_axi_bid;
    wire [1:0]                 dram_s_axi_bresp;
    wire                       dram_s_axi_bvalid;
    wire                       dram_s_axi_bready;
    
    // Read Address Channel
    wire [AXI4_ID_WIDTH-1:0]   dram_s_axi_arid;
    wire [ADDR_WIDTH-1:0]      dram_s_axi_araddr;
    wire [7:0]                 dram_s_axi_arlen;
    wire [2:0]                 dram_s_axi_arsize;
    wire [1:0]                 dram_s_axi_arburst;
    wire                       dram_s_axi_arvalid;
    wire                       dram_s_axi_arready;
    
    // Read Data Channel
    wire [AXI4_ID_WIDTH-1:0]   dram_s_axi_rid;
    wire [DATA_WIDTH-1:0]      dram_s_axi_rdata;
    wire [1:0]                 dram_s_axi_rresp;
    wire                       dram_s_axi_rlast;
    wire                       dram_s_axi_rvalid;
    wire                       dram_s_axi_rready;
    
    // ========== Additional wires for unused PicoRV32 ports ==========
    wire        mem_la_read;
    wire        mem_la_write;
    wire [31:0] mem_la_addr;
    wire [31:0] mem_la_wdata;
    wire [3:0]  mem_la_wstrb;
    
    wire        pcpi_valid;
    wire [31:0] pcpi_insn;
    wire [31:0] pcpi_rs1;
    wire [31:0] pcpi_rs2;
    
    wire [31:0] eoi;
    
    wire        trace_valid;
    wire [35:0] trace_data;
    
    // ========== Instantiate PicoRV32 CPU ==========
    picorv32 cpu (
        .clk(clk_sys),
        .resetn(reset_sys_n),
        .trap(trap),
        
        // Memory interface
        .mem_valid(mem_valid),
        .mem_instr(mem_instr),
        .mem_ready(mem_ready),
        .mem_addr(mem_addr),
        .mem_wdata(mem_wdata),
        .mem_wstrb(mem_wstrb),
        .mem_rdata(mem_rdata),
        
        // Look-ahead interface (unused)
        .mem_la_read(mem_la_read),
        .mem_la_write(mem_la_write),
        .mem_la_addr(mem_la_addr),
        .mem_la_wdata(mem_la_wdata),
        .mem_la_wstrb(mem_la_wstrb),
        
        // PCPI interface (unused since ENABLE_PCPI=0)
        .pcpi_valid(pcpi_valid),
        .pcpi_insn(pcpi_insn),
        .pcpi_rs1(pcpi_rs1),
        .pcpi_rs2(pcpi_rs2),
        .pcpi_wr(1'b0),
        .pcpi_rd(32'h0),
        .pcpi_wait(1'b0),
        .pcpi_ready(1'b0),
        
        // IRQ interface (unused since ENABLE_IRQ=0)
        .irq(32'h0),
        .eoi(eoi),
        
        // Trace interface (unused since ENABLE_TRACE=0)
        .trace_valid(trace_valid),
        .trace_data(trace_data)
    );
    
    // ========== Instantiate AXI4 Master Bridge for CPU ==========
    axi4_master cpu_axi_master (
        .aclk(clk_sys),
        .aresetn(reset_sys_n),
        
        // PicoRV32 memory interface
        .mem_valid(mem_valid),
        .mem_instr(mem_instr),
        .mem_ready(mem_ready),
        .mem_addr(mem_addr),
        .mem_wdata(mem_wdata),
        .mem_wstrb(mem_wstrb),
        .mem_rdata(mem_rdata),
        
        // AXI4 master interface
        .m_axi_awid(cpu_m_axi_awid),
        .m_axi_awaddr(cpu_m_axi_awaddr),
        .m_axi_awlen(cpu_m_axi_awlen),
        .m_axi_awsize(cpu_m_axi_awsize),
        .m_axi_awburst(cpu_m_axi_awburst),
        .m_axi_awvalid(cpu_m_axi_awvalid),
        .m_axi_awready(cpu_m_axi_awready),
        
        .m_axi_wdata(cpu_m_axi_wdata),
        .m_axi_wstrb(cpu_m_axi_wstrb),
        .m_axi_wlast(cpu_m_axi_wlast),
        .m_axi_wvalid(cpu_m_axi_wvalid),
        .m_axi_wready(cpu_m_axi_wready),
        
        .m_axi_bid(cpu_m_axi_bid),
        .m_axi_bresp(cpu_m_axi_bresp),
        .m_axi_bvalid(cpu_m_axi_bvalid),
        .m_axi_bready(cpu_m_axi_bready),
        
        .m_axi_arid(cpu_m_axi_arid),
        .m_axi_araddr(cpu_m_axi_araddr),
        .m_axi_arlen(cpu_m_axi_arlen),
        .m_axi_arsize(cpu_m_axi_arsize),
        .m_axi_arburst(cpu_m_axi_arburst),
        .m_axi_arvalid(cpu_m_axi_arvalid),
        .m_axi_arready(cpu_m_axi_arready),
        
        .m_axi_rid(cpu_m_axi_rid),
        .m_axi_rdata(cpu_m_axi_rdata),
        .m_axi_rresp(cpu_m_axi_rresp),
        .m_axi_rlast(cpu_m_axi_rlast),
        .m_axi_rvalid(cpu_m_axi_rvalid),
        .m_axi_rready(cpu_m_axi_rready)
    );

    // ========== Instantiate AXI4 Interconnect ==========
    axi_interconnect #(
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(DATA_WIDTH),
        .AXI4_ID_WIDTH(AXI4_ID_WIDTH)
    ) axi_interconnect_inst (
        // Common signals
        .ACLK(clk_sys),
        .ARESETN(reset_sys_n),
        
        // Slave Port 0: AXI4 from RISC-V (S0_AXI4_...)
        .S0_AXI4_AWID(cpu_m_axi_awid),
        .S0_AXI4_AWADDR(cpu_m_axi_awaddr),
        .S0_AXI4_AWLEN(cpu_m_axi_awlen),
        .S0_AXI4_AWSIZE(cpu_m_axi_awsize),
        .S0_AXI4_AWBURST(cpu_m_axi_awburst),
        .S0_AXI4_AWVALID(cpu_m_axi_awvalid),
        .S0_AXI4_AWREADY(cpu_m_axi_awready),
        
        .S0_AXI4_WDATA(cpu_m_axi_wdata),
        .S0_AXI4_WSTRB(cpu_m_axi_wstrb),
        .S0_AXI4_WLAST(cpu_m_axi_wlast),
        .S0_AXI4_WVALID(cpu_m_axi_wvalid),
        .S0_AXI4_WREADY(cpu_m_axi_wready),
        
        .S0_AXI4_BID(cpu_m_axi_bid),
        .S0_AXI4_BRESP(cpu_m_axi_bresp),
        .S0_AXI4_BVALID(cpu_m_axi_bvalid),
        .S0_AXI4_BREADY(cpu_m_axi_bready),
        
        .S0_AXI4_ARID(cpu_m_axi_arid),
        .S0_AXI4_ARADDR(cpu_m_axi_araddr),
        .S0_AXI4_ARLEN(cpu_m_axi_arlen),
        .S0_AXI4_ARSIZE(cpu_m_axi_arsize),
        .S0_AXI4_ARBURST(cpu_m_axi_arburst),
        .S0_AXI4_ARVALID(cpu_m_axi_arvalid),
        .S0_AXI4_ARREADY(cpu_m_axi_arready),
        
        .S0_AXI4_RID(cpu_m_axi_rid),
        .S0_AXI4_RDATA(cpu_m_axi_rdata),
        .S0_AXI4_RRESP(cpu_m_axi_rresp),
        .S0_AXI4_RLAST(cpu_m_axi_rlast),
        .S0_AXI4_RVALID(cpu_m_axi_rvalid),
        .S0_AXI4_RREADY(cpu_m_axi_rready),
        
        // Slave Port 1: AXI4 from SA (S1_AXI4_...)
        .S1_AXI4_AWID(sa_m_axi_awid),
        .S1_AXI4_AWADDR(sa_m_axi_awaddr),
        .S1_AXI4_AWLEN(sa_m_axi_awlen),
        .S1_AXI4_AWSIZE(sa_m_axi_awsize),
        .S1_AXI4_AWBURST(sa_m_axi_awburst),
        .S1_AXI4_AWVALID(sa_m_axi_awvalid),
        .S1_AXI4_AWREADY(sa_m_axi_awready),
        
        .S1_AXI4_WDATA(sa_m_axi_wdata),
        .S1_AXI4_WSTRB(sa_m_axi_wstrb),
        .S1_AXI4_WLAST(sa_m_axi_wlast),
        .S1_AXI4_WVALID(sa_m_axi_wvalid),
        .S1_AXI4_WREADY(sa_m_axi_wready),
        
        .S1_AXI4_BID(sa_m_axi_bid),
        .S1_AXI4_BRESP(sa_m_axi_bresp),
        .S1_AXI4_BVALID(sa_m_axi_bvalid),
        .S1_AXI4_BREADY(sa_m_axi_bready),
        
        .S1_AXI4_ARID(sa_m_axi_arid),
        .S1_AXI4_ARADDR(sa_m_axi_araddr),
        .S1_AXI4_ARLEN(sa_m_axi_arlen),
        .S1_AXI4_ARSIZE(sa_m_axi_arsize),
        .S1_AXI4_ARBURST(sa_m_axi_arburst),
        .S1_AXI4_ARVALID(sa_m_axi_arvalid),
        .S1_AXI4_ARREADY(sa_m_axi_arready),
        
        .S1_AXI4_RID(sa_m_axi_rid),
        .S1_AXI4_RDATA(sa_m_axi_rdata),
        .S1_AXI4_RRESP(sa_m_axi_rresp),
        .S1_AXI4_RLAST(sa_m_axi_rlast),
        .S1_AXI4_RVALID(sa_m_axi_rvalid),
        .S1_AXI4_RREADY(sa_m_axi_rready),
        
        // Master Port 0: AXI4-Lite to CORDIC (M0_AXI4LITE_...)
        .M0_AXI4LITE_AWADDR(cordic_axil_awaddr),
        .M0_AXI4LITE_AWPROT(cordic_axil_awprot),
        .M0_AXI4LITE_AWVALID(cordic_axil_awvalid),
        .M0_AXI4LITE_AWREADY(cordic_axil_awready),
        
        .M0_AXI4LITE_WDATA(cordic_axil_wdata),
        .M0_AXI4LITE_WSTRB(cordic_axil_wstrb),
        .M0_AXI4LITE_WVALID(cordic_axil_wvalid),
        .M0_AXI4LITE_WREADY(cordic_axil_wready),
        
        .M0_AXI4LITE_BRESP(cordic_axil_bresp),
        .M0_AXI4LITE_BVALID(cordic_axil_bvalid),
        .M0_AXI4LITE_BREADY(cordic_axil_bready),
        
        .M0_AXI4LITE_ARADDR(cordic_axil_araddr),
        .M0_AXI4LITE_ARPROT(cordic_axil_arprot),
        .M0_AXI4LITE_ARVALID(cordic_axil_arvalid),
        .M0_AXI4LITE_ARREADY(cordic_axil_arready),
        
        .M0_AXI4LITE_RDATA(cordic_axil_rdata),
        .M0_AXI4LITE_RRESP(cordic_axil_rresp),
        .M0_AXI4LITE_RVALID(cordic_axil_rvalid),
        .M0_AXI4LITE_RREADY(cordic_axil_rready),
        
        // Master Port 1: AXI4-Lite to SA (M1_AXI4LITE_...)
        .M1_AXI4LITE_AWADDR(sa_axil_awaddr),
        .M1_AXI4LITE_AWPROT(sa_axil_awprot),
        .M1_AXI4LITE_AWVALID(sa_axil_awvalid),
        .M1_AXI4LITE_AWREADY(sa_axil_awready),
        
        .M1_AXI4LITE_WDATA(sa_axil_wdata),
        .M1_AXI4LITE_WSTRB(sa_axil_wstrb),
        .M1_AXI4LITE_WVALID(sa_axil_wvalid),
        .M1_AXI4LITE_WREADY(sa_axil_wready),
        
        .M1_AXI4LITE_BRESP(sa_axil_bresp),
        .M1_AXI4LITE_BVALID(sa_axil_bvalid),
        .M1_AXI4LITE_BREADY(sa_axil_bready),
        
        .M1_AXI4LITE_ARADDR(sa_axil_araddr),
        .M1_AXI4LITE_ARPROT(sa_axil_arprot),
        .M1_AXI4LITE_ARVALID(sa_axil_arvalid),
        .M1_AXI4LITE_ARREADY(sa_axil_arready),
        
        .M1_AXI4LITE_RDATA(sa_axil_rdata),
        .M1_AXI4LITE_RRESP(sa_axil_rresp),
        .M1_AXI4LITE_RVALID(sa_axil_rvalid),
        .M1_AXI4LITE_RREADY(sa_axil_rready),
        
        // Master Port 2: AXI4 to DRAM Controller (M2_AXI4_...)
        .M2_AXI4_AWID(dram_s_axi_awid),
        .M2_AXI4_AWADDR(dram_s_axi_awaddr),
        .M2_AXI4_AWLEN(dram_s_axi_awlen),
        .M2_AXI4_AWSIZE(dram_s_axi_awsize),
        .M2_AXI4_AWBURST(dram_s_axi_awburst),
        .M2_AXI4_AWVALID(dram_s_axi_awvalid),
        .M2_AXI4_AWREADY(dram_s_axi_awready),
        
        .M2_AXI4_WDATA(dram_s_axi_wdata),
        .M2_AXI4_WSTRB(dram_s_axi_wstrb),
        .M2_AXI4_WLAST(dram_s_axi_wlast),
        .M2_AXI4_WVALID(dram_s_axi_wvalid),
        .M2_AXI4_WREADY(dram_s_axi_wready),
        
        .M2_AXI4_BID(dram_s_axi_bid),
        .M2_AXI4_BRESP(dram_s_axi_bresp),
        .M2_AXI4_BVALID(dram_s_axi_bvalid),
        .M2_AXI4_BREADY(dram_s_axi_bready),
        
        .M2_AXI4_ARID(dram_s_axi_arid),
        .M2_AXI4_ARADDR(dram_s_axi_araddr),
        .M2_AXI4_ARLEN(dram_s_axi_arlen),
        .M2_AXI4_ARSIZE(dram_s_axi_arsize),
        .M2_AXI4_ARBURST(dram_s_axi_arburst),
        .M2_AXI4_ARVALID(dram_s_axi_arvalid),
        .M2_AXI4_ARREADY(dram_s_axi_arready),
        
        .M2_AXI4_RID(dram_s_axi_rid),
        .M2_AXI4_RDATA(dram_s_axi_rdata),
        .M2_AXI4_RRESP(dram_s_axi_rresp),
        .M2_AXI4_RLAST(dram_s_axi_rlast),
        .M2_AXI4_RVALID(dram_s_axi_rvalid),
        .M2_AXI4_RREADY(dram_s_axi_rready)
    );
    
    // ========== Instantiate DRAM Controller ==========
    dram_controller #(
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(DATA_WIDTH),
        .AXI4_ID_WIDTH(AXI4_ID_WIDTH)
    ) dram_controller_inst (
        // Clock and Reset
        .clk(clk_sys),
        .rst_n(reset_sys_n),
        
        // AXI4 Slave Interface
        .M2_AXI4_AWID(dram_s_axi_awid),
        .M2_AXI4_AWADDR(dram_s_axi_awaddr),
        .M2_AXI4_AWLEN(dram_s_axi_awlen),
        .M2_AXI4_AWSIZE(dram_s_axi_awsize),
        .M2_AXI4_AWBURST(dram_s_axi_awburst),
        .M2_AXI4_AWVALID(dram_s_axi_awvalid),
        .M2_AXI4_AWREADY(dram_s_axi_awready),
        
        .M2_AXI4_WDATA(dram_s_axi_wdata),
        .M2_AXI4_WSTRB(dram_s_axi_wstrb),
        .M2_AXI4_WLAST(dram_s_axi_wlast),
        .M2_AXI4_WVALID(dram_s_axi_wvalid),
        .M2_AXI4_WREADY(dram_s_axi_wready),
        
        .M2_AXI4_BID(dram_s_axi_bid),
        .M2_AXI4_BRESP(dram_s_axi_bresp),
        .M2_AXI4_BVALID(dram_s_axi_bvalid),
        .M2_AXI4_BREADY(dram_s_axi_bready),
        
        .M2_AXI4_ARID(dram_s_axi_arid),
        .M2_AXI4_ARADDR(dram_s_axi_araddr),
        .M2_AXI4_ARLEN(dram_s_axi_arlen),
        .M2_AXI4_ARSIZE(dram_s_axi_arsize),
        .M2_AXI4_ARBURST(dram_s_axi_arburst),
        .M2_AXI4_ARVALID(dram_s_axi_arvalid),
        .M2_AXI4_ARREADY(dram_s_axi_arready),
        
        .M2_AXI4_RID(dram_s_axi_rid),
        .M2_AXI4_RDATA(dram_s_axi_rdata),
        .M2_AXI4_RRESP(dram_s_axi_rresp),
        .M2_AXI4_RLAST(dram_s_axi_rlast),
        .M2_AXI4_RVALID(dram_s_axi_rvalid),
        .M2_AXI4_RREADY(dram_s_axi_rready),
        
        // DRAM Physical Interface
        .dram_ck(dram_ck),
        .dram_cs(dram_cs),
        .dram_we(dram_we),
        .dram_ras(dram_ras),
        .dram_cas(dram_cas),
        .dram_addr(dram_addr),
        .dram_ba(dram_ba),
        .dram_dq(dram_dq),
        .dram_dm(dram_dm),
        .dram_dqs(dram_dqs)
    );

    // ========== Instantiate CORDIX ==========

    cordic_system cordic_inst (
        .aclk(clk_sys),
        .aresetn(reset_sys_n),
        .awaddr(cordic_axil_awaddr),
        .awvalid(cordic_axil_awvalid),
        .awready(cordic_axil_awready),
        .wdata(cordic_axil_wdata),
        .wstrb(cordic_axil_wstrb),
        .wvalid(cordic_axil_wvalid),
        .wready(cordic_axil_wready),
        .bresp(cordic_axil_bresp),
        .bvalid(cordic_axil_bvalid),
        .bready(cordic_axil_bready),
        .araddr(cordic_axil_araddr),
        .arvalid(cordic_axil_arvalid),
        .arready(cordic_axil_arready),
        .rdata(cordic_axil_rdata),
        .rresp(cordic_axil_rresp),
        .rvalid(cordic_axil_rvalid),
        .rready(cordic_axil_rready)
    );
    
    // ========== Tie off unused SA AXI4 Master signals ==========
    // Write Address Channel
    assign sa_m_axi_awid = {AXI4_ID_WIDTH{1'b0}};
    assign sa_m_axi_awaddr = {ADDR_WIDTH{1'b0}};
    assign sa_m_axi_awlen = 8'h00;
    assign sa_m_axi_awsize = 3'b000;
    assign sa_m_axi_awburst = 2'b00;
    assign sa_m_axi_awvalid = 1'b0;
    
    // Write Data Channel
    assign sa_m_axi_wdata = {DATA_WIDTH{1'b0}};
    assign sa_m_axi_wstrb = {(DATA_WIDTH/8){1'b0}};
    assign sa_m_axi_wlast = 1'b0;
    assign sa_m_axi_wvalid = 1'b0;
    
    // Write Response Channel
    assign sa_m_axi_bready = 1'b0;
    
    // Read Address Channel
    assign sa_m_axi_arid = {AXI4_ID_WIDTH{1'b0}};
    assign sa_m_axi_araddr = {ADDR_WIDTH{1'b0}};
    assign sa_m_axi_arlen = 8'h00;
    assign sa_m_axi_arsize = 3'b000;
    assign sa_m_axi_arburst = 2'b00;
    assign sa_m_axi_arvalid = 1'b0;
    
    // Read Data Channel
    assign sa_m_axi_rready = 1'b0;
    
    // ========== Tie off unused SA AXI4-Lite Control signals ==========
    // Write Address Channel
    assign sa_axil_awready = 1'b0;
    
    // Write Data Channel
    assign sa_axil_wready = 1'b0;
    
    // Write Response Channel
    assign sa_axil_bresp = 2'b00;
    assign sa_axil_bvalid = 1'b0;
    
    // Read Address Channel
    assign sa_axil_arready = 1'b0;
    
    // Read Data Channel
    assign sa_axil_rdata = {DATA_WIDTH{1'b0}};
    assign sa_axil_rresp = 2'b00;
    assign sa_axil_rvalid = 1'b0;
    
    // ========== Tie off unused PicoRV32 outputs ==========
    // Look-ahead interface outputs are not connected anywhere, so they're inherently floating
    // PCPI outputs are not connected since PCPI is disabled
    // IRQ eoi output is not used
    // Trace outputs are not used since tracing is disabled
    
    // Create dummy wires to absorb unused outputs if needed by synthesis tools
    wire dummy_absorb;
    assign dummy_absorb = mem_la_read | mem_la_write | (|mem_la_addr) | (|mem_la_wdata) | (|mem_la_wstrb) |
                         pcpi_valid | (|pcpi_insn) | (|pcpi_rs1) | (|pcpi_rs2) |
                         (|eoi) | trace_valid | (|trace_data);

endmodule
