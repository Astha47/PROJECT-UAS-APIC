VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO picorv32
  CLASS BLOCK ;
  FOREIGN picorv32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 477.045 BY 487.765 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 476.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 476.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 476.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 471.740 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 471.740 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 471.740 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 476.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 476.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 476.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 471.740 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 471.740 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 471.740 334.690 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END clk
  PIN eoi[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END eoi[0]
  PIN eoi[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 486.240 477.045 486.840 ;
    END
  END eoi[10]
  PIN eoi[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END eoi[11]
  PIN eoi[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 483.765 435.070 487.765 ;
    END
  END eoi[12]
  PIN eoi[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END eoi[13]
  PIN eoi[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 483.765 418.970 487.765 ;
    END
  END eoi[14]
  PIN eoi[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 483.765 444.730 487.765 ;
    END
  END eoi[15]
  PIN eoi[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 483.765 380.330 487.765 ;
    END
  END eoi[16]
  PIN eoi[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END eoi[17]
  PIN eoi[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 483.765 396.430 487.765 ;
    END
  END eoi[18]
  PIN eoi[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END eoi[19]
  PIN eoi[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END eoi[1]
  PIN eoi[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 483.765 64.770 487.765 ;
    END
  END eoi[20]
  PIN eoi[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 483.765 402.870 487.765 ;
    END
  END eoi[21]
  PIN eoi[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 483.765 39.010 487.765 ;
    END
  END eoi[22]
  PIN eoi[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END eoi[23]
  PIN eoi[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 442.040 477.045 442.640 ;
    END
  END eoi[24]
  PIN eoi[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 483.765 412.530 487.765 ;
    END
  END eoi[25]
  PIN eoi[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END eoi[26]
  PIN eoi[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 483.765 361.010 487.765 ;
    END
  END eoi[27]
  PIN eoi[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END eoi[28]
  PIN eoi[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END eoi[29]
  PIN eoi[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 483.765 389.990 487.765 ;
    END
  END eoi[2]
  PIN eoi[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 483.765 96.970 487.765 ;
    END
  END eoi[30]
  PIN eoi[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 476.040 477.045 476.640 ;
    END
  END eoi[31]
  PIN eoi[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END eoi[3]
  PIN eoi[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END eoi[4]
  PIN eoi[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 10.240 477.045 10.840 ;
    END
  END eoi[5]
  PIN eoi[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END eoi[6]
  PIN eoi[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END eoi[7]
  PIN eoi[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 483.765 409.310 487.765 ;
    END
  END eoi[8]
  PIN eoi[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 472.640 477.045 473.240 ;
    END
  END eoi[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END irq[15]
  PIN irq[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END irq[16]
  PIN irq[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END irq[17]
  PIN irq[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END irq[18]
  PIN irq[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END irq[19]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END irq[1]
  PIN irq[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END irq[20]
  PIN irq[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END irq[21]
  PIN irq[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END irq[22]
  PIN irq[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END irq[23]
  PIN irq[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END irq[24]
  PIN irq[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END irq[25]
  PIN irq[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END irq[26]
  PIN irq[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END irq[27]
  PIN irq[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END irq[28]
  PIN irq[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END irq[29]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END irq[2]
  PIN irq[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END irq[30]
  PIN irq[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END irq[31]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END irq[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 483.765 357.790 487.765 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 408.040 477.045 408.640 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 483.765 145.270 487.765 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 483.765 109.850 487.765 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 483.765 129.170 487.765 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 347.850 483.765 348.130 487.765 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 305.990 483.765 306.270 487.765 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 483.765 100.190 487.765 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 483.765 84.090 487.765 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 483.765 106.630 487.765 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 483.765 164.590 487.765 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 27.240 477.045 27.840 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 483.765 151.710 487.765 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 483.765 190.350 487.765 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 112.240 477.045 112.840 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 231.240 477.045 231.840 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 132.640 477.045 133.240 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END mem_addr[9]
  PIN mem_instr
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 309.210 483.765 309.490 487.765 ;
    END
  END mem_instr
  PIN mem_la_addr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END mem_la_addr[0]
  PIN mem_la_addr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END mem_la_addr[10]
  PIN mem_la_addr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END mem_la_addr[11]
  PIN mem_la_addr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END mem_la_addr[12]
  PIN mem_la_addr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END mem_la_addr[13]
  PIN mem_la_addr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END mem_la_addr[14]
  PIN mem_la_addr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END mem_la_addr[15]
  PIN mem_la_addr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END mem_la_addr[16]
  PIN mem_la_addr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END mem_la_addr[17]
  PIN mem_la_addr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END mem_la_addr[18]
  PIN mem_la_addr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END mem_la_addr[19]
  PIN mem_la_addr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END mem_la_addr[1]
  PIN mem_la_addr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END mem_la_addr[20]
  PIN mem_la_addr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 483.765 71.210 487.765 ;
    END
  END mem_la_addr[21]
  PIN mem_la_addr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 483.765 77.650 487.765 ;
    END
  END mem_la_addr[22]
  PIN mem_la_addr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 483.765 148.490 487.765 ;
    END
  END mem_la_addr[23]
  PIN mem_la_addr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 312.430 483.765 312.710 487.765 ;
    END
  END mem_la_addr[24]
  PIN mem_la_addr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 315.650 483.765 315.930 487.765 ;
    END
  END mem_la_addr[25]
  PIN mem_la_addr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 483.765 67.990 487.765 ;
    END
  END mem_la_addr[26]
  PIN mem_la_addr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 483.765 154.930 487.765 ;
    END
  END mem_la_addr[27]
  PIN mem_la_addr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 483.765 74.430 487.765 ;
    END
  END mem_la_addr[28]
  PIN mem_la_addr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 483.765 216.110 487.765 ;
    END
  END mem_la_addr[29]
  PIN mem_la_addr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 244.840 477.045 245.440 ;
    END
  END mem_la_addr[2]
  PIN mem_la_addr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 483.765 225.770 487.765 ;
    END
  END mem_la_addr[30]
  PIN mem_la_addr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 483.765 138.830 487.765 ;
    END
  END mem_la_addr[31]
  PIN mem_la_addr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 221.040 477.045 221.640 ;
    END
  END mem_la_addr[3]
  PIN mem_la_addr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 227.840 477.045 228.440 ;
    END
  END mem_la_addr[4]
  PIN mem_la_addr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 210.840 477.045 211.440 ;
    END
  END mem_la_addr[5]
  PIN mem_la_addr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END mem_la_addr[6]
  PIN mem_la_addr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END mem_la_addr[7]
  PIN mem_la_addr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END mem_la_addr[8]
  PIN mem_la_addr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END mem_la_addr[9]
  PIN mem_la_read
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 483.765 303.050 487.765 ;
    END
  END mem_la_read
  PIN mem_la_wdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 108.840 477.045 109.440 ;
    END
  END mem_la_wdata[0]
  PIN mem_la_wdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 323.040 477.045 323.640 ;
    END
  END mem_la_wdata[10]
  PIN mem_la_wdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 34.040 477.045 34.640 ;
    END
  END mem_la_wdata[11]
  PIN mem_la_wdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 44.240 477.045 44.840 ;
    END
  END mem_la_wdata[12]
  PIN mem_la_wdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 302.640 477.045 303.240 ;
    END
  END mem_la_wdata[13]
  PIN mem_la_wdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 78.240 477.045 78.840 ;
    END
  END mem_la_wdata[14]
  PIN mem_la_wdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 299.240 477.045 299.840 ;
    END
  END mem_la_wdata[15]
  PIN mem_la_wdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 265.240 477.045 265.840 ;
    END
  END mem_la_wdata[16]
  PIN mem_la_wdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 85.040 477.045 85.640 ;
    END
  END mem_la_wdata[17]
  PIN mem_la_wdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 88.440 477.045 89.040 ;
    END
  END mem_la_wdata[18]
  PIN mem_la_wdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 278.840 477.045 279.440 ;
    END
  END mem_la_wdata[19]
  PIN mem_la_wdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 251.640 477.045 252.240 ;
    END
  END mem_la_wdata[1]
  PIN mem_la_wdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 261.840 477.045 262.440 ;
    END
  END mem_la_wdata[20]
  PIN mem_la_wdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 255.040 477.045 255.640 ;
    END
  END mem_la_wdata[21]
  PIN mem_la_wdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 115.640 477.045 116.240 ;
    END
  END mem_la_wdata[22]
  PIN mem_la_wdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 387.640 477.045 388.240 ;
    END
  END mem_la_wdata[23]
  PIN mem_la_wdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 357.040 477.045 357.640 ;
    END
  END mem_la_wdata[24]
  PIN mem_la_wdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 380.840 477.045 381.440 ;
    END
  END mem_la_wdata[25]
  PIN mem_la_wdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 397.840 477.045 398.440 ;
    END
  END mem_la_wdata[26]
  PIN mem_la_wdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 343.440 477.045 344.040 ;
    END
  END mem_la_wdata[27]
  PIN mem_la_wdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 360.440 477.045 361.040 ;
    END
  END mem_la_wdata[28]
  PIN mem_la_wdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 479.440 477.045 480.040 ;
    END
  END mem_la_wdata[29]
  PIN mem_la_wdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 122.440 477.045 123.040 ;
    END
  END mem_la_wdata[2]
  PIN mem_la_wdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 377.440 477.045 378.040 ;
    END
  END mem_la_wdata[30]
  PIN mem_la_wdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 316.240 477.045 316.840 ;
    END
  END mem_la_wdata[31]
  PIN mem_la_wdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 125.840 477.045 126.440 ;
    END
  END mem_la_wdata[3]
  PIN mem_la_wdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 57.840 477.045 58.440 ;
    END
  END mem_la_wdata[4]
  PIN mem_la_wdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 119.040 477.045 119.640 ;
    END
  END mem_la_wdata[5]
  PIN mem_la_wdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 207.440 477.045 208.040 ;
    END
  END mem_la_wdata[6]
  PIN mem_la_wdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 170.040 477.045 170.640 ;
    END
  END mem_la_wdata[7]
  PIN mem_la_wdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 64.640 477.045 65.240 ;
    END
  END mem_la_wdata[8]
  PIN mem_la_wdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 71.440 477.045 72.040 ;
    END
  END mem_la_wdata[9]
  PIN mem_la_write
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 296.330 483.765 296.610 487.765 ;
    END
  END mem_la_write
  PIN mem_la_wstrb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 483.765 286.950 487.765 ;
    END
  END mem_la_wstrb[0]
  PIN mem_la_wstrb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 51.040 477.045 51.640 ;
    END
  END mem_la_wstrb[1]
  PIN mem_la_wstrb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 54.440 477.045 55.040 ;
    END
  END mem_la_wstrb[2]
  PIN mem_la_wstrb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 37.440 477.045 38.040 ;
    END
  END mem_la_wstrb[3]
  PIN mem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 270.570 483.765 270.850 487.765 ;
    END
  END mem_rdata[0]
  PIN mem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 167.530 483.765 167.810 487.765 ;
    END
  END mem_rdata[10]
  PIN mem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.410 483.765 180.690 487.765 ;
    END
  END mem_rdata[11]
  PIN mem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 93.470 483.765 93.750 487.765 ;
    END
  END mem_rdata[12]
  PIN mem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 141.770 483.765 142.050 487.765 ;
    END
  END mem_rdata[13]
  PIN mem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 415.470 483.765 415.750 487.765 ;
    END
  END mem_rdata[14]
  PIN mem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.970 483.765 174.250 487.765 ;
    END
  END mem_rdata[15]
  PIN mem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.130 483.765 103.410 487.765 ;
    END
  END mem_rdata[16]
  PIN mem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 119.230 483.765 119.510 487.765 ;
    END
  END mem_rdata[17]
  PIN mem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 177.190 483.765 177.470 487.765 ;
    END
  END mem_rdata[18]
  PIN mem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 132.110 483.765 132.390 487.765 ;
    END
  END mem_rdata[19]
  PIN mem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 351.070 483.765 351.350 487.765 ;
    END
  END mem_rdata[1]
  PIN mem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 431.570 483.765 431.850 487.765 ;
    END
  END mem_rdata[20]
  PIN mem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.030 483.765 87.310 487.765 ;
    END
  END mem_rdata[21]
  PIN mem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.850 483.765 187.130 487.765 ;
    END
  END mem_rdata[22]
  PIN mem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 267.350 483.765 267.630 487.765 ;
    END
  END mem_rdata[23]
  PIN mem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 280.230 483.765 280.510 487.765 ;
    END
  END mem_rdata[24]
  PIN mem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 322.090 483.765 322.370 487.765 ;
    END
  END mem_rdata[25]
  PIN mem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 367.170 483.765 367.450 487.765 ;
    END
  END mem_rdata[26]
  PIN mem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.190 483.765 338.470 487.765 ;
    END
  END mem_rdata[27]
  PIN mem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 273.790 483.765 274.070 487.765 ;
    END
  END mem_rdata[28]
  PIN mem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 341.410 483.765 341.690 487.765 ;
    END
  END mem_rdata[29]
  PIN mem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 421.910 483.765 422.190 487.765 ;
    END
  END mem_rdata[2]
  PIN mem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 363.950 483.765 364.230 487.765 ;
    END
  END mem_rdata[30]
  PIN mem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 328.530 483.765 328.810 487.765 ;
    END
  END mem_rdata[31]
  PIN mem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 260.910 483.765 261.190 487.765 ;
    END
  END mem_rdata[3]
  PIN mem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 370.390 483.765 370.670 487.765 ;
    END
  END mem_rdata[4]
  PIN mem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 264.130 483.765 264.410 487.765 ;
    END
  END mem_rdata[5]
  PIN mem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 373.610 483.765 373.890 487.765 ;
    END
  END mem_rdata[6]
  PIN mem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.870 483.765 158.150 487.765 ;
    END
  END mem_rdata[7]
  PIN mem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.090 483.765 161.370 487.765 ;
    END
  END mem_rdata[8]
  PIN mem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 483.765 135.610 487.765 ;
    END
  END mem_rdata[9]
  PIN mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 318.870 483.765 319.150 487.765 ;
    END
  END mem_ready
  PIN mem_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 283.450 483.765 283.730 487.765 ;
    END
  END mem_valid
  PIN mem_wdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 292.440 477.045 293.040 ;
    END
  END mem_wdata[0]
  PIN mem_wdata[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 326.440 477.045 327.040 ;
    END
  END mem_wdata[10]
  PIN mem_wdata[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 30.640 477.045 31.240 ;
    END
  END mem_wdata[11]
  PIN mem_wdata[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 47.640 477.045 48.240 ;
    END
  END mem_wdata[12]
  PIN mem_wdata[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 306.040 477.045 306.640 ;
    END
  END mem_wdata[13]
  PIN mem_wdata[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 285.640 477.045 286.240 ;
    END
  END mem_wdata[14]
  PIN mem_wdata[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 312.840 477.045 313.440 ;
    END
  END mem_wdata[15]
  PIN mem_wdata[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 272.040 477.045 272.640 ;
    END
  END mem_wdata[16]
  PIN mem_wdata[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 275.440 477.045 276.040 ;
    END
  END mem_wdata[17]
  PIN mem_wdata[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 95.240 477.045 95.840 ;
    END
  END mem_wdata[18]
  PIN mem_wdata[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 282.240 477.045 282.840 ;
    END
  END mem_wdata[19]
  PIN mem_wdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 459.040 477.045 459.640 ;
    END
  END mem_wdata[1]
  PIN mem_wdata[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 268.640 477.045 269.240 ;
    END
  END mem_wdata[20]
  PIN mem_wdata[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 258.440 477.045 259.040 ;
    END
  END mem_wdata[21]
  PIN mem_wdata[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 102.040 477.045 102.640 ;
    END
  END mem_wdata[22]
  PIN mem_wdata[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 336.640 477.045 337.240 ;
    END
  END mem_wdata[23]
  PIN mem_wdata[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 462.440 477.045 463.040 ;
    END
  END mem_wdata[24]
  PIN mem_wdata[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 428.440 477.045 429.040 ;
    END
  END mem_wdata[25]
  PIN mem_wdata[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 421.640 477.045 422.240 ;
    END
  END mem_wdata[26]
  PIN mem_wdata[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 469.240 477.045 469.840 ;
    END
  END mem_wdata[27]
  PIN mem_wdata[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 425.040 477.045 425.640 ;
    END
  END mem_wdata[28]
  PIN mem_wdata[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 445.440 477.045 446.040 ;
    END
  END mem_wdata[29]
  PIN mem_wdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 309.440 477.045 310.040 ;
    END
  END mem_wdata[2]
  PIN mem_wdata[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 329.840 477.045 330.440 ;
    END
  END mem_wdata[30]
  PIN mem_wdata[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 319.640 477.045 320.240 ;
    END
  END mem_wdata[31]
  PIN mem_wdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 350.240 477.045 350.840 ;
    END
  END mem_wdata[3]
  PIN mem_wdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 435.240 477.045 435.840 ;
    END
  END mem_wdata[4]
  PIN mem_wdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 404.640 477.045 405.240 ;
    END
  END mem_wdata[5]
  PIN mem_wdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 353.640 477.045 354.240 ;
    END
  END mem_wdata[6]
  PIN mem_wdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 455.640 477.045 456.240 ;
    END
  END mem_wdata[7]
  PIN mem_wdata[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 68.040 477.045 68.640 ;
    END
  END mem_wdata[8]
  PIN mem_wdata[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 74.840 477.045 75.440 ;
    END
  END mem_wdata[9]
  PIN mem_wstrb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 289.890 483.765 290.170 487.765 ;
    END
  END mem_wstrb[0]
  PIN mem_wstrb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 299.550 483.765 299.830 487.765 ;
    END
  END mem_wstrb[1]
  PIN mem_wstrb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 295.840 477.045 296.440 ;
    END
  END mem_wstrb[2]
  PIN mem_wstrb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 370.640 477.045 371.240 ;
    END
  END mem_wstrb[3]
  PIN pcpi_insn[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 483.765 277.290 487.765 ;
    END
  END pcpi_insn[0]
  PIN pcpi_insn[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 483.765 254.750 487.765 ;
    END
  END pcpi_insn[10]
  PIN pcpi_insn[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 241.590 483.765 241.870 487.765 ;
    END
  END pcpi_insn[11]
  PIN pcpi_insn[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 401.240 477.045 401.840 ;
    END
  END pcpi_insn[12]
  PIN pcpi_insn[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 418.240 477.045 418.840 ;
    END
  END pcpi_insn[13]
  PIN pcpi_insn[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 376.830 483.765 377.110 487.765 ;
    END
  END pcpi_insn[14]
  PIN pcpi_insn[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END pcpi_insn[15]
  PIN pcpi_insn[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 483.765 113.070 487.765 ;
    END
  END pcpi_insn[16]
  PIN pcpi_insn[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 483.765 80.870 487.765 ;
    END
  END pcpi_insn[17]
  PIN pcpi_insn[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 483.765 183.910 487.765 ;
    END
  END pcpi_insn[18]
  PIN pcpi_insn[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 483.765 196.790 487.765 ;
    END
  END pcpi_insn[19]
  PIN pcpi_insn[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 331.750 483.765 332.030 487.765 ;
    END
  END pcpi_insn[1]
  PIN pcpi_insn[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 483.765 222.550 487.765 ;
    END
  END pcpi_insn[20]
  PIN pcpi_insn[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 483.765 116.290 487.765 ;
    END
  END pcpi_insn[21]
  PIN pcpi_insn[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 483.765 193.570 487.765 ;
    END
  END pcpi_insn[22]
  PIN pcpi_insn[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 483.765 251.530 487.765 ;
    END
  END pcpi_insn[23]
  PIN pcpi_insn[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 257.690 483.765 257.970 487.765 ;
    END
  END pcpi_insn[24]
  PIN pcpi_insn[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 483.765 200.010 487.765 ;
    END
  END pcpi_insn[25]
  PIN pcpi_insn[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 483.765 212.890 487.765 ;
    END
  END pcpi_insn[26]
  PIN pcpi_insn[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 483.765 235.430 487.765 ;
    END
  END pcpi_insn[27]
  PIN pcpi_insn[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 483.765 232.210 487.765 ;
    END
  END pcpi_insn[28]
  PIN pcpi_insn[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 483.765 209.670 487.765 ;
    END
  END pcpi_insn[29]
  PIN pcpi_insn[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 483.765 122.730 487.765 ;
    END
  END pcpi_insn[2]
  PIN pcpi_insn[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 483.765 125.950 487.765 ;
    END
  END pcpi_insn[30]
  PIN pcpi_insn[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 483.765 206.450 487.765 ;
    END
  END pcpi_insn[31]
  PIN pcpi_insn[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 483.765 248.310 487.765 ;
    END
  END pcpi_insn[3]
  PIN pcpi_insn[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 483.765 238.650 487.765 ;
    END
  END pcpi_insn[4]
  PIN pcpi_insn[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 483.765 171.030 487.765 ;
    END
  END pcpi_insn[5]
  PIN pcpi_insn[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 483.765 203.230 487.765 ;
    END
  END pcpi_insn[6]
  PIN pcpi_insn[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 483.765 219.330 487.765 ;
    END
  END pcpi_insn[7]
  PIN pcpi_insn[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 228.710 483.765 228.990 487.765 ;
    END
  END pcpi_insn[8]
  PIN pcpi_insn[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 483.765 245.090 487.765 ;
    END
  END pcpi_insn[9]
  PIN pcpi_rd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END pcpi_rd[0]
  PIN pcpi_rd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END pcpi_rd[10]
  PIN pcpi_rd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END pcpi_rd[11]
  PIN pcpi_rd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END pcpi_rd[12]
  PIN pcpi_rd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END pcpi_rd[13]
  PIN pcpi_rd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END pcpi_rd[14]
  PIN pcpi_rd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END pcpi_rd[15]
  PIN pcpi_rd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END pcpi_rd[16]
  PIN pcpi_rd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END pcpi_rd[17]
  PIN pcpi_rd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END pcpi_rd[18]
  PIN pcpi_rd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END pcpi_rd[19]
  PIN pcpi_rd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END pcpi_rd[1]
  PIN pcpi_rd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END pcpi_rd[20]
  PIN pcpi_rd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END pcpi_rd[21]
  PIN pcpi_rd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END pcpi_rd[22]
  PIN pcpi_rd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END pcpi_rd[23]
  PIN pcpi_rd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END pcpi_rd[24]
  PIN pcpi_rd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END pcpi_rd[25]
  PIN pcpi_rd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END pcpi_rd[26]
  PIN pcpi_rd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END pcpi_rd[27]
  PIN pcpi_rd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END pcpi_rd[28]
  PIN pcpi_rd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END pcpi_rd[29]
  PIN pcpi_rd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END pcpi_rd[2]
  PIN pcpi_rd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END pcpi_rd[30]
  PIN pcpi_rd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END pcpi_rd[31]
  PIN pcpi_rd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END pcpi_rd[3]
  PIN pcpi_rd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END pcpi_rd[4]
  PIN pcpi_rd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END pcpi_rd[5]
  PIN pcpi_rd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END pcpi_rd[6]
  PIN pcpi_rd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END pcpi_rd[7]
  PIN pcpi_rd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END pcpi_rd[8]
  PIN pcpi_rd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END pcpi_rd[9]
  PIN pcpi_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END pcpi_ready
  PIN pcpi_rs1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 431.840 477.045 432.440 ;
    END
  END pcpi_rs1[0]
  PIN pcpi_rs1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 142.840 477.045 143.440 ;
    END
  END pcpi_rs1[10]
  PIN pcpi_rs1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END pcpi_rs1[11]
  PIN pcpi_rs1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END pcpi_rs1[12]
  PIN pcpi_rs1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END pcpi_rs1[13]
  PIN pcpi_rs1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END pcpi_rs1[14]
  PIN pcpi_rs1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END pcpi_rs1[15]
  PIN pcpi_rs1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END pcpi_rs1[16]
  PIN pcpi_rs1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END pcpi_rs1[17]
  PIN pcpi_rs1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END pcpi_rs1[18]
  PIN pcpi_rs1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END pcpi_rs1[19]
  PIN pcpi_rs1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 214.240 477.045 214.840 ;
    END
  END pcpi_rs1[1]
  PIN pcpi_rs1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END pcpi_rs1[20]
  PIN pcpi_rs1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END pcpi_rs1[21]
  PIN pcpi_rs1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END pcpi_rs1[22]
  PIN pcpi_rs1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END pcpi_rs1[23]
  PIN pcpi_rs1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 98.640 477.045 99.240 ;
    END
  END pcpi_rs1[24]
  PIN pcpi_rs1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 105.440 477.045 106.040 ;
    END
  END pcpi_rs1[25]
  PIN pcpi_rs1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 129.240 477.045 129.840 ;
    END
  END pcpi_rs1[26]
  PIN pcpi_rs1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 136.040 477.045 136.640 ;
    END
  END pcpi_rs1[27]
  PIN pcpi_rs1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 187.040 477.045 187.640 ;
    END
  END pcpi_rs1[28]
  PIN pcpi_rs1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 91.840 477.045 92.440 ;
    END
  END pcpi_rs1[29]
  PIN pcpi_rs1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 200.640 477.045 201.240 ;
    END
  END pcpi_rs1[2]
  PIN pcpi_rs1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 61.240 477.045 61.840 ;
    END
  END pcpi_rs1[30]
  PIN pcpi_rs1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 414.840 477.045 415.440 ;
    END
  END pcpi_rs1[31]
  PIN pcpi_rs1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 183.640 477.045 184.240 ;
    END
  END pcpi_rs1[3]
  PIN pcpi_rs1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 180.240 477.045 180.840 ;
    END
  END pcpi_rs1[4]
  PIN pcpi_rs1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 204.040 477.045 204.640 ;
    END
  END pcpi_rs1[5]
  PIN pcpi_rs1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 146.240 477.045 146.840 ;
    END
  END pcpi_rs1[6]
  PIN pcpi_rs1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 156.440 477.045 157.040 ;
    END
  END pcpi_rs1[7]
  PIN pcpi_rs1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 149.640 477.045 150.240 ;
    END
  END pcpi_rs1[8]
  PIN pcpi_rs1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END pcpi_rs1[9]
  PIN pcpi_rs2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 411.440 477.045 412.040 ;
    END
  END pcpi_rs2[0]
  PIN pcpi_rs2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 153.040 477.045 153.640 ;
    END
  END pcpi_rs2[10]
  PIN pcpi_rs2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 139.440 477.045 140.040 ;
    END
  END pcpi_rs2[11]
  PIN pcpi_rs2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 159.840 477.045 160.440 ;
    END
  END pcpi_rs2[12]
  PIN pcpi_rs2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 176.840 477.045 177.440 ;
    END
  END pcpi_rs2[13]
  PIN pcpi_rs2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 193.840 477.045 194.440 ;
    END
  END pcpi_rs2[14]
  PIN pcpi_rs2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 190.440 477.045 191.040 ;
    END
  END pcpi_rs2[15]
  PIN pcpi_rs2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 197.240 477.045 197.840 ;
    END
  END pcpi_rs2[16]
  PIN pcpi_rs2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 163.240 477.045 163.840 ;
    END
  END pcpi_rs2[17]
  PIN pcpi_rs2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 224.440 477.045 225.040 ;
    END
  END pcpi_rs2[18]
  PIN pcpi_rs2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 234.640 477.045 235.240 ;
    END
  END pcpi_rs2[19]
  PIN pcpi_rs2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 346.840 477.045 347.440 ;
    END
  END pcpi_rs2[1]
  PIN pcpi_rs2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 241.440 477.045 242.040 ;
    END
  END pcpi_rs2[20]
  PIN pcpi_rs2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 248.240 477.045 248.840 ;
    END
  END pcpi_rs2[21]
  PIN pcpi_rs2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 81.640 477.045 82.240 ;
    END
  END pcpi_rs2[22]
  PIN pcpi_rs2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 40.840 477.045 41.440 ;
    END
  END pcpi_rs2[23]
  PIN pcpi_rs2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 394.440 477.045 395.040 ;
    END
  END pcpi_rs2[24]
  PIN pcpi_rs2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 333.240 477.045 333.840 ;
    END
  END pcpi_rs2[25]
  PIN pcpi_rs2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 448.840 477.045 449.440 ;
    END
  END pcpi_rs2[26]
  PIN pcpi_rs2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 367.240 477.045 367.840 ;
    END
  END pcpi_rs2[27]
  PIN pcpi_rs2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 374.040 477.045 374.640 ;
    END
  END pcpi_rs2[28]
  PIN pcpi_rs2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 482.840 477.045 483.440 ;
    END
  END pcpi_rs2[29]
  PIN pcpi_rs2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 340.040 477.045 340.640 ;
    END
  END pcpi_rs2[2]
  PIN pcpi_rs2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 452.240 477.045 452.840 ;
    END
  END pcpi_rs2[30]
  PIN pcpi_rs2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 391.040 477.045 391.640 ;
    END
  END pcpi_rs2[31]
  PIN pcpi_rs2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 289.040 477.045 289.640 ;
    END
  END pcpi_rs2[3]
  PIN pcpi_rs2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 384.240 477.045 384.840 ;
    END
  END pcpi_rs2[4]
  PIN pcpi_rs2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 363.840 477.045 364.440 ;
    END
  END pcpi_rs2[5]
  PIN pcpi_rs2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 217.640 477.045 218.240 ;
    END
  END pcpi_rs2[6]
  PIN pcpi_rs2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 238.040 477.045 238.640 ;
    END
  END pcpi_rs2[7]
  PIN pcpi_rs2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 173.440 477.045 174.040 ;
    END
  END pcpi_rs2[8]
  PIN pcpi_rs2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 473.045 166.640 477.045 167.240 ;
    END
  END pcpi_rs2[9]
  PIN pcpi_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 483.765 383.550 487.765 ;
    END
  END pcpi_valid
  PIN pcpi_wait
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END pcpi_wait
  PIN pcpi_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END pcpi_wr
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END resetn
  PIN trace_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 465.840 477.045 466.440 ;
    END
  END trace_data[0]
  PIN trace_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END trace_data[10]
  PIN trace_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END trace_data[11]
  PIN trace_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 17.040 477.045 17.640 ;
    END
  END trace_data[12]
  PIN trace_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END trace_data[13]
  PIN trace_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END trace_data[14]
  PIN trace_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 483.765 344.910 487.765 ;
    END
  END trace_data[15]
  PIN trace_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END trace_data[16]
  PIN trace_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 483.765 460.830 487.765 ;
    END
  END trace_data[17]
  PIN trace_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 483.765 464.050 487.765 ;
    END
  END trace_data[18]
  PIN trace_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 438.640 477.045 439.240 ;
    END
  END trace_data[19]
  PIN trace_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END trace_data[1]
  PIN trace_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END trace_data[20]
  PIN trace_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 483.765 428.630 487.765 ;
    END
  END trace_data[21]
  PIN trace_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END trace_data[22]
  PIN trace_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 483.765 325.590 487.765 ;
    END
  END trace_data[23]
  PIN trace_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 483.765 354.570 487.765 ;
    END
  END trace_data[24]
  PIN trace_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 13.640 477.045 14.240 ;
    END
  END trace_data[25]
  PIN trace_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 473.045 20.440 477.045 21.040 ;
    END
  END trace_data[26]
  PIN trace_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 483.765 393.210 487.765 ;
    END
  END trace_data[27]
  PIN trace_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 483.765 399.650 487.765 ;
    END
  END trace_data[28]
  PIN trace_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END trace_data[29]
  PIN trace_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 483.765 406.090 487.765 ;
    END
  END trace_data[2]
  PIN trace_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 483.765 425.410 487.765 ;
    END
  END trace_data[30]
  PIN trace_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END trace_data[31]
  PIN trace_data[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END trace_data[32]
  PIN trace_data[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 483.765 61.550 487.765 ;
    END
  END trace_data[33]
  PIN trace_data[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END trace_data[34]
  PIN trace_data[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END trace_data[35]
  PIN trace_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END trace_data[3]
  PIN trace_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END trace_data[4]
  PIN trace_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END trace_data[5]
  PIN trace_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 483.765 386.770 487.765 ;
    END
  END trace_data[6]
  PIN trace_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 483.765 447.950 487.765 ;
    END
  END trace_data[7]
  PIN trace_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 483.765 335.250 487.765 ;
    END
  END trace_data[8]
  PIN trace_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 483.765 90.530 487.765 ;
    END
  END trace_data[9]
  PIN trace_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END trace_valid
  PIN trap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 293.110 483.765 293.390 487.765 ;
    END
  END trap
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 471.690 476.190 ;
      LAYER li1 ;
        RECT 5.520 10.795 471.500 476.085 ;
      LAYER met1 ;
        RECT 4.210 10.240 476.030 479.360 ;
      LAYER met2 ;
        RECT 0.550 483.485 38.450 486.725 ;
        RECT 39.290 483.485 60.990 486.725 ;
        RECT 61.830 483.485 64.210 486.725 ;
        RECT 65.050 483.485 67.430 486.725 ;
        RECT 68.270 483.485 70.650 486.725 ;
        RECT 71.490 483.485 73.870 486.725 ;
        RECT 74.710 483.485 77.090 486.725 ;
        RECT 77.930 483.485 80.310 486.725 ;
        RECT 81.150 483.485 83.530 486.725 ;
        RECT 84.370 483.485 86.750 486.725 ;
        RECT 87.590 483.485 89.970 486.725 ;
        RECT 90.810 483.485 93.190 486.725 ;
        RECT 94.030 483.485 96.410 486.725 ;
        RECT 97.250 483.485 99.630 486.725 ;
        RECT 100.470 483.485 102.850 486.725 ;
        RECT 103.690 483.485 106.070 486.725 ;
        RECT 106.910 483.485 109.290 486.725 ;
        RECT 110.130 483.485 112.510 486.725 ;
        RECT 113.350 483.485 115.730 486.725 ;
        RECT 116.570 483.485 118.950 486.725 ;
        RECT 119.790 483.485 122.170 486.725 ;
        RECT 123.010 483.485 125.390 486.725 ;
        RECT 126.230 483.485 128.610 486.725 ;
        RECT 129.450 483.485 131.830 486.725 ;
        RECT 132.670 483.485 135.050 486.725 ;
        RECT 135.890 483.485 138.270 486.725 ;
        RECT 139.110 483.485 141.490 486.725 ;
        RECT 142.330 483.485 144.710 486.725 ;
        RECT 145.550 483.485 147.930 486.725 ;
        RECT 148.770 483.485 151.150 486.725 ;
        RECT 151.990 483.485 154.370 486.725 ;
        RECT 155.210 483.485 157.590 486.725 ;
        RECT 158.430 483.485 160.810 486.725 ;
        RECT 161.650 483.485 164.030 486.725 ;
        RECT 164.870 483.485 167.250 486.725 ;
        RECT 168.090 483.485 170.470 486.725 ;
        RECT 171.310 483.485 173.690 486.725 ;
        RECT 174.530 483.485 176.910 486.725 ;
        RECT 177.750 483.485 180.130 486.725 ;
        RECT 180.970 483.485 183.350 486.725 ;
        RECT 184.190 483.485 186.570 486.725 ;
        RECT 187.410 483.485 189.790 486.725 ;
        RECT 190.630 483.485 193.010 486.725 ;
        RECT 193.850 483.485 196.230 486.725 ;
        RECT 197.070 483.485 199.450 486.725 ;
        RECT 200.290 483.485 202.670 486.725 ;
        RECT 203.510 483.485 205.890 486.725 ;
        RECT 206.730 483.485 209.110 486.725 ;
        RECT 209.950 483.485 212.330 486.725 ;
        RECT 213.170 483.485 215.550 486.725 ;
        RECT 216.390 483.485 218.770 486.725 ;
        RECT 219.610 483.485 221.990 486.725 ;
        RECT 222.830 483.485 225.210 486.725 ;
        RECT 226.050 483.485 228.430 486.725 ;
        RECT 229.270 483.485 231.650 486.725 ;
        RECT 232.490 483.485 234.870 486.725 ;
        RECT 235.710 483.485 238.090 486.725 ;
        RECT 238.930 483.485 241.310 486.725 ;
        RECT 242.150 483.485 244.530 486.725 ;
        RECT 245.370 483.485 247.750 486.725 ;
        RECT 248.590 483.485 250.970 486.725 ;
        RECT 251.810 483.485 254.190 486.725 ;
        RECT 255.030 483.485 257.410 486.725 ;
        RECT 258.250 483.485 260.630 486.725 ;
        RECT 261.470 483.485 263.850 486.725 ;
        RECT 264.690 483.485 267.070 486.725 ;
        RECT 267.910 483.485 270.290 486.725 ;
        RECT 271.130 483.485 273.510 486.725 ;
        RECT 274.350 483.485 276.730 486.725 ;
        RECT 277.570 483.485 279.950 486.725 ;
        RECT 280.790 483.485 283.170 486.725 ;
        RECT 284.010 483.485 286.390 486.725 ;
        RECT 287.230 483.485 289.610 486.725 ;
        RECT 290.450 483.485 292.830 486.725 ;
        RECT 293.670 483.485 296.050 486.725 ;
        RECT 296.890 483.485 299.270 486.725 ;
        RECT 300.110 483.485 302.490 486.725 ;
        RECT 303.330 483.485 305.710 486.725 ;
        RECT 306.550 483.485 308.930 486.725 ;
        RECT 309.770 483.485 312.150 486.725 ;
        RECT 312.990 483.485 315.370 486.725 ;
        RECT 316.210 483.485 318.590 486.725 ;
        RECT 319.430 483.485 321.810 486.725 ;
        RECT 322.650 483.485 325.030 486.725 ;
        RECT 325.870 483.485 328.250 486.725 ;
        RECT 329.090 483.485 331.470 486.725 ;
        RECT 332.310 483.485 334.690 486.725 ;
        RECT 335.530 483.485 337.910 486.725 ;
        RECT 338.750 483.485 341.130 486.725 ;
        RECT 341.970 483.485 344.350 486.725 ;
        RECT 345.190 483.485 347.570 486.725 ;
        RECT 348.410 483.485 350.790 486.725 ;
        RECT 351.630 483.485 354.010 486.725 ;
        RECT 354.850 483.485 357.230 486.725 ;
        RECT 358.070 483.485 360.450 486.725 ;
        RECT 361.290 483.485 363.670 486.725 ;
        RECT 364.510 483.485 366.890 486.725 ;
        RECT 367.730 483.485 370.110 486.725 ;
        RECT 370.950 483.485 373.330 486.725 ;
        RECT 374.170 483.485 376.550 486.725 ;
        RECT 377.390 483.485 379.770 486.725 ;
        RECT 380.610 483.485 382.990 486.725 ;
        RECT 383.830 483.485 386.210 486.725 ;
        RECT 387.050 483.485 389.430 486.725 ;
        RECT 390.270 483.485 392.650 486.725 ;
        RECT 393.490 483.485 395.870 486.725 ;
        RECT 396.710 483.485 399.090 486.725 ;
        RECT 399.930 483.485 402.310 486.725 ;
        RECT 403.150 483.485 405.530 486.725 ;
        RECT 406.370 483.485 408.750 486.725 ;
        RECT 409.590 483.485 411.970 486.725 ;
        RECT 412.810 483.485 415.190 486.725 ;
        RECT 416.030 483.485 418.410 486.725 ;
        RECT 419.250 483.485 421.630 486.725 ;
        RECT 422.470 483.485 424.850 486.725 ;
        RECT 425.690 483.485 428.070 486.725 ;
        RECT 428.910 483.485 431.290 486.725 ;
        RECT 432.130 483.485 434.510 486.725 ;
        RECT 435.350 483.485 444.170 486.725 ;
        RECT 445.010 483.485 447.390 486.725 ;
        RECT 448.230 483.485 460.270 486.725 ;
        RECT 461.110 483.485 463.490 486.725 ;
        RECT 464.330 483.485 476.000 486.725 ;
        RECT 0.550 4.280 476.000 483.485 ;
        RECT 0.650 4.000 3.030 4.280 ;
        RECT 3.870 4.000 6.250 4.280 ;
        RECT 7.090 4.000 9.470 4.280 ;
        RECT 10.310 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 86.750 4.280 ;
        RECT 87.590 4.000 89.970 4.280 ;
        RECT 90.810 4.000 93.190 4.280 ;
        RECT 94.030 4.000 96.410 4.280 ;
        RECT 97.250 4.000 99.630 4.280 ;
        RECT 100.470 4.000 102.850 4.280 ;
        RECT 103.690 4.000 106.070 4.280 ;
        RECT 106.910 4.000 109.290 4.280 ;
        RECT 110.130 4.000 112.510 4.280 ;
        RECT 113.350 4.000 115.730 4.280 ;
        RECT 116.570 4.000 118.950 4.280 ;
        RECT 119.790 4.000 122.170 4.280 ;
        RECT 123.010 4.000 125.390 4.280 ;
        RECT 126.230 4.000 128.610 4.280 ;
        RECT 129.450 4.000 131.830 4.280 ;
        RECT 132.670 4.000 135.050 4.280 ;
        RECT 135.890 4.000 138.270 4.280 ;
        RECT 139.110 4.000 141.490 4.280 ;
        RECT 142.330 4.000 144.710 4.280 ;
        RECT 145.550 4.000 147.930 4.280 ;
        RECT 148.770 4.000 151.150 4.280 ;
        RECT 151.990 4.000 154.370 4.280 ;
        RECT 155.210 4.000 157.590 4.280 ;
        RECT 158.430 4.000 160.810 4.280 ;
        RECT 161.650 4.000 164.030 4.280 ;
        RECT 164.870 4.000 167.250 4.280 ;
        RECT 168.090 4.000 170.470 4.280 ;
        RECT 171.310 4.000 173.690 4.280 ;
        RECT 174.530 4.000 176.910 4.280 ;
        RECT 177.750 4.000 180.130 4.280 ;
        RECT 180.970 4.000 183.350 4.280 ;
        RECT 184.190 4.000 186.570 4.280 ;
        RECT 187.410 4.000 189.790 4.280 ;
        RECT 190.630 4.000 193.010 4.280 ;
        RECT 193.850 4.000 196.230 4.280 ;
        RECT 197.070 4.000 199.450 4.280 ;
        RECT 200.290 4.000 202.670 4.280 ;
        RECT 203.510 4.000 205.890 4.280 ;
        RECT 206.730 4.000 209.110 4.280 ;
        RECT 209.950 4.000 212.330 4.280 ;
        RECT 213.170 4.000 215.550 4.280 ;
        RECT 216.390 4.000 218.770 4.280 ;
        RECT 219.610 4.000 221.990 4.280 ;
        RECT 222.830 4.000 225.210 4.280 ;
        RECT 226.050 4.000 228.430 4.280 ;
        RECT 229.270 4.000 231.650 4.280 ;
        RECT 232.490 4.000 234.870 4.280 ;
        RECT 235.710 4.000 238.090 4.280 ;
        RECT 238.930 4.000 241.310 4.280 ;
        RECT 242.150 4.000 244.530 4.280 ;
        RECT 245.370 4.000 247.750 4.280 ;
        RECT 248.590 4.000 250.970 4.280 ;
        RECT 251.810 4.000 254.190 4.280 ;
        RECT 255.030 4.000 257.410 4.280 ;
        RECT 258.250 4.000 260.630 4.280 ;
        RECT 261.470 4.000 263.850 4.280 ;
        RECT 264.690 4.000 267.070 4.280 ;
        RECT 267.910 4.000 270.290 4.280 ;
        RECT 271.130 4.000 273.510 4.280 ;
        RECT 274.350 4.000 276.730 4.280 ;
        RECT 277.570 4.000 279.950 4.280 ;
        RECT 280.790 4.000 283.170 4.280 ;
        RECT 284.010 4.000 286.390 4.280 ;
        RECT 287.230 4.000 289.610 4.280 ;
        RECT 290.450 4.000 292.830 4.280 ;
        RECT 293.670 4.000 296.050 4.280 ;
        RECT 296.890 4.000 299.270 4.280 ;
        RECT 300.110 4.000 302.490 4.280 ;
        RECT 303.330 4.000 305.710 4.280 ;
        RECT 306.550 4.000 308.930 4.280 ;
        RECT 309.770 4.000 312.150 4.280 ;
        RECT 312.990 4.000 315.370 4.280 ;
        RECT 316.210 4.000 318.590 4.280 ;
        RECT 319.430 4.000 321.810 4.280 ;
        RECT 322.650 4.000 325.030 4.280 ;
        RECT 325.870 4.000 328.250 4.280 ;
        RECT 329.090 4.000 331.470 4.280 ;
        RECT 332.310 4.000 334.690 4.280 ;
        RECT 335.530 4.000 337.910 4.280 ;
        RECT 338.750 4.000 341.130 4.280 ;
        RECT 341.970 4.000 344.350 4.280 ;
        RECT 345.190 4.000 347.570 4.280 ;
        RECT 348.410 4.000 350.790 4.280 ;
        RECT 351.630 4.000 389.430 4.280 ;
        RECT 390.270 4.000 392.650 4.280 ;
        RECT 393.490 4.000 418.410 4.280 ;
        RECT 419.250 4.000 421.630 4.280 ;
        RECT 422.470 4.000 424.850 4.280 ;
        RECT 425.690 4.000 437.730 4.280 ;
        RECT 438.570 4.000 453.830 4.280 ;
        RECT 454.670 4.000 476.000 4.280 ;
      LAYER met3 ;
        RECT 0.525 485.840 472.645 486.705 ;
        RECT 0.525 483.840 475.575 485.840 ;
        RECT 0.525 482.440 472.645 483.840 ;
        RECT 0.525 480.440 475.575 482.440 ;
        RECT 0.525 479.040 472.645 480.440 ;
        RECT 0.525 477.040 475.575 479.040 ;
        RECT 0.525 475.640 472.645 477.040 ;
        RECT 0.525 473.640 475.575 475.640 ;
        RECT 0.525 472.240 472.645 473.640 ;
        RECT 0.525 470.240 475.575 472.240 ;
        RECT 4.400 468.840 472.645 470.240 ;
        RECT 0.525 466.840 475.575 468.840 ;
        RECT 4.400 465.440 472.645 466.840 ;
        RECT 0.525 463.440 475.575 465.440 ;
        RECT 0.525 462.040 472.645 463.440 ;
        RECT 0.525 460.040 475.575 462.040 ;
        RECT 4.400 458.640 472.645 460.040 ;
        RECT 0.525 456.640 475.575 458.640 ;
        RECT 0.525 455.240 472.645 456.640 ;
        RECT 0.525 453.240 475.575 455.240 ;
        RECT 0.525 451.840 472.645 453.240 ;
        RECT 0.525 449.840 475.575 451.840 ;
        RECT 0.525 448.440 472.645 449.840 ;
        RECT 0.525 446.440 475.575 448.440 ;
        RECT 0.525 445.040 472.645 446.440 ;
        RECT 0.525 443.040 475.575 445.040 ;
        RECT 0.525 441.640 472.645 443.040 ;
        RECT 0.525 439.640 475.575 441.640 ;
        RECT 0.525 438.240 472.645 439.640 ;
        RECT 0.525 436.240 475.575 438.240 ;
        RECT 0.525 434.840 472.645 436.240 ;
        RECT 0.525 432.840 475.575 434.840 ;
        RECT 0.525 431.440 472.645 432.840 ;
        RECT 0.525 429.440 475.575 431.440 ;
        RECT 0.525 428.040 472.645 429.440 ;
        RECT 0.525 426.040 475.575 428.040 ;
        RECT 0.525 424.640 472.645 426.040 ;
        RECT 0.525 422.640 475.575 424.640 ;
        RECT 0.525 421.240 472.645 422.640 ;
        RECT 0.525 419.240 475.575 421.240 ;
        RECT 0.525 417.840 472.645 419.240 ;
        RECT 0.525 415.840 475.575 417.840 ;
        RECT 0.525 414.440 472.645 415.840 ;
        RECT 0.525 412.440 475.575 414.440 ;
        RECT 0.525 411.040 472.645 412.440 ;
        RECT 0.525 409.040 475.575 411.040 ;
        RECT 0.525 407.640 472.645 409.040 ;
        RECT 0.525 405.640 475.575 407.640 ;
        RECT 0.525 404.240 472.645 405.640 ;
        RECT 0.525 402.240 475.575 404.240 ;
        RECT 0.525 400.840 472.645 402.240 ;
        RECT 0.525 398.840 475.575 400.840 ;
        RECT 0.525 397.440 472.645 398.840 ;
        RECT 0.525 395.440 475.575 397.440 ;
        RECT 0.525 394.040 472.645 395.440 ;
        RECT 0.525 392.040 475.575 394.040 ;
        RECT 0.525 390.640 472.645 392.040 ;
        RECT 0.525 388.640 475.575 390.640 ;
        RECT 0.525 387.240 472.645 388.640 ;
        RECT 0.525 385.240 475.575 387.240 ;
        RECT 0.525 383.840 472.645 385.240 ;
        RECT 0.525 381.840 475.575 383.840 ;
        RECT 0.525 380.440 472.645 381.840 ;
        RECT 0.525 378.440 475.575 380.440 ;
        RECT 0.525 377.040 472.645 378.440 ;
        RECT 0.525 375.040 475.575 377.040 ;
        RECT 0.525 373.640 472.645 375.040 ;
        RECT 0.525 371.640 475.575 373.640 ;
        RECT 0.525 370.240 472.645 371.640 ;
        RECT 0.525 368.240 475.575 370.240 ;
        RECT 0.525 366.840 472.645 368.240 ;
        RECT 0.525 364.840 475.575 366.840 ;
        RECT 0.525 363.440 472.645 364.840 ;
        RECT 0.525 361.440 475.575 363.440 ;
        RECT 0.525 360.040 472.645 361.440 ;
        RECT 0.525 358.040 475.575 360.040 ;
        RECT 0.525 356.640 472.645 358.040 ;
        RECT 0.525 354.640 475.575 356.640 ;
        RECT 0.525 353.240 472.645 354.640 ;
        RECT 0.525 351.240 475.575 353.240 ;
        RECT 0.525 349.840 472.645 351.240 ;
        RECT 0.525 347.840 475.575 349.840 ;
        RECT 0.525 346.440 472.645 347.840 ;
        RECT 0.525 344.440 475.575 346.440 ;
        RECT 0.525 343.040 472.645 344.440 ;
        RECT 0.525 341.040 475.575 343.040 ;
        RECT 0.525 339.640 472.645 341.040 ;
        RECT 0.525 337.640 475.575 339.640 ;
        RECT 0.525 336.240 472.645 337.640 ;
        RECT 0.525 334.240 475.575 336.240 ;
        RECT 0.525 332.840 472.645 334.240 ;
        RECT 0.525 330.840 475.575 332.840 ;
        RECT 0.525 329.440 472.645 330.840 ;
        RECT 0.525 327.440 475.575 329.440 ;
        RECT 0.525 326.040 472.645 327.440 ;
        RECT 0.525 324.040 475.575 326.040 ;
        RECT 0.525 322.640 472.645 324.040 ;
        RECT 0.525 320.640 475.575 322.640 ;
        RECT 0.525 319.240 472.645 320.640 ;
        RECT 0.525 317.240 475.575 319.240 ;
        RECT 0.525 315.840 472.645 317.240 ;
        RECT 0.525 313.840 475.575 315.840 ;
        RECT 0.525 312.440 472.645 313.840 ;
        RECT 0.525 310.440 475.575 312.440 ;
        RECT 0.525 309.040 472.645 310.440 ;
        RECT 0.525 307.040 475.575 309.040 ;
        RECT 0.525 305.640 472.645 307.040 ;
        RECT 0.525 303.640 475.575 305.640 ;
        RECT 0.525 302.240 472.645 303.640 ;
        RECT 0.525 300.240 475.575 302.240 ;
        RECT 0.525 298.840 472.645 300.240 ;
        RECT 0.525 296.840 475.575 298.840 ;
        RECT 0.525 295.440 472.645 296.840 ;
        RECT 0.525 293.440 475.575 295.440 ;
        RECT 0.525 292.040 472.645 293.440 ;
        RECT 0.525 290.040 475.575 292.040 ;
        RECT 4.400 288.640 472.645 290.040 ;
        RECT 0.525 286.640 475.575 288.640 ;
        RECT 4.400 285.240 472.645 286.640 ;
        RECT 0.525 283.240 475.575 285.240 ;
        RECT 0.525 281.840 472.645 283.240 ;
        RECT 0.525 279.840 475.575 281.840 ;
        RECT 0.525 278.440 472.645 279.840 ;
        RECT 0.525 276.440 475.575 278.440 ;
        RECT 0.525 275.040 472.645 276.440 ;
        RECT 0.525 273.040 475.575 275.040 ;
        RECT 0.525 271.640 472.645 273.040 ;
        RECT 0.525 269.640 475.575 271.640 ;
        RECT 0.525 268.240 472.645 269.640 ;
        RECT 0.525 266.240 475.575 268.240 ;
        RECT 4.400 264.840 472.645 266.240 ;
        RECT 0.525 262.840 475.575 264.840 ;
        RECT 4.400 261.440 472.645 262.840 ;
        RECT 0.525 259.440 475.575 261.440 ;
        RECT 4.400 258.040 472.645 259.440 ;
        RECT 0.525 256.040 475.575 258.040 ;
        RECT 0.525 254.640 472.645 256.040 ;
        RECT 0.525 252.640 475.575 254.640 ;
        RECT 0.525 251.240 472.645 252.640 ;
        RECT 0.525 249.240 475.575 251.240 ;
        RECT 4.400 247.840 472.645 249.240 ;
        RECT 0.525 245.840 475.575 247.840 ;
        RECT 4.400 244.440 472.645 245.840 ;
        RECT 0.525 242.440 475.575 244.440 ;
        RECT 0.525 241.040 472.645 242.440 ;
        RECT 0.525 239.040 475.575 241.040 ;
        RECT 0.525 237.640 472.645 239.040 ;
        RECT 0.525 235.640 475.575 237.640 ;
        RECT 4.400 234.240 472.645 235.640 ;
        RECT 0.525 232.240 475.575 234.240 ;
        RECT 4.400 230.840 472.645 232.240 ;
        RECT 0.525 228.840 475.575 230.840 ;
        RECT 0.525 227.440 472.645 228.840 ;
        RECT 0.525 225.440 475.575 227.440 ;
        RECT 0.525 224.040 472.645 225.440 ;
        RECT 0.525 222.040 475.575 224.040 ;
        RECT 4.400 220.640 472.645 222.040 ;
        RECT 0.525 218.640 475.575 220.640 ;
        RECT 4.400 217.240 472.645 218.640 ;
        RECT 0.525 215.240 475.575 217.240 ;
        RECT 0.525 213.840 472.645 215.240 ;
        RECT 0.525 211.840 475.575 213.840 ;
        RECT 4.400 210.440 472.645 211.840 ;
        RECT 0.525 208.440 475.575 210.440 ;
        RECT 4.400 207.040 472.645 208.440 ;
        RECT 0.525 205.040 475.575 207.040 ;
        RECT 0.525 203.640 472.645 205.040 ;
        RECT 0.525 201.640 475.575 203.640 ;
        RECT 0.525 200.240 472.645 201.640 ;
        RECT 0.525 198.240 475.575 200.240 ;
        RECT 0.525 196.840 472.645 198.240 ;
        RECT 0.525 194.840 475.575 196.840 ;
        RECT 0.525 193.440 472.645 194.840 ;
        RECT 0.525 191.440 475.575 193.440 ;
        RECT 0.525 190.040 472.645 191.440 ;
        RECT 0.525 188.040 475.575 190.040 ;
        RECT 0.525 186.640 472.645 188.040 ;
        RECT 0.525 184.640 475.575 186.640 ;
        RECT 0.525 183.240 472.645 184.640 ;
        RECT 0.525 181.240 475.575 183.240 ;
        RECT 0.525 179.840 472.645 181.240 ;
        RECT 0.525 177.840 475.575 179.840 ;
        RECT 0.525 176.440 472.645 177.840 ;
        RECT 0.525 174.440 475.575 176.440 ;
        RECT 0.525 173.040 472.645 174.440 ;
        RECT 0.525 171.040 475.575 173.040 ;
        RECT 0.525 169.640 472.645 171.040 ;
        RECT 0.525 167.640 475.575 169.640 ;
        RECT 0.525 166.240 472.645 167.640 ;
        RECT 0.525 164.240 475.575 166.240 ;
        RECT 0.525 162.840 472.645 164.240 ;
        RECT 0.525 160.840 475.575 162.840 ;
        RECT 0.525 159.440 472.645 160.840 ;
        RECT 0.525 157.440 475.575 159.440 ;
        RECT 0.525 156.040 472.645 157.440 ;
        RECT 0.525 154.040 475.575 156.040 ;
        RECT 0.525 152.640 472.645 154.040 ;
        RECT 0.525 150.640 475.575 152.640 ;
        RECT 0.525 149.240 472.645 150.640 ;
        RECT 0.525 147.240 475.575 149.240 ;
        RECT 0.525 145.840 472.645 147.240 ;
        RECT 0.525 143.840 475.575 145.840 ;
        RECT 0.525 142.440 472.645 143.840 ;
        RECT 0.525 140.440 475.575 142.440 ;
        RECT 0.525 139.040 472.645 140.440 ;
        RECT 0.525 137.040 475.575 139.040 ;
        RECT 0.525 135.640 472.645 137.040 ;
        RECT 0.525 133.640 475.575 135.640 ;
        RECT 0.525 132.240 472.645 133.640 ;
        RECT 0.525 130.240 475.575 132.240 ;
        RECT 0.525 128.840 472.645 130.240 ;
        RECT 0.525 126.840 475.575 128.840 ;
        RECT 0.525 125.440 472.645 126.840 ;
        RECT 0.525 123.440 475.575 125.440 ;
        RECT 0.525 122.040 472.645 123.440 ;
        RECT 0.525 120.040 475.575 122.040 ;
        RECT 0.525 118.640 472.645 120.040 ;
        RECT 0.525 116.640 475.575 118.640 ;
        RECT 0.525 115.240 472.645 116.640 ;
        RECT 0.525 113.240 475.575 115.240 ;
        RECT 0.525 111.840 472.645 113.240 ;
        RECT 0.525 109.840 475.575 111.840 ;
        RECT 0.525 108.440 472.645 109.840 ;
        RECT 0.525 106.440 475.575 108.440 ;
        RECT 0.525 105.040 472.645 106.440 ;
        RECT 0.525 103.040 475.575 105.040 ;
        RECT 0.525 101.640 472.645 103.040 ;
        RECT 0.525 99.640 475.575 101.640 ;
        RECT 0.525 98.240 472.645 99.640 ;
        RECT 0.525 96.240 475.575 98.240 ;
        RECT 0.525 94.840 472.645 96.240 ;
        RECT 0.525 92.840 475.575 94.840 ;
        RECT 0.525 91.440 472.645 92.840 ;
        RECT 0.525 89.440 475.575 91.440 ;
        RECT 0.525 88.040 472.645 89.440 ;
        RECT 0.525 86.040 475.575 88.040 ;
        RECT 0.525 84.640 472.645 86.040 ;
        RECT 0.525 82.640 475.575 84.640 ;
        RECT 0.525 81.240 472.645 82.640 ;
        RECT 0.525 79.240 475.575 81.240 ;
        RECT 0.525 77.840 472.645 79.240 ;
        RECT 0.525 75.840 475.575 77.840 ;
        RECT 0.525 74.440 472.645 75.840 ;
        RECT 0.525 72.440 475.575 74.440 ;
        RECT 0.525 71.040 472.645 72.440 ;
        RECT 0.525 69.040 475.575 71.040 ;
        RECT 0.525 67.640 472.645 69.040 ;
        RECT 0.525 65.640 475.575 67.640 ;
        RECT 4.400 64.240 472.645 65.640 ;
        RECT 0.525 62.240 475.575 64.240 ;
        RECT 0.525 60.840 472.645 62.240 ;
        RECT 0.525 58.840 475.575 60.840 ;
        RECT 0.525 57.440 472.645 58.840 ;
        RECT 0.525 55.440 475.575 57.440 ;
        RECT 4.400 54.040 472.645 55.440 ;
        RECT 0.525 52.040 475.575 54.040 ;
        RECT 4.400 50.640 472.645 52.040 ;
        RECT 0.525 48.640 475.575 50.640 ;
        RECT 0.525 47.240 472.645 48.640 ;
        RECT 0.525 45.240 475.575 47.240 ;
        RECT 4.400 43.840 472.645 45.240 ;
        RECT 0.525 41.840 475.575 43.840 ;
        RECT 4.400 40.440 472.645 41.840 ;
        RECT 0.525 38.440 475.575 40.440 ;
        RECT 4.400 37.040 472.645 38.440 ;
        RECT 0.525 35.040 475.575 37.040 ;
        RECT 4.400 33.640 472.645 35.040 ;
        RECT 0.525 31.640 475.575 33.640 ;
        RECT 0.525 30.240 472.645 31.640 ;
        RECT 0.525 28.240 475.575 30.240 ;
        RECT 4.400 26.840 472.645 28.240 ;
        RECT 0.525 24.840 475.575 26.840 ;
        RECT 4.400 23.440 475.575 24.840 ;
        RECT 0.525 21.440 475.575 23.440 ;
        RECT 4.400 20.040 472.645 21.440 ;
        RECT 0.525 18.040 475.575 20.040 ;
        RECT 4.400 16.640 472.645 18.040 ;
        RECT 0.525 14.640 475.575 16.640 ;
        RECT 4.400 13.240 472.645 14.640 ;
        RECT 0.525 11.240 475.575 13.240 ;
        RECT 4.400 9.840 472.645 11.240 ;
        RECT 0.525 7.840 475.575 9.840 ;
        RECT 4.400 6.975 475.575 7.840 ;
      LAYER met4 ;
        RECT 23.295 19.895 23.940 474.465 ;
        RECT 26.340 19.895 174.240 474.465 ;
        RECT 176.640 19.895 177.540 474.465 ;
        RECT 179.940 19.895 327.840 474.465 ;
        RECT 330.240 19.895 331.140 474.465 ;
        RECT 333.540 19.895 469.825 474.465 ;
      LAYER met5 ;
        RECT 122.940 364.700 367.420 373.100 ;
  END
END picorv32
END LIBRARY

