* NGSPICE file created from picorv32.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt picorv32 VGND VPWR clk eoi[0] eoi[10] eoi[11] eoi[12] eoi[13] eoi[14] eoi[15]
+ eoi[16] eoi[17] eoi[18] eoi[19] eoi[1] eoi[20] eoi[21] eoi[22] eoi[23] eoi[24] eoi[25]
+ eoi[26] eoi[27] eoi[28] eoi[29] eoi[2] eoi[30] eoi[31] eoi[3] eoi[4] eoi[5] eoi[6]
+ eoi[7] eoi[8] eoi[9] irq[0] irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[16]
+ irq[17] irq[18] irq[19] irq[1] irq[20] irq[21] irq[22] irq[23] irq[24] irq[25] irq[26]
+ irq[27] irq[28] irq[29] irq[2] irq[30] irq[31] irq[3] irq[4] irq[5] irq[6] irq[7]
+ irq[8] irq[9] mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12] mem_addr[13] mem_addr[14]
+ mem_addr[15] mem_addr[16] mem_addr[17] mem_addr[18] mem_addr[19] mem_addr[1] mem_addr[20]
+ mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[24] mem_addr[25] mem_addr[26] mem_addr[27]
+ mem_addr[28] mem_addr[29] mem_addr[2] mem_addr[30] mem_addr[31] mem_addr[3] mem_addr[4]
+ mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_instr mem_la_addr[0]
+ mem_la_addr[10] mem_la_addr[11] mem_la_addr[12] mem_la_addr[13] mem_la_addr[14]
+ mem_la_addr[15] mem_la_addr[16] mem_la_addr[17] mem_la_addr[18] mem_la_addr[19]
+ mem_la_addr[1] mem_la_addr[20] mem_la_addr[21] mem_la_addr[22] mem_la_addr[23] mem_la_addr[24]
+ mem_la_addr[25] mem_la_addr[26] mem_la_addr[27] mem_la_addr[28] mem_la_addr[29]
+ mem_la_addr[2] mem_la_addr[30] mem_la_addr[31] mem_la_addr[3] mem_la_addr[4] mem_la_addr[5]
+ mem_la_addr[6] mem_la_addr[7] mem_la_addr[8] mem_la_addr[9] mem_la_read mem_la_wdata[0]
+ mem_la_wdata[10] mem_la_wdata[11] mem_la_wdata[12] mem_la_wdata[13] mem_la_wdata[14]
+ mem_la_wdata[15] mem_la_wdata[16] mem_la_wdata[17] mem_la_wdata[18] mem_la_wdata[19]
+ mem_la_wdata[1] mem_la_wdata[20] mem_la_wdata[21] mem_la_wdata[22] mem_la_wdata[23]
+ mem_la_wdata[24] mem_la_wdata[25] mem_la_wdata[26] mem_la_wdata[27] mem_la_wdata[28]
+ mem_la_wdata[29] mem_la_wdata[2] mem_la_wdata[30] mem_la_wdata[31] mem_la_wdata[3]
+ mem_la_wdata[4] mem_la_wdata[5] mem_la_wdata[6] mem_la_wdata[7] mem_la_wdata[8]
+ mem_la_wdata[9] mem_la_write mem_la_wstrb[0] mem_la_wstrb[1] mem_la_wstrb[2] mem_la_wstrb[3]
+ mem_rdata[0] mem_rdata[10] mem_rdata[11] mem_rdata[12] mem_rdata[13] mem_rdata[14]
+ mem_rdata[15] mem_rdata[16] mem_rdata[17] mem_rdata[18] mem_rdata[19] mem_rdata[1]
+ mem_rdata[20] mem_rdata[21] mem_rdata[22] mem_rdata[23] mem_rdata[24] mem_rdata[25]
+ mem_rdata[26] mem_rdata[27] mem_rdata[28] mem_rdata[29] mem_rdata[2] mem_rdata[30]
+ mem_rdata[31] mem_rdata[3] mem_rdata[4] mem_rdata[5] mem_rdata[6] mem_rdata[7] mem_rdata[8]
+ mem_rdata[9] mem_ready mem_valid mem_wdata[0] mem_wdata[10] mem_wdata[11] mem_wdata[12]
+ mem_wdata[13] mem_wdata[14] mem_wdata[15] mem_wdata[16] mem_wdata[17] mem_wdata[18]
+ mem_wdata[19] mem_wdata[1] mem_wdata[20] mem_wdata[21] mem_wdata[22] mem_wdata[23]
+ mem_wdata[24] mem_wdata[25] mem_wdata[26] mem_wdata[27] mem_wdata[28] mem_wdata[29]
+ mem_wdata[2] mem_wdata[30] mem_wdata[31] mem_wdata[3] mem_wdata[4] mem_wdata[5]
+ mem_wdata[6] mem_wdata[7] mem_wdata[8] mem_wdata[9] mem_wstrb[0] mem_wstrb[1] mem_wstrb[2]
+ mem_wstrb[3] pcpi_insn[0] pcpi_insn[10] pcpi_insn[11] pcpi_insn[12] pcpi_insn[13]
+ pcpi_insn[14] pcpi_insn[15] pcpi_insn[16] pcpi_insn[17] pcpi_insn[18] pcpi_insn[19]
+ pcpi_insn[1] pcpi_insn[20] pcpi_insn[21] pcpi_insn[22] pcpi_insn[23] pcpi_insn[24]
+ pcpi_insn[25] pcpi_insn[26] pcpi_insn[27] pcpi_insn[28] pcpi_insn[29] pcpi_insn[2]
+ pcpi_insn[30] pcpi_insn[31] pcpi_insn[3] pcpi_insn[4] pcpi_insn[5] pcpi_insn[6]
+ pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_rd[0] pcpi_rd[10] pcpi_rd[11] pcpi_rd[12]
+ pcpi_rd[13] pcpi_rd[14] pcpi_rd[15] pcpi_rd[16] pcpi_rd[17] pcpi_rd[18] pcpi_rd[19]
+ pcpi_rd[1] pcpi_rd[20] pcpi_rd[21] pcpi_rd[22] pcpi_rd[23] pcpi_rd[24] pcpi_rd[25]
+ pcpi_rd[26] pcpi_rd[27] pcpi_rd[28] pcpi_rd[29] pcpi_rd[2] pcpi_rd[30] pcpi_rd[31]
+ pcpi_rd[3] pcpi_rd[4] pcpi_rd[5] pcpi_rd[6] pcpi_rd[7] pcpi_rd[8] pcpi_rd[9] pcpi_ready
+ pcpi_rs1[0] pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14] pcpi_rs1[15]
+ pcpi_rs1[16] pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20] pcpi_rs1[21]
+ pcpi_rs1[22] pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27] pcpi_rs1[28]
+ pcpi_rs1[29] pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4] pcpi_rs1[5]
+ pcpi_rs1[6] pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10] pcpi_rs2[11]
+ pcpi_rs2[12] pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17] pcpi_rs2[18]
+ pcpi_rs2[19] pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23] pcpi_rs2[24]
+ pcpi_rs2[25] pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2] pcpi_rs2[30]
+ pcpi_rs2[31] pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7] pcpi_rs2[8]
+ pcpi_rs2[9] pcpi_valid pcpi_wait pcpi_wr resetn trace_data[0] trace_data[10] trace_data[11]
+ trace_data[12] trace_data[13] trace_data[14] trace_data[15] trace_data[16] trace_data[17]
+ trace_data[18] trace_data[19] trace_data[1] trace_data[20] trace_data[21] trace_data[22]
+ trace_data[23] trace_data[24] trace_data[25] trace_data[26] trace_data[27] trace_data[28]
+ trace_data[29] trace_data[2] trace_data[30] trace_data[31] trace_data[32] trace_data[33]
+ trace_data[34] trace_data[35] trace_data[3] trace_data[4] trace_data[5] trace_data[6]
+ trace_data[7] trace_data[8] trace_data[9] trace_valid trap
XFILLER_67_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06883_ net850 _02480_ _02478_ _02472_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__a211o_1
X_09671_ _04460_ _02479_ net848 _04424_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_143_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08622_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__inv_2
XANTENNA__09304__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08553_ genblk1.genblk1.pcpi_mul.next_rs2\[12\] net1091 genblk1.genblk1.pcpi_mul.rd\[11\]
+ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__a21o_1
XANTENNA__09287__A1 _03844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07504_ _02983_ _02995_ _03031_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__o31a_1
X_08484_ genblk1.genblk1.pcpi_mul.rd\[0\] genblk1.genblk1.pcpi_mul.next_rs2\[1\] net1101
+ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_18_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07435_ count_instr\[51\] net1132 net1142 count_cycle\[51\] VGND VGND VPWR VPWR _02969_
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1071_A net1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1169_A net1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12043__B1 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07366_ net1071 _02895_ _02896_ _02904_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__a31o_1
XANTENNA__13240__C1 net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09105_ net1840 net354 net505 VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__mux2_1
XANTENNA__11141__Y _05820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09995__C1 _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07297_ _02811_ _02839_ net1060 VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__o21a_1
XFILLER_164_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09036_ net408 net2513 net513 VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__mux2_1
XANTENNA__07470__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout796_A net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11149__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13496__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold340 cpuregs\[29\]\[27\] VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08014__A2 net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1124_X net1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold351 cpuregs\[8\]\[21\] VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold362 genblk1.genblk1.pcpi_mul.pcpi_rd\[19\] VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 cpuregs\[31\]\[18\] VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold384 cpuregs\[10\]\[21\] VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout963_A net965 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold395 cpuregs\[16\]\[17\] VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 net821 VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout831 net834 VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__clkbuf_4
X_09938_ net3017 net879 _04710_ _04714_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__a22o_1
XANTENNA__10109__B1 net1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout842 _02702_ VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__buf_2
Xfanout853 net854 VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__buf_2
Xfanout864 net865 VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout875 net876 VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__buf_2
Xfanout886 net891 VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__buf_2
XANTENNA_fanout751_X net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09869_ net1128 _04441_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__nand2_1
Xfanout897 net898 VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__clkbuf_4
Xhold1040 cpuregs\[11\]\[17\] VGND VGND VPWR VPWR net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout849_X net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11321__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11744__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1051 cpuregs\[7\]\[16\] VGND VGND VPWR VPWR net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _01423_ VGND VGND VPWR VPWR net2376 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ genblk2.pcpi_div.divisor\[27\] genblk2.pcpi_div.dividend\[27\] VGND VGND
+ VPWR VPWR _06371_ sky130_fd_sc_hd__nand2b_1
X_12880_ mem_rdata_q\[17\] net9 net962 VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__mux2_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1073 cpuregs\[2\]\[7\] VGND VGND VPWR VPWR net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 instr_fence VGND VGND VPWR VPWR net2398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09214__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1095 genblk1.genblk1.pcpi_mul.next_rs1\[1\] VGND VGND VPWR VPWR net2409 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ genblk2.pcpi_div.dividend\[11\] genblk2.pcpi_div.divisor\[11\] VGND VGND
+ VPWR VPWR _06302_ sky130_fd_sc_hd__and2b_1
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14550_ clknet_leaf_187_clk _00936_ VGND VGND VPWR VPWR cpuregs\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ net2698 net116 net729 VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__mux2_1
XANTENNA__11085__B2 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13501_ net1519 net348 net419 VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__mux2_1
X_10713_ net789 _05398_ _05400_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__or4_1
X_14481_ clknet_leaf_95_clk _00870_ VGND VGND VPWR VPWR instr_sh sky130_fd_sc_hd__dfxtp_1
XANTENNA__12575__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11693_ net1859 net409 net373 VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13432_ net1188 _04883_ net760 VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__a21o_1
XFILLER_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10644_ cpuregs\[28\]\[8\] cpuregs\[29\]\[8\] net670 VGND VGND VPWR VPWR _05336_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10575_ cpuregs\[22\]\[6\] cpuregs\[23\]\[6\] net671 VGND VGND VPWR VPWR _05269_
+ sky130_fd_sc_hd__mux2_1
X_13363_ net958 _05008_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__and3_1
XFILLER_154_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15102_ clknet_leaf_15_clk _01454_ VGND VGND VPWR VPWR cpuregs\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12314_ net1146 decoded_imm_j\[16\] net970 mem_rdata_q\[16\] VGND VGND VPWR VPWR
+ _06636_ sky130_fd_sc_hd__a22o_1
X_13294_ _04928_ _04978_ _04982_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__and3_1
XANTENNA__12337__A1 decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12337__B2 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15033_ clknet_leaf_136_clk net1327 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_12245_ genblk2.pcpi_div.divisor\[8\] net379 net366 net2661 VGND VGND VPWR VPWR _01114_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10348__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14799__Q decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ net751 net3000 VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__nor2_1
X_11127_ cpuregs\[24\]\[21\] net658 VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11058_ cpuregs\[30\]\[19\] cpuregs\[31\]\[19\] net681 VGND VGND VPWR VPWR _05739_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07516__A1 net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11654__S net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13435__A is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10009_ count_cycle\[4\] _04771_ count_cycle\[5\] VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__a21o_1
XFILLER_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10520__B1 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09124__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14817_ clknet_leaf_79_clk _01169_ VGND VGND VPWR VPWR decoded_imm\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14748_ clknet_leaf_157_clk _01133_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08963__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14679_ clknet_leaf_153_clk _01064_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14369__CLK clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07220_ count_instr\[37\] net1130 net1135 count_instr\[5\] VGND VGND VPWR VPWR _02768_
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12025__B1 net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07151_ count_cycle\[0\] net975 VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__or2_1
XFILLER_158_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11402__B net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07082_ net1121 _02644_ net2766 VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_35_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__B2 net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11542__A_N net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07984_ _03311_ _03496_ net771 VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__o21ai_1
X_09723_ _04427_ _04428_ _04488_ _04429_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__a31o_1
X_06935_ genblk2.pcpi_div.dividend\[2\] _02518_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout377_A net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09654_ _04422_ _04453_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__or2_1
XFILLER_95_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06866_ instr_lw net410 _02460_ instr_sw net850 VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__a221o_1
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09034__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08605_ genblk1.genblk1.pcpi_mul.next_rs2\[20\] net1098 genblk1.genblk1.pcpi_mul.rd\[19\]
+ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__a21o_1
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09585_ net2865 _04417_ net1238 VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__o21ai_1
X_06797_ net1026 VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__inv_2
XFILLER_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12264__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08536_ genblk1.genblk1.pcpi_mul.next_rs2\[9\] net1095 _03918_ _03920_ VGND VGND
+ VPWR VPWR _03922_ sky130_fd_sc_hd__and4_1
XFILLER_168_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12395__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A _02083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08467_ net285 net2493 net531 VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__mux2_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1074_X net1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout809_A net812 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07418_ _02951_ _02952_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__nand2_1
X_08398_ _03808_ _03809_ net767 VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07349_ genblk1.genblk1.pcpi_mul.pcpi_rd\[13\] genblk2.pcpi_div.pcpi_rd\[13\] net1110
+ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__mux2_1
XANTENNA__11224__D1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10209__A decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_X net1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ net833 _05061_ _05063_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__a211o_1
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12319__A1 decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11739__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_X net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09019_ net299 net2078 net518 VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__mux2_1
X_10291_ decoded_imm\[19\] net1012 VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__nand2_1
X_12030_ net722 _06484_ net1019 VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09209__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold170 cpuregs\[12\]\[1\] VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 net165 VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_151_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold192 cpuregs\[12\]\[23\] VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__A1 net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07746__B2 decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout650 net654 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout661 net663 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkbuf_4
Xfanout672 net679 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_2
X_13981_ clknet_leaf_199_clk _00435_ VGND VGND VPWR VPWR cpuregs\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout683 net696 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__buf_2
Xfanout694 net695 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__buf_2
XANTENNA__13255__A net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12932_ net1066 reg_sh\[1\] reg_sh\[0\] decoded_imm_j\[1\] _02701_ VGND VGND VPWR
+ VPWR _02121_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_166_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15651_ clknet_leaf_70_clk _01987_ VGND VGND VPWR VPWR cpuregs\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12863_ net1 net2699 _02450_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__mux2_1
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14602_ clknet_leaf_156_clk _00988_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dfxtp_1
X_11814_ _06280_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12255__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15582_ clknet_leaf_35_clk _01918_ VGND VGND VPWR VPWR cpuregs\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12794_ genblk1.genblk1.pcpi_mul.mul_counter\[5\] _06670_ VGND VGND VPWR VPWR _02115_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10805__A1 net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14533_ clknet_leaf_82_clk _00922_ VGND VGND VPWR VPWR decoded_imm\[0\] sky130_fd_sc_hd__dfxtp_2
X_11745_ net1447 net98 net727 VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__mux2_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07399__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12007__B1 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14464_ clknet_leaf_64_clk _00853_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dfxtp_1
X_11676_ net2658 net747 _06230_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__o21a_1
XFILLER_30_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12558__A1 net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13415_ net992 net760 VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__or2_1
XANTENNA__11222__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10627_ cpuregs\[6\]\[8\] cpuregs\[7\]\[8\] net677 VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14395_ clknet_leaf_84_clk _00816_ VGND VGND VPWR VPWR latched_is_lb sky130_fd_sc_hd__dfxtp_1
XANTENNA__08226__A2 net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13346_ net959 _02258_ _02259_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__and3_1
XANTENNA__07904__A_N net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10558_ cpuregs\[14\]\[6\] cpuregs\[15\]\[6\] net673 VGND VGND VPWR VPWR _05252_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11649__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11565__A_N mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13277_ _02194_ _02195_ _02199_ net395 net1032 VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__o32a_1
X_10489_ cpuregs\[28\]\[1\] cpuregs\[29\]\[1\] net683 VGND VGND VPWR VPWR _05188_
+ sky130_fd_sc_hd__mux2_1
X_15016_ clknet_leaf_106_clk net2957 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09119__S net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12228_ net750 _06606_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__nor2_1
XANTENNA__08023__S net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12730__B2 net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ genblk2.pcpi_div.quotient_msk\[18\] net377 net365 net2839 VGND VGND VPWR
+ VPWR _01060_ sky130_fd_sc_hd__a22o_1
XANTENNA__10741__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08958__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06960__A2 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11297__B2 net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12246__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09370_ net2092 net540 net400 VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__mux2_1
X_08321_ net768 _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__and2b_2
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13104__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08252_ reg_out\[3\] reg_next_pc\[3\] net922 VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07203_ net4 net21 net1048 VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__mux2_1
XFILLER_165_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08183_ _03266_ net929 net966 VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__a21o_1
XANTENNA__08217__A2 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12943__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13210__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07134_ net1050 net1054 VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__and2_1
XANTENNA__09818__A decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08281__X net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07065_ net1117 _02628_ genblk2.pcpi_div.quotient\[21\] VGND VGND VPWR VPWR _02630_
+ sky130_fd_sc_hd__a21oi_1
Xoutput220 net1003 VGND VGND VPWR VPWR pcpi_rs1[25] sky130_fd_sc_hd__buf_2
XFILLER_161_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10980__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput231 net231 VGND VGND VPWR VPWR pcpi_rs1[6] sky130_fd_sc_hd__buf_2
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput242 net242 VGND VGND VPWR VPWR pcpi_rs2[16] sky130_fd_sc_hd__buf_2
XANTENNA__09029__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput253 net253 VGND VGND VPWR VPWR pcpi_rs2[26] sky130_fd_sc_hd__buf_2
Xoutput264 net264 VGND VGND VPWR VPWR pcpi_rs2[7] sky130_fd_sc_hd__buf_2
XFILLER_160_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout494_A _04286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1201_A net1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout661_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07967_ _03424_ _03481_ net989 VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__mux2_1
XFILLER_28_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout759_A _04884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11294__S net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09706_ _04499_ _04501_ net2593 net876 VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a2bb2o_1
X_06918_ net1237 net3031 VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__and2_1
XFILLER_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07898_ _03364_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__nand2_1
X_09637_ reg_pc\[24\] net881 _04445_ net851 VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__a22o_1
X_06849_ net1232 _02451_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout926_A net927 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10211__B net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1191_X net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12237__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09568_ count_instr\[56\] count_instr\[55\] count_instr\[54\] _04403_ VGND VGND VPWR
+ VPWR _04408_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_65_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08456__X _03857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07801__A net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08519_ net892 _03905_ _03907_ net2773 net1201 VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__a32o_1
X_09499_ net2805 _04362_ net1239 VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__o21ai_1
XFILLER_169_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13014__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11530_ mem_rdata_q\[23\] net2053 net737 VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__mux2_1
XANTENNA__07664__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11461_ cpuregs\[19\]\[30\] net636 net598 VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__o21a_1
XANTENNA__09405__A1 net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12853__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13200_ net1051 decoded_imm\[0\] _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__o21a_1
X_10412_ net254 _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__or2_1
XANTENNA__11212__A1 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14180_ clknet_leaf_109_clk _00634_ VGND VGND VPWR VPWR count_instr\[51\] sky130_fd_sc_hd__dfxtp_1
X_11392_ cpuregs\[16\]\[28\] net688 VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__or2_1
XFILLER_136_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13131_ latched_rd\[4\] latched_rd\[3\] latched_rd\[2\] VGND VGND VPWR VPWR _02127_
+ sky130_fd_sc_hd__nand3b_1
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10343_ cpuregs\[14\]\[31\] cpuregs\[15\]\[31\] net695 VGND VGND VPWR VPWR _05049_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13062_ net2498 net85 net534 VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__mux2_1
X_10274_ _04933_ _04979_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__or2_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12013_ net721 _06470_ net1024 VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11993__A net1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12712__B2 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07195__A2 net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout480 net483 VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout491 _04287_ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_4
XANTENNA__11279__A1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13964_ clknet_leaf_51_clk _00418_ VGND VGND VPWR VPWR cpuregs\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10402__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input10_X net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12915_ net326 net2278 net457 VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__mux2_1
XANTENNA__10487__C1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output211_A net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13895_ clknet_leaf_60_clk _00349_ VGND VGND VPWR VPWR cpuregs\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15634_ clknet_leaf_198_clk _01970_ VGND VGND VPWR VPWR cpuregs\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12846_ net339 net2176 net459 VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__mux2_1
XFILLER_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15565_ clknet_leaf_20_clk _01901_ VGND VGND VPWR VPWR cpuregs\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12777_ net1220 genblk1.genblk1.pcpi_mul.next_rs1\[45\] net2517 net909 net765 VGND
+ VGND VPWR VPWR _01416_ sky130_fd_sc_hd__a221o_1
XANTENNA__11233__A net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14516_ clknet_leaf_77_clk _00905_ VGND VGND VPWR VPWR decoded_imm_j\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _02363_ net1089 net1232 VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_155_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15496_ clknet_leaf_131_clk _01832_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dfxtp_1
X_14447_ clknet_leaf_98_clk _00836_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11659_ decoded_imm_j\[17\] net9 net546 VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__mux2_1
XANTENNA__12400__A0 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09947__A2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14378_ clknet_leaf_131_clk _00799_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dfxtp_2
XANTENNA__07958__A1 net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold906 cpuregs\[9\]\[4\] VGND VGND VPWR VPWR net2220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold917 cpuregs\[3\]\[12\] VGND VGND VPWR VPWR net2231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__B2 net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold928 cpuregs\[6\]\[7\] VGND VGND VPWR VPWR net2242 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ net960 _04991_ _02244_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__nor3_1
Xhold939 cpuregs\[7\]\[30\] VGND VGND VPWR VPWR net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07158__A reg_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12703__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12703__B2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08870_ genblk1.genblk1.pcpi_mul.rd\[60\] genblk1.genblk1.pcpi_mul.rdx\[60\] VGND
+ VGND VPWR VPWR _04204_ sky130_fd_sc_hd__nand2_1
XFILLER_85_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1606 genblk2.pcpi_div.quotient_msk\[8\] VGND VGND VPWR VPWR net2920 sky130_fd_sc_hd__dlygate4sd3_1
X_07821_ _03337_ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nor2_1
Xhold1617 genblk1.genblk1.pcpi_mul.rd\[35\] VGND VGND VPWR VPWR net2931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 genblk1.genblk1.pcpi_mul.next_rs2\[41\] VGND VGND VPWR VPWR net2942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1639 genblk1.genblk1.pcpi_mul.next_rs2\[36\] VGND VGND VPWR VPWR net2953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12003__S net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07752_ net252 net1002 VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__nand2_1
X_07683_ net798 _03202_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__or2_1
XANTENNA__12938__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09422_ count_instr\[3\] count_instr\[2\] _04303_ _04312_ VGND VGND VPWR VPWR _04313_
+ sky130_fd_sc_hd__and4_1
XANTENNA__11690__A1 net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09312__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09353_ net1675 net314 net477 VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__mux2_1
XANTENNA__09635__B2 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08304_ reg_out\[29\] reg_next_pc\[29\] net924 VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09284_ net1500 net316 net486 VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__mux2_1
X_08235_ net1177 net244 net940 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__mux2_1
XFILLER_165_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1151_A net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A _04279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13195__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09938__A2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08166_ _03657_ _03658_ _03653_ VGND VGND VPWR VPWR alu_out\[25\] sky130_fd_sc_hd__o21ai_1
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07117_ net1123 genblk2.pcpi_div.quotient\[29\] _02671_ _02673_ net952 VGND VGND
+ VPWR VPWR _02674_ sky130_fd_sc_hd__a311o_1
XANTENNA__08071__B1 net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08097_ _03339_ _03595_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__o21a_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout1037_X net1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07048_ genblk2.pcpi_div.dividend\[18\] net1114 _02614_ net947 VGND VGND VPWR VPWR
+ _02616_ sky130_fd_sc_hd__a31o_1
Xclkload90 clknet_leaf_141_clk VGND VGND VPWR VPWR clkload90/Y sky130_fd_sc_hd__clkinv_2
XFILLER_115_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout876_A net882 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12702__A _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1204_X net1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_X net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12170__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout664_X net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08999_ net537 net1964 net516 VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__mux2_1
XFILLER_88_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13009__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10222__A decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10961_ cpuregs\[1\]\[17\] net621 net605 _05643_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout831_X net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12848__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07334__C1 _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11130__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11752__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12700_ _02384_ net912 VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__nor2_1
X_13680_ clknet_leaf_144_clk _00134_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_10892_ cpuregs\[8\]\[15\] net648 VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__or2_1
XANTENNA__09222__S net495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12631_ _02394_ net911 VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15350_ clknet_leaf_42_clk _01690_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_1
X_12562_ genblk2.pcpi_div.divisor\[60\] net874 _02042_ _02043_ VGND VGND VPWR VPWR
+ _02044_ sky130_fd_sc_hd__o22a_1
X_14301_ clknet_leaf_126_clk _00755_ VGND VGND VPWR VPWR count_cycle\[46\] sky130_fd_sc_hd__dfxtp_1
X_11513_ net2737 mem_rdata_q\[6\] net746 VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__mux2_1
XFILLER_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ clknet_leaf_199_clk _01622_ VGND VGND VPWR VPWR cpuregs\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12583__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _05105_ net718 net1163 VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14232_ clknet_leaf_173_clk _00686_ VGND VGND VPWR VPWR reg_next_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_11444_ cpuregs\[3\]\[30\] net636 net598 _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__o211a_1
XFILLER_137_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11199__S net821 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08062__B1 net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14163_ clknet_leaf_126_clk net2583 VGND VGND VPWR VPWR count_instr\[34\] sky130_fd_sc_hd__dfxtp_1
X_11375_ cpuregs\[8\]\[28\] net689 VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13114_ net341 net2270 net435 VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__mux2_1
X_10326_ _04895_ _05031_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__nor2_1
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14094_ clknet_leaf_39_clk _00548_ VGND VGND VPWR VPWR cpuregs\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output259_A net259 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ net1477 net68 net534 VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__mux2_1
XFILLER_79_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10257_ _04943_ _04962_ _04941_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__o21ai_1
Xfanout1220 net1221 VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__buf_2
XFILLER_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07168__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12161__A2 net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07706__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1231 net1241 VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__buf_2
X_10188_ decoded_imm\[29\] net994 VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__nor2_1
XANTENNA__08301__S net983 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14996_ clknet_leaf_148_clk _01348_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13947_ clknet_leaf_197_clk _00401_ VGND VGND VPWR VPWR cpuregs\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11662__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_185_clk _00332_ VGND VGND VPWR VPWR cpuregs\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09132__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15617_ clknet_leaf_48_clk _01953_ VGND VGND VPWR VPWR cpuregs\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12829_ net279 net2119 net466 VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__mux2_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11424__A1 net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15548_ clknet_leaf_43_clk _01884_ VGND VGND VPWR VPWR cpuregs\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12621__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08971__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_150_clk sky130_fd_sc_hd__clkbuf_8
X_15479_ clknet_leaf_10_clk _01815_ VGND VGND VPWR VPWR cpuregs\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13177__A1 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08020_ _03350_ _03352_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__nand2_1
Xhold703 cpuregs\[25\]\[23\] VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 cpuregs\[3\]\[20\] VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 cpuregs\[4\]\[27\] VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10935__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold736 cpuregs\[2\]\[3\] VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 cpuregs\[31\]\[31\] VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 cpuregs\[16\]\[24\] VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _04742_ _04743_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__nor2_1
Xhold769 cpuregs\[6\]\[8\] VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ _04200_ _04202_ _04199_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12522__A net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12152__A2 net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09307__S net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08853_ genblk1.genblk1.pcpi_mul.rd\[57\] genblk1.genblk1.pcpi_mul.next_rs2\[58\]
+ net1105 VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nand3_1
Xhold1403 genblk2.pcpi_div.divisor\[4\] VGND VGND VPWR VPWR net2717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 genblk2.pcpi_div.divisor\[14\] VGND VGND VPWR VPWR net2728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 genblk1.genblk1.pcpi_mul.pcpi_rd\[11\] VGND VGND VPWR VPWR net2739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14510__Q decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1436 genblk2.pcpi_div.quotient_msk\[2\] VGND VGND VPWR VPWR net2750 sky130_fd_sc_hd__dlygate4sd3_1
X_07804_ net1158 net1008 VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__or2_1
Xhold1447 genblk2.pcpi_div.quotient\[20\] VGND VGND VPWR VPWR net2761 sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ _04131_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__inv_2
Xhold1458 genblk1.genblk1.pcpi_mul.next_rs1\[0\] VGND VGND VPWR VPWR net2772 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1469 count_cycle\[50\] VGND VGND VPWR VPWR net2783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07735_ net835 _03249_ _03251_ _03253_ net794 VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07316__C1 _02853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1199_A net1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11663__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07666_ cpuregs\[27\]\[2\] net641 net601 _03186_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__o211a_1
XFILLER_52_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10696__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09042__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09405_ net1089 net1186 count_instr\[0\] VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a21o_1
XFILLER_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07597_ count_instr\[62\] net1133 net1141 count_cycle\[62\] VGND VGND VPWR VPWR _03120_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout624_A net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1310 VGND VGND VPWR VPWR picorv32_1310/HI trace_data[32] sky130_fd_sc_hd__conb_1
X_09336_ net1394 net542 net476 VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__mux2_1
XANTENNA__13499__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout412_X net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09267_ net1517 net574 net487 VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_141_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_141_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1154_X net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11601__A net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08218_ net1180 net1059 net1168 net942 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__a22o_1
X_09198_ net2199 net585 net494 VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11179__B1 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11320__B net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08149_ _03323_ _03327_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__and2_1
XFILLER_136_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11160_ net783 _05828_ _05837_ net778 VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__o211a_1
XANTENNA__07252__D1 net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout781_X net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout879_X net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11747__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10111_ count_cycle\[41\] _04836_ count_cycle\[42\] VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__a21o_1
XFILLER_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11091_ net798 _05768_ _05770_ net838 VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a211o_1
XFILLER_122_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12432__A net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ count_cycle\[16\] count_cycle\[17\] VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__and2_1
XANTENNA__09217__S net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12143__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold30 cpuregs\[30\]\[12\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold41 _01377_ VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11048__A net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14850_ clknet_leaf_56_clk _01202_ VGND VGND VPWR VPWR cpuregs\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07245__B decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold52 net59 VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold63 cpuregs\[26\]\[4\] VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 cpuregs\[26\]\[17\] VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold85 cpuregs\[14\]\[2\] VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 cpuregs\[24\]\[25\] VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_48_clk _00255_ VGND VGND VPWR VPWR cpuregs\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_input18_A mem_rdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14781_ clknet_leaf_155_clk _00036_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12578__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11993_ net1030 _06453_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11103__B1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13263__A net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13732_ clknet_leaf_112_clk _00186_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11654__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10944_ cpuregs\[30\]\[16\] cpuregs\[31\]\[16\] net656 VGND VGND VPWR VPWR _05628_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10457__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07322__A2 decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13663_ clknet_leaf_120_clk _00117_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10875_ net828 _05556_ _05558_ _05560_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__a211o_1
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15402_ clknet_leaf_179_clk _01741_ VGND VGND VPWR VPWR cpuregs\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12614_ net1200 net2902 net893 net2914 _02056_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__a221o_1
XFILLER_169_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11406__B2 net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13594_ net1322 VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_152_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15333_ clknet_leaf_159_clk _01673_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_1
XANTENNA__08283__A0 net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12545_ genblk2.pcpi_div.divisor\[56\] net874 _02029_ _02030_ VGND VGND VPWR VPWR
+ _02031_ sky130_fd_sc_hd__o22a_1
XFILLER_157_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_132_clk sky130_fd_sc_hd__clkbuf_8
X_15264_ clknet_leaf_52_clk _01605_ VGND VGND VPWR VPWR cpuregs\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12476_ net2599 net386 _06701_ _06702_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_113_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14215_ clknet_leaf_75_clk _00669_ VGND VGND VPWR VPWR reg_pc\[23\] sky130_fd_sc_hd__dfxtp_2
X_11427_ _06096_ _06097_ net808 VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08035__B1 net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15195_ clknet_leaf_19_clk _01544_ VGND VGND VPWR VPWR cpuregs\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14146_ clknet_leaf_110_clk net2562 VGND VGND VPWR VPWR count_instr\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output86_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11358_ cpuregs\[19\]\[27\] net638 net599 VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__o21a_1
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12119__C1 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11657__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10309_ _04906_ _04907_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__or2_1
XFILLER_141_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14077_ clknet_leaf_198_clk _00531_ VGND VGND VPWR VPWR cpuregs\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07707__Y _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11289_ _05945_ _05946_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__a21oi_2
X_13028_ net304 net2330 net446 VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_199_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_199_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11342__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1050 net214 VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1062 VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__clkbuf_2
Xfanout1072 net1073 VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__buf_2
XFILLER_120_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1083 net1084 VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08966__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1094 net1109 VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__buf_2
XFILLER_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14979_ clknet_leaf_112_clk _01331_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_07520_ _03046_ _03047_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11645__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07451_ _02977_ _02982_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15161__Q mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07602__C _03124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14419__D alu_out\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07382_ net1063 net1020 _02919_ net1078 _02915_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__a221o_1
X_09121_ net1959 net294 net506 VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12517__A net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13112__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09052_ net301 net2167 net514 VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__mux2_1
X_08003_ _03352_ net934 VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__nor2_1
XANTENNA__14505__Q instr_rdinstrh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12951__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold500 cpuregs\[10\]\[23\] VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 cpuregs\[31\]\[4\] VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 genblk1.genblk1.pcpi_mul.next_rs1\[30\] VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold533 cpuregs\[28\]\[7\] VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 cpuregs\[27\]\[8\] VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 cpuregs\[23\]\[17\] VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 cpuregs\[23\]\[11\] VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold577 cpuregs\[4\]\[19\] VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 cpuregs\[10\]\[25\] VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13348__A net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09954_ _04448_ _04719_ net985 VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__o21a_1
XFILLER_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold599 cpuregs\[5\]\[18\] VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09037__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08905_ net1210 net2706 net899 _04229_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__a22o_1
X_09885_ _04629_ _04640_ _04641_ _04654_ _04652_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__a41o_1
Xhold1200 cpuregs\[1\]\[30\] VGND VGND VPWR VPWR net2514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A _03761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1211 cpuregs\[3\]\[31\] VGND VGND VPWR VPWR net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1222 genblk2.pcpi_div.divisor\[44\] VGND VGND VPWR VPWR net2536 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ _04175_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__inv_2
Xhold1233 cpuregs\[30\]\[26\] VGND VGND VPWR VPWR net2547 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1244 count_instr\[1\] VGND VGND VPWR VPWR net2558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1255 reg_next_pc\[16\] VGND VGND VPWR VPWR net2569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07552__A2 net1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1266 _01106_ VGND VGND VPWR VPWR net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1277 _00636_ VGND VGND VPWR VPWR net2591 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__inv_2
XFILLER_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12398__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1288 genblk2.pcpi_div.quotient_msk\[0\] VGND VGND VPWR VPWR net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _00825_ VGND VGND VPWR VPWR net2613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout839_A _03136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07718_ _03234_ _03236_ net785 VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__a21o_1
XANTENNA__10439__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08698_ _04056_ _04058_ _04051_ _04054_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_24_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07649_ net986 decoded_imm_j\[4\] _03168_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__o21a_2
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10660_ net1076 decoded_imm\[8\] VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__or2_1
XFILLER_167_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08265__A0 net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09319_ net1401 net319 net479 VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10591_ cpuregs\[0\]\[7\] net673 VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_114_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_167_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12427__A net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13022__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12330_ net1148 decoded_imm_j\[9\] net744 VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__and3_1
XFILLER_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08116__S net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout996_X net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12261_ net2692 net381 net369 net2775 VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__a22o_1
XANTENNA__12861__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14000_ clknet_leaf_29_clk _00454_ VGND VGND VPWR VPWR cpuregs\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11212_ net785 _05879_ _05888_ net776 VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__o211a_1
XFILLER_123_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12192_ net749 _06588_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__nor2_1
XANTENNA__10375__A1 net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput42 net42 VGND VGND VPWR VPWR mem_addr[17] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VGND VGND VPWR VPWR mem_addr[28] sky130_fd_sc_hd__buf_2
X_11143_ net1082 _05820_ net856 VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__a21oi_1
Xoutput64 net64 VGND VGND VPWR VPWR mem_addr[9] sky130_fd_sc_hd__buf_2
XFILLER_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput75 net75 VGND VGND VPWR VPWR mem_la_addr[19] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VGND VGND VPWR VPWR mem_la_addr[2] sky130_fd_sc_hd__buf_2
Xoutput97 net1180 VGND VGND VPWR VPWR mem_la_wdata[0] sky130_fd_sc_hd__buf_2
X_11074_ cpuregs\[24\]\[20\] net658 VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__or2_1
XFILLER_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14902_ clknet_leaf_143_clk _01254_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_10025_ count_cycle\[10\] _04781_ count_cycle\[11\] VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__a21o_1
XFILLER_37_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07543__X _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14833_ clknet_leaf_187_clk _01185_ VGND VGND VPWR VPWR cpuregs\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output124_A net1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11506__A _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14764_ clknet_leaf_170_clk _00018_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ net1039 _06434_ net726 VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__o21a_1
XANTENNA__10410__A net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13715_ clknet_leaf_144_clk _00169_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10927_ cpuregs\[12\]\[16\] cpuregs\[13\]\[16\] net655 VGND VGND VPWR VPWR _05611_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14695_ clknet_leaf_138_clk _01080_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13646_ clknet_leaf_146_clk _00100_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10858_ cpuregs\[11\]\[14\] net620 net590 _05543_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__o211a_1
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_105_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_8
X_13577_ net310 net2230 net413 VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__mux2_1
X_10789_ _05475_ _05476_ net809 VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__mux2_1
XFILLER_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15316_ clknet_leaf_8_clk _01656_ VGND VGND VPWR VPWR cpuregs\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12528_ net247 _02017_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__xor2_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15247_ clknet_leaf_40_clk _01588_ VGND VGND VPWR VPWR cpuregs\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12459_ _06689_ net2551 net383 VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__mux2_1
XFILLER_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15178_ clknet_leaf_89_clk _01527_ VGND VGND VPWR VPWR mem_rdata_q\[29\] sky130_fd_sc_hd__dfxtp_2
XFILLER_141_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14129_ clknet_leaf_83_clk _00583_ VGND VGND VPWR VPWR count_instr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout309 net311 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_1
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06951_ genblk2.pcpi_div.dividend\[5\] _02531_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15156__Q mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11315__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09670_ _04467_ _04468_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__and2_1
X_06882_ net1182 net1149 VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08621_ _03985_ _03988_ _03990_ _03992_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13107__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08552_ genblk1.genblk1.pcpi_mul.rd\[11\] genblk1.genblk1.pcpi_mul.next_rs2\[12\]
+ net1091 VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nand3_1
XFILLER_51_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07503_ _03007_ _03019_ _03031_ _03009_ _03020_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__o221a_1
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12291__A1 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12946__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08483_ net1199 net2759 net916 net1181 VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07434_ net11 net939 net936 VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09320__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12043__A1 net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07365_ _02898_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_4_8_0_clk_X clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_A _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_A net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10054__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09104_ net1568 net405 net505 VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__mux2_1
X_07296_ net19 _02689_ _02694_ net2 _02812_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__o221a_1
X_09035_ net521 net2143 net513 VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1231_A net1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold330 net149 VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 cpuregs\[28\]\[18\] VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 cpuregs\[20\]\[24\] VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net696 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_A net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold363 cpuregs\[14\]\[1\] VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 genblk1.genblk1.pcpi_mul.next_rs1\[5\] VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold385 cpuregs\[8\]\[2\] VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 cpuregs\[14\]\[7\] VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout810 net812 VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__buf_4
XFILLER_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout821 _03142_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__buf_2
X_09937_ net1185 _04446_ _04713_ net849 VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_70_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout832 net833 VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__clkbuf_4
Xfanout843 net844 VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__buf_2
XFILLER_132_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11306__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout854 net855 VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__clkbuf_2
Xfanout865 net866 VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout876 net882 VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__clkbuf_4
Xfanout887 net891 VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__clkbuf_2
X_09868_ net2578 net877 _04650_ net847 VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__a22o_1
Xfanout898 _03879_ VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__clkbuf_2
Xhold1030 cpuregs\[9\]\[2\] VGND VGND VPWR VPWR net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 cpuregs\[23\]\[28\] VGND VGND VPWR VPWR net2355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1052 cpuregs\[18\]\[8\] VGND VGND VPWR VPWR net2366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07804__A net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08819_ _04160_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__inv_2
Xhold1063 cpuregs\[9\]\[24\] VGND VGND VPWR VPWR net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 cpuregs\[18\]\[14\] VGND VGND VPWR VPWR net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09799_ _04435_ _04577_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__xnor2_1
Xhold1085 cpuregs\[11\]\[29\] VGND VGND VPWR VPWR net2399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13017__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ genblk2.pcpi_div.divisor\[11\] genblk2.pcpi_div.dividend\[11\] VGND VGND
+ VPWR VPWR _06301_ sky130_fd_sc_hd__nand2b_1
Xhold1096 _01371_ VGND VGND VPWR VPWR net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10230__A decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10817__C1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11761_ net1807 net115 net729 VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout911_X net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12282__A1 net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12856__S net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12282__B2 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11760__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13500_ net1975 net352 net419 VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__mux2_1
X_10712_ cpuregs\[11\]\[10\] net625 net593 _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__o211a_1
XFILLER_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14480_ clknet_leaf_96_clk _00869_ VGND VGND VPWR VPWR instr_sb sky130_fd_sc_hd__dfxtp_1
XANTENNA__11490__C1 net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11692_ net1858 net522 net373 VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__mux2_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09230__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13431_ _04896_ _05030_ _02334_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08238__A0 net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10643_ cpuregs\[30\]\[8\] cpuregs\[31\]\[8\] net670 VGND VGND VPWR VPWR _05335_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12034__A1 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13362_ _05003_ _05005_ _05007_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__o21ai_1
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10574_ net830 _05263_ _05265_ _05267_ net790 VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15101_ clknet_leaf_38_clk _01453_ VGND VGND VPWR VPWR cpuregs\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ decoded_imm\[17\] net743 _06632_ _06635_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__o22a_1
XANTENNA__12591__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13293_ _02208_ _02209_ _02213_ net395 net205 VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__o32a_1
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07538__X _03065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15032_ clknet_leaf_136_clk net1332 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09738__B1 _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12337__A2 net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12244_ net2715 net382 net366 genblk2.pcpi_div.divisor\[8\] VGND VGND VPWR VPWR _01113_
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ genblk2.pcpi_div.quotient_msk\[1\] net277 net2999 VGND VGND VPWR VPWR _06580_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__10405__A net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11126_ _05803_ _05804_ net810 VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__mux2_1
XFILLER_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output241_A net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ net831 _05733_ _05735_ _05737_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_108_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ net3039 _04771_ _04773_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_160_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13435__B _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14816_ clknet_leaf_79_clk _01168_ VGND VGND VPWR VPWR decoded_imm\[6\] sky130_fd_sc_hd__dfxtp_2
X_14747_ clknet_leaf_158_clk net2744 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11959_ _06312_ _06313_ _06314_ _06325_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__a211o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14678_ clknet_leaf_162_clk _01063_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09140__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08229__B1 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12025__A1 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13629_ clknet_leaf_120_clk _00083_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09977__B1 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07150_ net1073 net1084 net1068 net1061 VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__or4_1
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10587__A1 net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11784__B1 _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07081_ genblk2.pcpi_div.quotient\[21\] genblk2.pcpi_div.quotient\[22\] _02628_ VGND
+ VGND VPWR VPWR _02644_ sky130_fd_sc_hd__or3_1
XANTENNA__07452__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11536__A0 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07983_ net1143 _03426_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__a21o_1
X_09722_ _04427_ _04428_ _04429_ _04488_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__nand4_2
XFILLER_68_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06934_ genblk2.pcpi_div.dividend\[1\] genblk2.pcpi_div.dividend\[0\] net1126 VGND
+ VGND VPWR VPWR _02518_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08279__X net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09315__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09901__B1 net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09653_ _04422_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__nand2_1
XFILLER_95_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06865_ _02370_ net1208 VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__nor2_1
XFILLER_55_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10511__A1 net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08604_ genblk1.genblk1.pcpi_mul.rd\[19\] genblk1.genblk1.pcpi_mul.next_rs2\[20\]
+ net1099 VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__nand3_1
XFILLER_82_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09584_ count_instr\[62\] count_instr\[61\] count_instr\[60\] _04413_ VGND VGND VPWR
+ VPWR _04418_ sky130_fd_sc_hd__and4_1
X_06796_ net1028 VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__inv_2
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08535_ genblk1.genblk1.pcpi_mul.next_rs2\[9\] net1094 _03918_ _03920_ VGND VGND
+ VPWR VPWR _03921_ sky130_fd_sc_hd__a22o_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08466_ _03861_ _03864_ net769 VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__mux2_1
XFILLER_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09050__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ reg_pc\[18\] decoded_imm\[18\] VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__or2_1
XANTENNA__13213__B1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08397_ reg_pc\[16\] _03805_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__xor2_1
XFILLER_149_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout1067_X net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07348_ count_cycle\[13\] net971 net841 _02887_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o211a_1
XFILLER_109_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07279_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1234_X net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09018_ net304 net2195 net519 VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__mux2_1
XANTENNA__11527__A0 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10290_ _04915_ _04992_ _04914_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__a21o_1
XFILLER_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold160 cpuregs\[31\]\[2\] VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__A decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold171 cpuregs\[15\]\[4\] VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 genblk1.genblk1.pcpi_mul.pcpi_rd\[30\] VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold193 cpuregs\[20\]\[7\] VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout861_X net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10750__A1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_X net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout640 net641 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 net654 VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__buf_2
XANTENNA__11755__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout662 net663 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__dlymetal6s2s_1
X_13980_ clknet_leaf_197_clk _00434_ VGND VGND VPWR VPWR cpuregs\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xfanout673 net676 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__buf_2
XFILLER_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12440__A net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout684 net687 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_2
XANTENNA__09225__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout695 net696 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__buf_2
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12931_ net3016 _02502_ _05169_ _02120_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__o22a_1
XFILLER_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10502__B2 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12862_ net278 net2466 net461 VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__mux2_1
X_15650_ clknet_leaf_46_clk _01986_ VGND VGND VPWR VPWR cpuregs\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ genblk2.pcpi_div.dividend\[18\] genblk2.pcpi_div.divisor\[18\] VGND VGND
+ VPWR VPWR _06284_ sky130_fd_sc_hd__nand2b_1
X_14601_ clknet_leaf_145_clk _00987_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dfxtp_1
XFILLER_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15581_ clknet_leaf_17_clk _01917_ VGND VGND VPWR VPWR cpuregs\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12793_ net1215 net1961 net1582 net906 net762 VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ clknet_leaf_81_clk _00921_ VGND VGND VPWR VPWR decoded_imm_j\[3\] sky130_fd_sc_hd__dfxtp_2
X_11744_ net1635 net128 net730 VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__mux2_1
XFILLER_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10805__A2 _05491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07667__D1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14463_ clknet_leaf_64_clk _00852_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dfxtp_1
XANTENNA__12007__A1 net1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11675_ is_alu_reg_imm _06179_ net737 instr_jalr VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__a211o_1
X_13414_ net569 _05999_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__nor2_1
XFILLER_139_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10626_ net1169 net854 _05317_ _05318_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__a22o_1
XFILLER_168_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14394_ clknet_leaf_85_clk _00815_ VGND VGND VPWR VPWR latched_is_lh sky130_fd_sc_hd__dfxtp_1
XFILLER_155_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13345_ _05000_ _05004_ _04996_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07434__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10557_ _05248_ _05250_ net781 VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__a21o_1
XANTENNA__11230__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11518__A0 mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08304__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13276_ net556 _02175_ _02196_ _02198_ net391 VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__a311o_1
X_10488_ cpuregs\[30\]\[1\] cpuregs\[31\]\[1\] net686 VGND VGND VPWR VPWR _05187_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12334__B decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15015_ clknet_leaf_106_clk net2946 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_12227_ net3072 net275 net2854 VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09924__A net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12158_ net2856 net378 net365 net2893 VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__a22o_1
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__06945__B1 net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11109_ cpuregs\[4\]\[21\] net684 VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__or2_1
XFILLER_111_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12089_ net1006 _06528_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__or2_1
XANTENNA__09135__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11297__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_56_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08974__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13443__B1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08320_ reg_out\[0\] alu_out_q\[0\] net1155 VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__mux2_1
XFILLER_33_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08251_ net1045 _03709_ net981 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_31_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_969 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07202_ net1074 _02749_ _02750_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__and3_1
XANTENNA__11206__C1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08182_ net771 _03671_ _03672_ _03668_ VGND VGND VPWR VPWR alu_out\[27\] sky130_fd_sc_hd__a31o_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07133_ _02685_ _02687_ net948 VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11221__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13120__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07178__X _02729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07064_ net1124 genblk2.pcpi_div.quotient\[21\] _02628_ VGND VGND VPWR VPWR _02629_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11509__A0 net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput210 net1019 VGND VGND VPWR VPWR pcpi_rs1[16] sky130_fd_sc_hd__buf_2
Xoutput221 net1001 VGND VGND VPWR VPWR pcpi_rs1[26] sky130_fd_sc_hd__buf_2
Xoutput232 net1037 VGND VGND VPWR VPWR pcpi_rs1[7] sky130_fd_sc_hd__buf_2
XANTENNA__14513__Q decoded_imm_j\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput243 net243 VGND VGND VPWR VPWR pcpi_rs2[17] sky130_fd_sc_hd__buf_2
XANTENNA__07338__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput254 net254 VGND VGND VPWR VPWR pcpi_rs2[27] sky130_fd_sc_hd__buf_2
XFILLER_99_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput265 net1168 VGND VGND VPWR VPWR pcpi_rs2[8] sky130_fd_sc_hd__buf_2
XANTENNA__07189__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12721__A2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout487_A _04288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13356__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07966_ _03277_ _03284_ _03474_ _03276_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__a31o_1
XFILLER_102_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09045__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09705_ net1183 _04427_ _04500_ _02489_ net846 VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__o221ai_1
X_06917_ net1061 _02483_ _02494_ _02506_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__a31o_1
XFILLER_28_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07897_ _03360_ _03414_ _03411_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_94_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout275_X net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_A net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09636_ _03840_ reg_next_pc\[24\] net926 VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__mux2_2
X_06848_ _02419_ _02447_ net965 _02448_ mem_do_rinst VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__a32o_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09567_ _04406_ _04407_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__nor2_1
X_06779_ net1061 VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout442_X net442 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13434__B1 _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10919__S net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1184_X net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09102__A1 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08518_ _03906_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__inv_2
XANTENNA__11445__C1 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07801__B net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09498_ count_instr\[31\] count_instr\[30\] count_instr\[29\] _04358_ VGND VGND VPWR
+ VPWR _04363_ sky130_fd_sc_hd__and4_2
XFILLER_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11996__B1 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08449_ reg_pc\[26\] _03847_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout707_X net707 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11460_ cpuregs\[17\]\[30\] net636 net612 _06129_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__o211a_1
XFILLER_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08472__X _03870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09405__A2 net1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10411_ net253 _05115_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__or2_1
XFILLER_125_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11391_ _06061_ _06062_ net817 VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__mux2_1
XFILLER_99_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13030__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13130_ net281 net2378 net438 VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__mux2_1
X_10342_ net833 _05043_ _05047_ net784 VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__a211o_1
XFILLER_125_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13061_ net1556 net84 net533 VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__mux2_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10273_ _04929_ _04930_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__nand2_1
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12012_ net1027 _06464_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__or2_1
XFILLER_151_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13266__A net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout470 _02051_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__buf_2
Xfanout481 _04291_ VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 net493 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_4
X_13963_ clknet_leaf_66_clk _00417_ VGND VGND VPWR VPWR cpuregs\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10402__B net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13553__X _02358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12914_ net331 net2153 net455 VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__mux2_1
X_13894_ clknet_leaf_30_clk _00348_ VGND VGND VPWR VPWR cpuregs\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12845_ net344 net2380 net460 VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__mux2_1
X_15633_ clknet_leaf_191_clk _01969_ VGND VGND VPWR VPWR cpuregs\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output204_A net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12776_ net1220 net2107 net2541 net909 net765 VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__a221o_1
XFILLER_14_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15564_ clknet_leaf_21_clk _01900_ VGND VGND VPWR VPWR cpuregs\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11987__B1 net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07203__S net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11727_ net1208 _02487_ _06149_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__or3_2
X_14515_ clknet_leaf_77_clk _00904_ VGND VGND VPWR VPWR decoded_imm_j\[12\] sky130_fd_sc_hd__dfxtp_1
X_15495_ clknet_leaf_131_clk _01831_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_155_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14446_ clknet_leaf_98_clk _00835_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dfxtp_2
X_11658_ decoded_imm_j\[16\] net8 net546 VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__mux2_1
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10609_ cpuregs\[16\]\[7\] net665 VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__or2_1
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14377_ clknet_leaf_78_clk _00798_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dfxtp_2
XFILLER_155_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11589_ net2864 net562 _06184_ _06192_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__a22o_1
Xhold907 cpuregs\[1\]\[7\] VGND VGND VPWR VPWR net2221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__A2 net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold918 cpuregs\[17\]\[8\] VGND VGND VPWR VPWR net2232 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ _04987_ _04989_ _04990_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_133_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold929 cpuregs\[9\]\[5\] VGND VGND VPWR VPWR net2243 sky130_fd_sc_hd__dlygate4sd3_1
X_13259_ net1038 net753 net556 _02161_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o211a_1
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08969__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12164__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10714__A1 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07820_ net244 net1014 VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__nor2_1
XFILLER_111_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1607 genblk1.genblk1.pcpi_mul.rd\[27\] VGND VGND VPWR VPWR net2921 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12080__A net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1618 instr_sh VGND VGND VPWR VPWR net2932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1629 _01347_ VGND VGND VPWR VPWR net2943 sky130_fd_sc_hd__dlygate4sd3_1
X_07751_ net252 net1002 VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__or2_1
XANTENNA__15164__Q mem_rdata_q\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10478__B1 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07682_ cpuregs\[12\]\[3\] cpuregs\[13\]\[3\] net660 VGND VGND VPWR VPWR _03202_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09421_ count_instr\[5\] count_instr\[4\] VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__and2_1
XFILLER_65_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13115__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09352_ net1438 net319 net476 VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__mux2_1
XANTENNA__09635__A2 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08303_ net996 _03735_ net982 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__mux2_2
XANTENNA__11978__B1 net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_150_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14508__Q decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ net2201 net320 net484 VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__mux2_1
XANTENNA__12954__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08843__B1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08234_ net1178 net1160 net940 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08165_ _03272_ _03656_ _03465_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout402_A _04293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07116_ net1122 genblk2.pcpi_div.quotient\[28\] genblk2.pcpi_div.quotient\[29\] _02670_
+ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__a211oi_1
XANTENNA_clkbuf_leaf_165_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07949__A2 _03457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08096_ _03339_ _03595_ _03465_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__a21oi_1
Xclkload80 clknet_leaf_133_clk VGND VGND VPWR VPWR clkload80/Y sky130_fd_sc_hd__bufinv_16
X_07047_ net1114 _02614_ net3021 VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__a21oi_1
Xclkload91 clknet_leaf_142_clk VGND VGND VPWR VPWR clkload91/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_X net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12702__B net912 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A _05082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08998_ net541 net2067 net517 VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__mux2_1
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ net3052 _03457_ _03461_ _03466_ VGND VGND VPWR VPWR alu_out\[0\] sky130_fd_sc_hd__a211o_1
XANTENNA__12458__B2 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10222__B net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10960_ cpuregs\[0\]\[17\] net656 VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__or2_1
XANTENNA__07371__X _02909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09619_ reg_pc\[15\] net876 _04436_ net846 VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__a22o_1
X_10891_ net796 _05573_ _05575_ net822 VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout824_X net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13407__B1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13025__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12630_ net2993 net885 _02064_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_80_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12561_ _02399_ _05117_ net720 _05083_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__a31o_1
XFILLER_34_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07637__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11512_ net2980 mem_rdata_q\[5\] net746 VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__mux2_1
XFILLER_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14300_ clknet_leaf_126_clk _00754_ VGND VGND VPWR VPWR count_cycle\[45\] sky130_fd_sc_hd__dfxtp_1
X_15280_ clknet_leaf_191_clk _01621_ VGND VGND VPWR VPWR cpuregs\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12492_ net1163 net715 _05105_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_22_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14231_ clknet_leaf_173_clk _00685_ VGND VGND VPWR VPWR reg_next_pc\[8\] sky130_fd_sc_hd__dfxtp_1
X_11443_ cpuregs\[2\]\[30\] net691 VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__or2_1
XFILLER_138_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08062__A1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14162_ clknet_leaf_126_clk _00616_ VGND VGND VPWR VPWR count_instr\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11374_ net817 _06043_ _06045_ net832 VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_78_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13113_ net346 net2126 net436 VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__mux2_1
X_10325_ decoded_imm\[28\] net996 _04896_ _05030_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__a22o_1
X_14093_ clknet_leaf_56_clk _00547_ VGND VGND VPWR VPWR cpuregs\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12146__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09474__A net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13044_ net1347 net67 net534 VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ _04945_ _04947_ _04960_ _04946_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__a31o_1
Xfanout1210 net1222 VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__buf_2
Xfanout1221 net1222 VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_91_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1232 net1233 VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__buf_2
XFILLER_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10187_ _04891_ _04892_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__or2_1
XANTENNA__10413__A net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11228__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_19_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14995_ clknet_leaf_148_clk net2943 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11943__S net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_13946_ clknet_leaf_198_clk _00400_ VGND VGND VPWR VPWR cpuregs\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_13877_ clknet_leaf_188_clk _00331_ VGND VGND VPWR VPWR cpuregs\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15616_ clknet_leaf_34_clk _01952_ VGND VGND VPWR VPWR cpuregs\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12828_ net284 net2128 net466 VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__mux2_1
XFILLER_61_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15547_ clknet_leaf_15_clk _01883_ VGND VGND VPWR VPWR cpuregs\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12759_ net1450 net905 _02113_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__a21o_1
XANTENNA__12621__B2 net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15478_ clknet_leaf_9_clk _01814_ VGND VGND VPWR VPWR cpuregs\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11250__Y _05926_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14429_ clknet_leaf_67_clk alu_out\[29\] VGND VGND VPWR VPWR alu_out_q\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11188__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold704 cpuregs\[25\]\[24\] VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 cpuregs\[27\]\[12\] VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15159__Q mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold726 cpuregs\[27\]\[28\] VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 cpuregs\[2\]\[27\] VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_139_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09970_ net1129 _04450_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__nor2_1
Xhold748 cpuregs\[10\]\[22\] VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 cpuregs\[31\]\[19\] VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09002__A0 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08921_ net1211 net2670 net900 _04237_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a22o_1
XFILLER_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06801__A net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12522__B net716 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08852_ genblk1.genblk1.pcpi_mul.rd\[57\] genblk1.genblk1.pcpi_mul.next_rs2\[58\]
+ net1105 VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__and3_1
Xhold1404 _01109_ VGND VGND VPWR VPWR net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 net191 VGND VGND VPWR VPWR net2729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11360__A1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07803_ net1158 net1007 VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__nor2_1
Xhold1426 reg_next_pc\[4\] VGND VGND VPWR VPWR net2740 sky130_fd_sc_hd__dlygate4sd3_1
X_08783_ _04123_ _04126_ _04128_ _04129_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__o211a_1
Xhold1437 _01043_ VGND VGND VPWR VPWR net2751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1448 _06599_ VGND VGND VPWR VPWR net2762 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12949__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
Xhold1459 genblk1.genblk1.pcpi_mul.rd\[5\] VGND VGND VPWR VPWR net2773 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08108__A2 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07734_ cpuregs\[27\]\[4\] net631 net595 _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__o211a_1
XFILLER_84_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08287__X net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09323__S net482 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07632__A net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07665_ cpuregs\[26\]\[2\] net700 VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__or2_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09404_ net1233 _02439_ _02440_ _04300_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1094_A net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07596_ net359 _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__nor2_1
Xpicorv32_1300 VGND VGND VPWR VPWR picorv32_1300/HI trace_data[22] sky130_fd_sc_hd__conb_1
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_1311 VGND VGND VPWR VPWR picorv32_1311/HI trace_data[33] sky130_fd_sc_hd__conb_1
X_09335_ net1359 net573 net477 VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__mux2_1
XANTENNA__07619__A1 net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11415__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10993__A net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net620 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10623__B1 _05315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09266_ net1651 net577 net485 VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__mux2_1
XFILLER_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08217_ net1181 net1056 net265 net1054 VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a22o_1
X_09197_ net1539 net586 net494 VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__mux2_1
XANTENNA__11179__A1 net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08044__A1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08148_ _03592_ _03608_ _03610_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_95_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_A _02379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07252__C1 net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload180 clknet_leaf_100_clk VGND VGND VPWR VPWR clkload180/X sky130_fd_sc_hd__clkbuf_8
X_08079_ _03346_ net928 net967 VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10110_ net3067 _04836_ _04838_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__o21a_1
XANTENNA__07807__A net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11090_ cpuregs\[5\]\[20\] net624 net811 _05769_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout774_X net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10504__Y _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ count_cycle\[16\] _04791_ net2787 VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_73_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10233__A decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold20 net64 VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 net63 VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 cpuregs\[28\]\[25\] VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 cpuregs\[12\]\[10\] VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 cpuregs\[28\]\[23\] VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12859__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11763__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold75 genblk1.genblk1.pcpi_mul.pcpi_rd\[24\] VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 cpuregs\[24\]\[22\] VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_34_clk _00254_ VGND VGND VPWR VPWR cpuregs\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold97 cpuregs\[26\]\[6\] VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ clknet_leaf_157_clk _00035_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[27\]
+ sky130_fd_sc_hd__dfxtp_2
X_11992_ net1032 _06448_ net723 VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__o21a_1
XANTENNA__11103__A1 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09233__S net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10943_ net824 _05622_ _05624_ _05626_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__a211o_1
X_13731_ clknet_leaf_112_clk _00185_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07261__B decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10874_ cpuregs\[18\]\[14\] net553 _05559_ net780 VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__o22a_1
X_13662_ clknet_leaf_116_clk _00116_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_15401_ clknet_leaf_24_clk _01740_ VGND VGND VPWR VPWR cpuregs\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12613_ genblk1.genblk1.pcpi_mul.mul_waiting net1224 net1172 VGND VGND VPWR VPWR
+ _02056_ sky130_fd_sc_hd__and3_1
X_13593_ net1318 VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12594__S net470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11406__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15332_ clknet_leaf_57_clk _01672_ VGND VGND VPWR VPWR cpuregs\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12544_ _02396_ _05114_ net719 net866 VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__a31o_1
XFILLER_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12475_ net868 _06699_ _06700_ net386 VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__a31oi_1
X_15263_ clknet_leaf_33_clk _01604_ VGND VGND VPWR VPWR cpuregs\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10408__A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11426_ cpuregs\[22\]\[29\] cpuregs\[23\]\[29\] net706 VGND VGND VPWR VPWR _06097_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08035__A1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14214_ clknet_leaf_76_clk _00668_ VGND VGND VPWR VPWR reg_pc\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15194_ clknet_leaf_5_clk _01543_ VGND VGND VPWR VPWR cpuregs\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10917__A1 net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14145_ clknet_leaf_110_clk _00599_ VGND VGND VPWR VPWR count_instr\[16\] sky130_fd_sc_hd__dfxtp_1
X_11357_ cpuregs\[17\]\[27\] net638 net613 _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__o211a_1
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12623__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10308_ _04906_ _04908_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__and2b_1
XANTENNA_output79_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14076_ clknet_leaf_191_clk _00530_ VGND VGND VPWR VPWR cpuregs\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11288_ net775 _05954_ _05962_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__and3_1
XFILLER_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ net305 net2377 net445 VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__mux2_1
X_10239_ decoded_imm\[5\] net1040 VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__nand2_1
Xfanout1040 net1041 VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__clkbuf_4
Xfanout1051 net1052 VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__clkbuf_4
Xfanout1062 cpu_state\[7\] VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__clkbuf_4
Xfanout1073 net1074 VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__clkbuf_4
XFILLER_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1084 net1085 VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1095 net1109 VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlymetal6s2s_1
X_14978_ clknet_leaf_112_clk _01330_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09143__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13929_ clknet_leaf_48_clk _00383_ VGND VGND VPWR VPWR cpuregs\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07450_ _02982_ _02977_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08982__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07381_ genblk1.genblk1.pcpi_mul.pcpi_rd\[15\] genblk2.pcpi_div.pcpi_rd\[15\] net1110
+ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__mux2_1
X_09120_ net2219 net298 net507 VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__mux2_1
XANTENNA__10605__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12517__B net716 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09051_ net306 net2095 net514 VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__mux2_1
XFILLER_129_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12009__S net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08002_ _03511_ _03512_ _03507_ VGND VGND VPWR VPWR alu_out\[7\] sky130_fd_sc_hd__o21ai_1
Xhold501 cpuregs\[10\]\[17\] VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 cpuregs\[30\]\[22\] VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 cpuregs\[25\]\[21\] VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11030__B1 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold534 cpuregs\[3\]\[6\] VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07234__C1 net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold545 cpuregs\[27\]\[9\] VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10752__S net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold556 cpuregs\[16\]\[9\] VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06802__Y _02410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11581__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09318__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold567 cpuregs\[6\]\[4\] VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07627__A net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold578 cpuregs\[22\]\[13\] VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold589 cpuregs\[28\]\[31\] VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _04448_ _04719_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__nand2_1
XANTENNA__13348__B net759 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08904_ _04002_ _04004_ _04001_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__a21bo_1
X_09884_ _04630_ _04640_ _04654_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout1107_A net1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1201 genblk1.genblk1.pcpi_mul.mul_counter\[6\] VGND VGND VPWR VPWR net2515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_4_0_clk_X clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11333__B2 net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1212 cpuregs\[17\]\[0\] VGND VGND VPWR VPWR net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 cpuregs\[18\]\[5\] VGND VGND VPWR VPWR net2537 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ _04167_ _04170_ _04172_ _04173_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__o211a_1
Xhold1234 net151 VGND VGND VPWR VPWR net2548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout567_A net570 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1245 genblk1.genblk1.pcpi_mul.rd\[20\] VGND VGND VPWR VPWR net2559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 genblk2.pcpi_div.divisor\[34\] VGND VGND VPWR VPWR net2570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13364__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08766_ genblk1.genblk1.pcpi_mul.rd\[44\] genblk1.genblk1.pcpi_mul.rdx\[44\] VGND
+ VGND VPWR VPWR _04116_ sky130_fd_sc_hd__nand2_1
Xhold1267 genblk2.pcpi_div.divisor\[54\] VGND VGND VPWR VPWR net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 genblk1.genblk1.pcpi_mul.rd\[8\] VGND VGND VPWR VPWR net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 _01042_ VGND VGND VPWR VPWR net2603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09829__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09053__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07717_ cpuregs\[1\]\[4\] net551 _03235_ net807 net835 VGND VGND VPWR VPWR _03236_
+ sky130_fd_sc_hd__a221o_1
X_08697_ genblk1.genblk1.pcpi_mul.rd\[33\] genblk1.genblk1.pcpi_mul.next_rs2\[34\]
+ net1101 VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout734_A net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07648_ net986 decoded_imm_j\[4\] _03168_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_24_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07579_ _03099_ _03100_ _03101_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout522_X net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09318_ net1390 net321 net479 VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10590_ _05281_ _05282_ net815 VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__mux2_1
XFILLER_167_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09249_ net1440 net324 net490 VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__mux2_1
XFILLER_166_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10228__A decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12260_ genblk2.pcpi_div.divisor\[23\] net381 net369 net2692 VGND VGND VPWR VPWR
+ _01129_ sky130_fd_sc_hd__a22o_1
XANTENNA__08017__A1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11211_ net788 _05883_ _05885_ _05887_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_75_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12191_ net2756 net274 net2877 VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10375__A2 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09228__S net495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput43 net43 VGND VGND VPWR VPWR mem_addr[18] sky130_fd_sc_hd__buf_2
X_11142_ net1080 decoded_imm\[21\] VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__or2_1
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput54 net54 VGND VGND VPWR VPWR mem_addr[29] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VGND VGND VPWR VPWR mem_instr sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR mem_la_addr[20] sky130_fd_sc_hd__buf_2
Xoutput87 net87 VGND VGND VPWR VPWR mem_la_addr[30] sky130_fd_sc_hd__buf_2
XFILLER_150_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11073_ _05751_ _05752_ net810 VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__mux2_1
XFILLER_122_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput98 net98 VGND VGND VPWR VPWR mem_la_wdata[10] sky130_fd_sc_hd__buf_2
XANTENNA__11324__A1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input30_A mem_rdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09752__A decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14901_ clknet_leaf_143_clk _01253_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_10024_ net3054 _04781_ _04783_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__o21a_1
XANTENNA__12589__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14832_ clknet_leaf_184_clk _01184_ VGND VGND VPWR VPWR cpuregs\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14763_ clknet_leaf_152_clk _00017_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _06329_ _06331_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_106_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10410__B net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08087__B net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13714_ clknet_leaf_121_clk _00168_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10926_ cpuregs\[14\]\[16\] cpuregs\[15\]\[16\] net657 VGND VGND VPWR VPWR _05610_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14694_ clknet_leaf_138_clk _01079_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10857_ cpuregs\[10\]\[14\] net653 VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__or2_1
X_13645_ clknet_leaf_147_clk _00099_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12588__A0 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08307__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10788_ cpuregs\[4\]\[12\] cpuregs\[5\]\[12\] net652 VGND VGND VPWR VPWR _05476_
+ sky130_fd_sc_hd__mux2_1
X_13576_ net312 net2407 net413 VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__mux2_1
XANTENNA__10599__C1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15315_ clknet_leaf_4_clk _01655_ VGND VGND VPWR VPWR cpuregs\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11260__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12527_ net245 _05111_ net718 VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_10_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15246_ clknet_leaf_16_clk _01587_ VGND VGND VPWR VPWR cpuregs\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12458_ _06687_ _06688_ genblk2.pcpi_div.divisor\[37\] net865 VGND VGND VPWR VPWR
+ _06689_ sky130_fd_sc_hd__a2bb2o_1
X_11409_ cpuregs\[12\]\[29\] cpuregs\[13\]\[29\] net704 VGND VGND VPWR VPWR _06080_
+ sky130_fd_sc_hd__mux2_1
X_15177_ clknet_leaf_89_clk _01526_ VGND VGND VPWR VPWR mem_rdata_q\[28\] sky130_fd_sc_hd__dfxtp_2
X_12389_ net1418 net280 net363 VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__mux2_1
XFILLER_125_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12760__B1 net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09138__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14128_ clknet_leaf_91_clk _00582_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06950_ genblk2.pcpi_div.dividend\[4\] _02528_ net1125 VGND VGND VPWR VPWR _02531_
+ sky130_fd_sc_hd__o21ai_1
X_14059_ clknet_leaf_66_clk _00513_ VGND VGND VPWR VPWR cpuregs\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08977__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12512__B1 net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09662__A net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06881_ _02380_ net985 VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__nor2_4
XANTENNA__08192__B1 net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ _03990_ _03992_ _03985_ _03988_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__a211o_1
XFILLER_39_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08551_ net887 _03932_ _03934_ net2628 net1197 VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__a32o_1
XFILLER_82_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15172__Q mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07502_ _03008_ _03021_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__or2_1
X_08482_ net1215 net1582 net762 VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__a21o_1
XFILLER_51_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07433_ _02951_ _02956_ _02965_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__a21o_1
XFILLER_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12528__A net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13123__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08247__A1 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07364_ net1064 net1022 _02902_ net1079 _02901_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__a221o_1
XANTENNA__13240__A1 net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09103_ net1773 net407 net505 VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__mux2_1
XANTENNA__14516__Q decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09995__A1 net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07295_ net991 _02836_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__or3_1
XANTENNA__12962__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout315_A _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_A net1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09034_ net527 net2221 net512 VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__mux2_1
XFILLER_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07470__A2 net1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold320 cpuregs\[14\]\[8\] VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 cpuregs\[26\]\[21\] VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold342 cpuregs\[31\]\[15\] VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1224_A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold353 cpuregs\[22\]\[15\] VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09048__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold364 cpuregs\[15\]\[23\] VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 cpuregs\[22\]\[12\] VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold386 net164 VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 net802 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__clkbuf_4
Xfanout811 net812 VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__buf_2
Xhold397 cpuregs\[13\]\[21\] VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout822 net823 VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09936_ _04711_ _04712_ _02489_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_70_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1012_X net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout833 net834 VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__clkbuf_4
Xfanout844 _02702_ VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout855 _05134_ VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__clkbuf_4
Xfanout866 _05083_ VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout851_A net852 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout877 net882 VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout472_X net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09867_ _04440_ _04649_ net1187 VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__mux2_1
Xhold1020 cpuregs\[9\]\[27\] VGND VGND VPWR VPWR net2334 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net890 VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__buf_2
XANTENNA__08183__B1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1031 cpuregs\[19\]\[7\] VGND VGND VPWR VPWR net2345 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A _02509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout899 net900 VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__buf_2
Xhold1042 cpuregs\[5\]\[21\] VGND VGND VPWR VPWR net2356 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13059__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1053 genblk1.genblk1.pcpi_mul.next_rs1\[58\] VGND VGND VPWR VPWR net2367 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07804__B net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08818_ genblk1.genblk1.pcpi_mul.rd\[52\] genblk1.genblk1.pcpi_mul.rdx\[52\] VGND
+ VGND VPWR VPWR _04160_ sky130_fd_sc_hd__nand2_1
Xhold1064 cpuregs\[11\]\[31\] VGND VGND VPWR VPWR net2378 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _04577_ _04435_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__nand2b_1
Xhold1075 cpuregs\[12\]\[28\] VGND VGND VPWR VPWR net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__B1 net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1086 instr_add VGND VGND VPWR VPWR net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 cpuregs\[1\]\[19\] VGND VGND VPWR VPWR net2411 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ genblk1.genblk1.pcpi_mul.rd\[41\] genblk1.genblk1.pcpi_mul.next_rs2\[42\]
+ net1092 VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__nand3_1
XFILLER_27_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10230__B net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11760_ net1669 net114 net729 VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12282__A2 net1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10711_ cpuregs\[10\]\[10\] net666 VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__or2_1
XFILLER_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07820__A net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11691_ net1796 net524 net373 VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__mux2_1
XFILLER_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12438__A net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13033__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13430_ _04896_ _05030_ net958 VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__o21ai_1
X_10642_ net781 _05324_ _05333_ net777 VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__o211a_1
XANTENNA__08238__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _02268_ _02269_ _02273_ net397 net1012 VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__o32a_1
X_10573_ cpuregs\[27\]\[6\] net629 net595 _05266_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__o211a_1
XFILLER_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15100_ clknet_leaf_3_clk _01452_ VGND VGND VPWR VPWR cpuregs\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12312_ net1147 decoded_imm_j\[17\] net970 mem_rdata_q\[17\] VGND VGND VPWR VPWR
+ _06635_ sky130_fd_sc_hd__a22o_1
X_13292_ net556 _02189_ _02210_ _02212_ net391 VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__a311o_1
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09738__A1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12243_ genblk2.pcpi_div.divisor\[6\] net382 net371 net2715 VGND VGND VPWR VPWR _01112_
+ sky130_fd_sc_hd__a22o_1
X_15031_ clknet_leaf_137_clk _01383_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12174_ net751 _06579_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_147_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10405__B net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11125_ cpuregs\[28\]\[21\] cpuregs\[29\]\[21\] net658 VGND VGND VPWR VPWR _05804_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11056_ cpuregs\[18\]\[19\] net554 _05736_ net784 VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_108_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output234_A net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10007_ count_cycle\[4\] _04771_ net1205 VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_160_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10421__A _02379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07206__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14815_ clknet_leaf_79_clk _01167_ VGND VGND VPWR VPWR decoded_imm\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14746_ clknet_leaf_158_clk _01131_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13470__A1 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11958_ net1043 net726 _06423_ net866 VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__a31oi_1
XFILLER_60_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_103_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10909_ cpuregs\[17\]\[15\] net617 net603 _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_15_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14677_ clknet_leaf_162_clk _01062_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11889_ _06283_ _06285_ _06287_ _06289_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08229__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13628_ clknet_leaf_102_clk _00082_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09977__A1 net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13559_ net542 net2417 net411 VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__mux2_1
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11784__A1 net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10587__A2 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07988__B1 net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07080_ net948 _02641_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__or3_1
XANTENNA__09657__A decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07452__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15229_ clknet_leaf_23_clk _01570_ VGND VGND VPWR VPWR cpuregs\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10339__A2 net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__15167__Q mem_rdata_q\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07982_ net988 _03303_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__and3_1
X_09721_ _04513_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__xnor2_1
X_06933_ net1126 genblk2.pcpi_div.quotient\[2\] _02515_ net953 VGND VGND VPWR VPWR
+ _02517_ sky130_fd_sc_hd__a31o_1
XFILLER_68_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08165__B1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13118__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06864_ net1208 _02464_ _02465_ _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__or4_1
XANTENNA__12022__S net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09652_ net1182 net1148 decoded_imm_j\[1\] VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__and3_1
XANTENNA__10511__A2 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08603_ net892 _03976_ _03978_ net2632 net1200 VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__a32o_1
X_09583_ _04417_ net1238 _04416_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__and3b_1
X_06795_ net1031 VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__inv_2
XANTENNA__12957__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08534_ genblk1.genblk1.pcpi_mul.rd\[8\] genblk1.genblk1.pcpi_mul.rdx\[8\] VGND VGND
+ VPWR VPWR _03920_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_121_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08295__X net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12264__A2 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09331__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07640__A net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08465_ _03862_ _03863_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__nor2_1
XANTENNA__07676__C1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_A net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_A net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07416_ reg_pc\[18\] decoded_imm\[18\] VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08396_ reg_out\[16\] alu_out_q\[16\] net1154 VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__mux2_1
XFILLER_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13213__B2 net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07428__C1 _02961_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07347_ net1140 count_cycle\[45\] net977 _02886_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__a211o_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07278_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nor2_1
X_09017_ net305 net1901 net518 VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout899_A net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1227_X net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold150 net60 VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold161 cpuregs\[21\]\[15\] VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 cpuregs\[28\]\[14\] VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 cpuregs\[30\]\[6\] VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 net141 VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout630 net631 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkbuf_4
Xfanout641 net645 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_2
XFILLER_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout652 net654 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_2
X_09919_ _04695_ _04696_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__xnor2_1
Xfanout663 net679 VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__buf_2
XANTENNA__08410__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_X net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout674 net676 VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08156__B1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout685 net687 VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__buf_2
XANTENNA__11337__A net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13028__S net446 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12930_ net1066 _02385_ decoded_imm_j\[11\] _02701_ net710 VGND VGND VPWR VPWR _02120_
+ sky130_fd_sc_hd__a221o_1
Xfanout696 net707 VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10241__A decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11160__C1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10502__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12861_ net283 net2295 net461 VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__mux2_1
XFILLER_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14600_ clknet_leaf_118_clk _00986_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _06279_ _06281_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ clknet_leaf_42_clk _01916_ VGND VGND VPWR VPWR cpuregs\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12792_ net1215 genblk1.genblk1.pcpi_mul.next_rs1\[60\] net1961 net906 net762 VGND
+ VGND VPWR VPWR _01431_ sky130_fd_sc_hd__a221o_1
XANTENNA__12255__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09241__S net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ clknet_leaf_73_clk _00920_ VGND VGND VPWR VPWR decoded_imm_j\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_159_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11743_ net1495 net127 net730 VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14462_ clknet_leaf_64_clk _00851_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dfxtp_1
XANTENNA__12007__A2 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13204__A1 net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11674_ net2671 net737 _06229_ is_alu_reg_imm VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__a22o_1
XFILLER_168_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09959__A1 net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11215__B1 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13413_ net961 _05026_ _02318_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__nor3_1
XANTENNA__06890__B1 _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10625_ net1077 decoded_imm\[7\] net860 VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__o21a_1
X_14393_ clknet_leaf_87_clk _00814_ VGND VGND VPWR VPWR decoder_pseudo_trigger sky130_fd_sc_hd__dfxtp_1
X_10556_ cpuregs\[1\]\[6\] net549 _05249_ net802 net830 VGND VGND VPWR VPWR _05250_
+ sky130_fd_sc_hd__a221o_1
X_13344_ _04996_ _05000_ _05004_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__or3_1
XANTENNA__07434__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13275_ net708 _02173_ _02197_ net564 reg_pc\[9\] VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__a32o_1
X_10487_ net792 _05185_ _05177_ net778 VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__o211a_1
X_15014_ clknet_leaf_107_clk _01366_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_12_0_clk_X clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12226_ net750 net2596 VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__nor2_1
XFILLER_97_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12157_ net2776 net378 net366 net2856 VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__a22o_1
XFILLER_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06945__A1 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11108_ cpuregs\[6\]\[21\] cpuregs\[7\]\[21\] net685 VGND VGND VPWR VPWR _05787_
+ sky130_fd_sc_hd__mux2_1
X_12088_ _06269_ _06368_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08320__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11039_ net831 _05715_ _05719_ net784 VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__a211o_1
XFILLER_65_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13443__A1 net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12246__A2 net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09151__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14729_ clknet_leaf_170_clk _01114_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08250_ reg_out\[2\] reg_next_pc\[2\] net923 VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07201_ _02745_ _02747_ _02748_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_138_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08181_ _03291_ _03670_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand2_1
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11757__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07132_ genblk2.pcpi_div.quotient\[31\] _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__xor2_1
XFILLER_119_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07425__A2 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06804__A net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07063_ genblk2.pcpi_div.quotient\[20\] _02625_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__or2_1
XFILLER_134_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput200 net200 VGND VGND VPWR VPWR pcpi_insn[7] sky130_fd_sc_hd__buf_2
Xoutput211 net1016 VGND VGND VPWR VPWR pcpi_rs1[17] sky130_fd_sc_hd__buf_2
Xoutput222 net999 VGND VGND VPWR VPWR pcpi_rs1[27] sky130_fd_sc_hd__buf_2
Xoutput233 net1034 VGND VGND VPWR VPWR pcpi_rs1[8] sky130_fd_sc_hd__buf_2
Xoutput244 net244 VGND VGND VPWR VPWR pcpi_rs2[18] sky130_fd_sc_hd__buf_2
XANTENNA__07189__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput255 net255 VGND VGND VPWR VPWR pcpi_rs2[28] sky130_fd_sc_hd__buf_2
XANTENNA__10045__B _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07189__B2 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput266 net1167 VGND VGND VPWR VPWR pcpi_rs2[9] sky130_fd_sc_hd__buf_2
XFILLER_114_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09326__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06936__B2 net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07635__A net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13356__B _05748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07965_ _03274_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout382_A net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09704_ _04427_ _04488_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__xor2_1
X_06916_ net1088 _02492_ _02494_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__and3_1
X_07896_ _03351_ _03413_ _03412_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09635_ net3059 net881 _04444_ net851 VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__a22o_1
X_06847_ net33 net134 VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__nand2_2
XFILLER_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout647_A net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13372__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09566_ net3013 _04404_ net1240 VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12237__A2 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06778_ net2768 VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__inv_2
XANTENNA__13434__A1 net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09061__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10248__A1 net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08517_ _03897_ _03900_ _03902_ _03904_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__o211a_1
X_09497_ _04362_ net1239 _04361_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout814_A net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_X net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11996__A1 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_X net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08448_ reg_out\[26\] alu_out_q\[26\] net1155 VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__mux2_1
XFILLER_11_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07664__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08379_ net351 net2370 net528 VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout602_X net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12716__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11620__A mem_rdata_q\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10410_ net252 net251 _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__or3_1
XFILLER_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11390_ cpuregs\[20\]\[28\] cpuregs\[21\]\[28\] net688 VGND VGND VPWR VPWR _06062_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08405__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10341_ cpuregs\[3\]\[31\] net638 net599 _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__o211a_1
XANTENNA__10236__A decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13060_ net1614 net83 net533 VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__mux2_1
X_10272_ _04929_ _04931_ _04930_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10708__C1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12011_ _06297_ _06346_ _06352_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__and3_1
XANTENNA__13370__B1 net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09236__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 _02118_ VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__buf_2
XFILLER_120_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout471 net472 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__buf_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout482 _04291_ VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13962_ clknet_leaf_52_clk _00416_ VGND VGND VPWR VPWR cpuregs\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xfanout493 _04286_ VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_4
XFILLER_74_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09877__B1 net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10487__A1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12913_ net335 net2449 net455 VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__mux2_1
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12597__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13893_ clknet_leaf_30_clk _00347_ VGND VGND VPWR VPWR cpuregs\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13282__A net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15632_ clknet_leaf_190_clk _01968_ VGND VGND VPWR VPWR cpuregs\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12844_ net347 net2245 net459 VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__mux2_1
XFILLER_64_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13425__A1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15563_ clknet_leaf_22_clk _01899_ VGND VGND VPWR VPWR cpuregs\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12775_ net1220 genblk1.genblk1.pcpi_mul.next_rs1\[43\] net2107 net909 net764 VGND
+ VGND VPWR VPWR _01414_ sky130_fd_sc_hd__a221o_1
XANTENNA__08301__A0 net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11987__A1 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14514_ clknet_leaf_79_clk _00903_ VGND VGND VPWR VPWR decoded_imm_j\[10\] sky130_fd_sc_hd__dfxtp_1
X_11726_ net1834 _06241_ net536 VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__mux2_1
X_15494_ clknet_leaf_56_clk _01830_ VGND VGND VPWR VPWR cpuregs\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14445_ clknet_leaf_98_clk _00834_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dfxtp_2
X_11657_ decoded_imm_j\[15\] net7 net546 VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__mux2_1
XANTENNA__11739__A1 net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10608_ _05299_ _05300_ net814 VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__mux2_1
X_14376_ clknet_leaf_132_clk _00797_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dfxtp_4
X_11588_ net3024 net561 net732 _06192_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__a22o_1
XFILLER_155_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13327_ _02238_ _02242_ _02243_ net395 net1020 VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__o32a_1
Xhold908 cpuregs\[18\]\[22\] VGND VGND VPWR VPWR net2222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 genblk1.genblk1.pcpi_mul.next_rs1\[47\] VGND VGND VPWR VPWR net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ cpuregs\[22\]\[5\] cpuregs\[23\]\[5\] net678 VGND VGND VPWR VPWR _05234_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13258_ net1044 net753 _02182_ net708 VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__o211a_1
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13361__B1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12209_ net2893 net270 net2926 VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10433__X _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ net1604 net308 net428 VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__mux2_1
XANTENNA__09146__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1608 instr_andi VGND VGND VPWR VPWR net2922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1619 genblk2.pcpi_div.quotient\[8\] VGND VGND VPWR VPWR net2933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07750_ _03266_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__nand2_1
XFILLER_37_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07681_ cpuregs\[14\]\[3\] cpuregs\[15\]\[3\] net660 VGND VGND VPWR VPWR _03201_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09420_ count_instr\[5\] _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__or2_1
XANTENNA__12219__A2 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09351_ net1630 net322 net476 VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__mux2_1
XANTENNA__15180__Q mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08302_ reg_out\[28\] reg_next_pc\[28\] net925 VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__mux2_1
X_09282_ net1822 net324 net486 VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__mux2_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08233_ net1180 net1161 net940 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__mux2_1
XFILLER_165_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10650__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12536__A net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08164_ _03272_ _03656_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__nor2_1
XFILLER_147_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07115_ net952 _02668_ _02669_ _02671_ _02672_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__a32o_1
XFILLER_109_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08095_ _03589_ _03594_ net989 VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__mux2_1
XANTENNA__12970__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08071__A2 net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1137_A net1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_152_clk VGND VGND VPWR VPWR clkload70/Y sky130_fd_sc_hd__clkinv_4
X_07046_ genblk2.pcpi_div.dividend\[17\] _02603_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__or2_1
Xclkload81 clknet_leaf_134_clk VGND VGND VPWR VPWR clkload81/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_161_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload92 clknet_leaf_143_clk VGND VGND VPWR VPWR clkload92/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13352__B1 net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10490__S net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10166__B1 net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11363__C1 net858 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09056__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07365__A _02898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout385_X net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08997_ net572 net1927 net518 VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__mux2_1
XFILLER_69_970 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07948_ net929 net771 _03279_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout931_A _03462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_X net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07879_ net1160 _02408_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__or2_1
XANTENNA__11130__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11615__A mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09618_ _03803_ reg_next_pc\[15\] net920 VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__mux2_1
XANTENNA__13407__A1 net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10890_ net809 _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__or2_1
X_09549_ _02373_ _04393_ _04395_ net1214 VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_80_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout817_X net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12560_ _05117_ net720 _02399_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11511_ net2636 mem_rdata_q\[4\] net746 VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__mux2_1
XANTENNA__10665__S net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12491_ net2669 net386 _06713_ _06714_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13041__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14230_ clknet_leaf_174_clk _00684_ VGND VGND VPWR VPWR reg_next_pc\[7\] sky130_fd_sc_hd__dfxtp_1
X_11442_ cpuregs\[1\]\[30\] net637 net612 _06111_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__o211a_1
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10929__C1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11373_ net805 _06044_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14161_ clknet_leaf_126_clk _00615_ VGND VGND VPWR VPWR count_instr\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10324_ _04898_ _05026_ _05027_ _04897_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__o31a_1
X_13112_ net349 net2138 net435 VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__mux2_1
XANTENNA__07270__B1 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14092_ clknet_leaf_51_clk _00546_ VGND VGND VPWR VPWR cpuregs\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ net1419 net66 net535 VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__mux2_1
X_10255_ _04947_ _04960_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__nand2_1
Xfanout1200 net1204 VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__buf_2
XANTENNA__07275__A _02814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1211 net1222 VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10186_ decoded_imm\[30\] net992 VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__nor2_1
Xfanout1222 _02378_ VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__buf_2
Xfanout1233 net1234 VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10413__B net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14994_ clknet_leaf_148_clk _01346_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[41\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout290 _03860_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_1
XANTENNA__11657__A0 decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13945_ clknet_leaf_190_clk _00399_ VGND VGND VPWR VPWR cpuregs\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkload6_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13876_ clknet_leaf_178_clk _00330_ VGND VGND VPWR VPWR cpuregs\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15615_ clknet_leaf_71_clk _01951_ VGND VGND VPWR VPWR cpuregs\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10880__A1 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12827_ net285 net1724 net465 VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__mux2_1
XFILLER_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15546_ clknet_leaf_12_clk _01882_ VGND VGND VPWR VPWR cpuregs\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12758_ net1216 genblk1.genblk1.pcpi_mul.next_rs1\[28\] net917 net995 VGND VGND VPWR
+ VPWR _02113_ sky130_fd_sc_hd__a22o_1
XANTENNA__07628__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10632__A1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11709_ net2442 net304 net375 VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15477_ clknet_leaf_195_clk _01813_ VGND VGND VPWR VPWR cpuregs\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12689_ net1203 genblk1.genblk1.pcpi_mul.next_rs2\[54\] net895 net2905 net713 VGND
+ VGND VPWR VPWR _01359_ sky130_fd_sc_hd__a221o_1
X_14428_ clknet_leaf_67_clk alu_out\[28\] VGND VGND VPWR VPWR alu_out_q\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold705 cpuregs\[16\]\[10\] VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__A2 net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14359_ clknet_leaf_80_clk _00780_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
Xhold716 cpuregs\[5\]\[12\] VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold727 cpuregs\[8\]\[22\] VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09665__A decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold738 cpuregs\[27\]\[22\] VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 cpuregs\[4\]\[1\] VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12137__A1 net1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08920_ _04178_ _04180_ _04177_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__a21bo_1
XFILLER_69_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10604__A net790 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08851_ genblk1.genblk1.pcpi_mul.next_rs2\[58\] net1105 genblk1.genblk1.pcpi_mul.rd\[57\]
+ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__a21o_1
XANTENNA__15175__Q mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1405 genblk2.pcpi_div.divisor\[16\] VGND VGND VPWR VPWR net2719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1416 genblk1.genblk1.pcpi_mul.next_rs2\[28\] VGND VGND VPWR VPWR net2730 sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ net1158 net1007 VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__nand2_1
Xhold1427 reg_next_pc\[13\] VGND VGND VPWR VPWR net2741 sky130_fd_sc_hd__dlygate4sd3_1
X_08782_ _04128_ _04129_ _04123_ _04126_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__a211o_1
Xhold1438 genblk1.genblk1.pcpi_mul.next_rs2\[19\] VGND VGND VPWR VPWR net2752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1449 genblk1.genblk1.pcpi_mul.next_rs2\[20\] VGND VGND VPWR VPWR net2763 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09604__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11648__A0 decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07733_ cpuregs\[26\]\[4\] net698 VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__or2_1
XANTENNA__13126__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11435__A net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07632__B net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07664_ cpuregs\[25\]\[2\] net641 net614 _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__o211a_1
X_09403_ net267 net1233 _02437_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__and3_1
XFILLER_38_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14519__Q decoded_imm_j\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07595_ net24 net939 net937 VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12965__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09069__A1 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A _03802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1301 VGND VGND VPWR VPWR picorv32_1301/HI trace_data[23] sky130_fd_sc_hd__conb_1
XANTENNA_fanout1087_A cpu_state\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_1312 VGND VGND VPWR VPWR picorv32_1312/HI trace_data[34] sky130_fd_sc_hd__conb_1
X_09334_ net1706 net577 net476 VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__mux2_1
XANTENNA__07619__A2 decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10993__B _05675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_0_0_clk_X clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09265_ net1830 net581 net487 VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout512_A net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08216_ net1050 net1053 _02688_ net940 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__a211o_2
XFILLER_154_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09196_ _04275_ _04281_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__nor2_2
XANTENNA__11179__A2 _05855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08147_ net966 _03640_ _03293_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout1042_X net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload170 clknet_leaf_88_clk VGND VGND VPWR VPWR clkload170/Y sky130_fd_sc_hd__clkinv_4
X_08078_ net771 _03578_ _03579_ _03573_ VGND VGND VPWR VPWR alu_out\[16\] sky130_fd_sc_hd__a31o_1
Xclkload181 clknet_leaf_101_clk VGND VGND VPWR VPWR clkload181/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout881_A net882 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12128__A1 net993 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07029_ genblk2.pcpi_div.quotient\[14\] genblk2.pcpi_div.quotient\[15\] _02587_ VGND
+ VGND VPWR VPWR _02599_ sky130_fd_sc_hd__or3_1
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07807__B net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10040_ net2988 _04791_ _04793_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_73_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07555__A1 net1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10233__B net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold10 cpuregs\[0\]\[19\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__A2 net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold21 genblk1.genblk1.pcpi_mul.next_rs1\[10\] VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07555__B2 net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold32 cpuregs\[30\]\[18\] VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold43 cpuregs\[24\]\[9\] VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 cpuregs\[24\]\[17\] VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 cpuregs\[24\]\[14\] VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 cpuregs\[24\]\[20\] VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold87 cpuregs\[24\]\[21\] VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold98 cpuregs\[12\]\[25\] VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ genblk2.pcpi_div.dividend\[9\] net271 _06452_ VGND VGND VPWR VPWR _01018_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout934_X net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08197__Y alu_out\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13036__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13730_ clknet_leaf_116_clk _00184_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10942_ cpuregs\[18\]\[16\] net552 _05625_ net779 VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__o22a_1
XFILLER_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13661_ clknet_leaf_108_clk _00115_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10873_ cpuregs\[19\]\[14\] net625 net593 VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__o21a_1
XFILLER_44_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15400_ clknet_leaf_30_clk _01739_ VGND VGND VPWR VPWR cpuregs\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12612_ net1200 net2914 net893 genblk1.genblk1.pcpi_mul.next_rs2\[4\] _02055_ VGND
+ VGND VPWR VPWR _01310_ sky130_fd_sc_hd__a221o_1
XANTENNA__11999__B net1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13592_ net1317 VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15331_ clknet_leaf_54_clk _01671_ VGND VGND VPWR VPWR cpuregs\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12543_ _05114_ net719 _02396_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12176__A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15262_ clknet_leaf_41_clk _01603_ VGND VGND VPWR VPWR cpuregs\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12474_ net2533 net868 VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14213_ clknet_leaf_76_clk _00667_ VGND VGND VPWR VPWR reg_pc\[21\] sky130_fd_sc_hd__dfxtp_1
X_11425_ cpuregs\[20\]\[29\] cpuregs\[21\]\[29\] net706 VGND VGND VPWR VPWR _06096_
+ sky130_fd_sc_hd__mux2_1
X_15193_ clknet_leaf_4_clk _01542_ VGND VGND VPWR VPWR cpuregs\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ clknet_leaf_110_clk _00598_ VGND VGND VPWR VPWR count_instr\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11356_ cpuregs\[16\]\[27\] net692 VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__or2_1
XANTENNA__12623__B net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12119__B2 net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13316__B1 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10307_ _04908_ _05012_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nand2_1
X_14075_ clknet_leaf_197_clk _00529_ VGND VGND VPWR VPWR cpuregs\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11287_ net836 _05957_ _05959_ _05961_ net794 VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__a2111o_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ net308 net2465 net444 VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__mux2_1
X_10238_ decoded_imm\[5\] net1040 VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__and2_1
Xfanout1030 net204 VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11342__A2 net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1041 net230 VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__buf_2
XFILLER_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10169_ count_cycle\[61\] net2991 _04873_ _04876_ net1209 VGND VGND VPWR VPWR _00771_
+ sky130_fd_sc_hd__a311oi_1
Xfanout1052 net1053 VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08388__X _03802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1063 net1064 VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__buf_2
Xfanout1074 cpu_state\[4\] VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1085 net1086 VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1096 net1100 VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__buf_2
X_14977_ clknet_leaf_116_clk _01329_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13928_ clknet_leaf_33_clk _00382_ VGND VGND VPWR VPWR cpuregs\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_164_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13859_ clknet_leaf_12_clk _00313_ VGND VGND VPWR VPWR cpuregs\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12055__B1 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07380_ count_cycle\[15\] net971 VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__or2_1
XFILLER_148_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_179_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15529_ clknet_leaf_19_clk _01865_ VGND VGND VPWR VPWR cpuregs\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_09050_ net309 net2422 net513 VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08001_ _03318_ _03510_ _03465_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold502 cpuregs\[16\]\[12\] VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 net44 VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 cpuregs\[8\]\[29\] VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11030__A1 net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07234__B1 net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06812__A net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold535 cpuregs\[26\]\[11\] VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 cpuregs\[13\]\[22\] VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 cpuregs\[30\]\[5\] VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__A2 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold568 cpuregs\[21\]\[22\] VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _04723_ _04724_ _04725_ net1150 VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__o31ai_1
Xhold579 cpuregs\[10\]\[11\] VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07627__B net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10334__A is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08903_ net1202 net2621 net896 _04228_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09883_ _04662_ _04663_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__nor2_1
XANTENNA__11333__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1202 _00195_ VGND VGND VPWR VPWR net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08834_ _04172_ _04173_ _04167_ _04170_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__a211o_1
Xhold1213 genblk1.genblk1.pcpi_mul.rs2\[63\] VGND VGND VPWR VPWR net2527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1224 cpuregs\[21\]\[1\] VGND VGND VPWR VPWR net2538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10988__B net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1235 genblk1.genblk1.pcpi_mul.pcpi_rd\[12\] VGND VGND VPWR VPWR net2549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 reg_next_pc\[7\] VGND VGND VPWR VPWR net2560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09334__S net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1257 genblk2.pcpi_div.divisor\[38\] VGND VGND VPWR VPWR net2571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13364__B _05784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08765_ net1193 net2967 net886 _04115_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout462_A _02118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1268 count_instr\[34\] VGND VGND VPWR VPWR net2582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1279 reg_next_pc\[6\] VGND VGND VPWR VPWR net2593 sky130_fd_sc_hd__dlygate4sd3_1
X_07716_ cpuregs\[2\]\[4\] cpuregs\[3\]\[4\] net697 VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__mux2_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08696_ genblk1.genblk1.pcpi_mul.rd\[33\] genblk1.genblk1.pcpi_mul.next_rs2\[34\]
+ net1101 VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__and3_1
XFILLER_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07647_ net1080 decoded_imm_j\[19\] VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__or2_1
XFILLER_26_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13380__A net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07578_ _03099_ _03100_ _03101_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o21bai_1
X_09317_ net2271 net325 net481 VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__mux2_1
XFILLER_167_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout515_X net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09248_ net1810 net328 net488 VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__mux2_1
XFILLER_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10228__B net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
X_09179_ net342 net2037 net497 VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__mux2_1
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11210_ cpuregs\[11\]\[23\] net623 net592 _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_75_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12190_ net749 net2934 VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07818__A net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11572__A2 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11141_ _05793_ _05802_ _05819_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__a21oi_4
Xoutput44 net44 VGND VGND VPWR VPWR mem_addr[19] sky130_fd_sc_hd__buf_2
XANTENNA__10244__A net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput55 net55 VGND VGND VPWR VPWR mem_addr[2] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VGND VGND VPWR VPWR mem_la_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput77 net77 VGND VGND VPWR VPWR mem_la_addr[21] sky130_fd_sc_hd__buf_2
X_11072_ cpuregs\[28\]\[20\] cpuregs\[29\]\[20\] net661 VGND VGND VPWR VPWR _05752_
+ sky130_fd_sc_hd__mux2_1
Xoutput88 net88 VGND VGND VPWR VPWR mem_la_addr[31] sky130_fd_sc_hd__buf_2
XANTENNA__07528__A1 net1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput99 net99 VGND VGND VPWR VPWR mem_la_wdata[11] sky130_fd_sc_hd__buf_2
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12473__B1_N net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11774__S net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07528__B2 net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14900_ clknet_leaf_143_clk _01252_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_10023_ count_cycle\[10\] _04781_ net1205 VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_158_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09244__S net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input23_A mem_rdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14831_ clknet_leaf_184_clk _01183_ VGND VGND VPWR VPWR cpuregs\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14762_ clknet_leaf_137_clk _00047_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11974_ genblk2.pcpi_div.dividend\[6\] _06438_ net276 VGND VGND VPWR VPWR _01015_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12488__B1_N net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13713_ clknet_leaf_119_clk _00167_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10925_ net825 _05604_ _05608_ net782 VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__a211o_1
X_14693_ clknet_leaf_139_clk _01078_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13290__A net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13644_ clknet_leaf_151_clk _00098_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10856_ cpuregs\[9\]\[14\] net619 net604 _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__o211a_1
XANTENNA__13234__C1 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_167_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ net316 net2374 net413 VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__mux2_1
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10787_ cpuregs\[6\]\[12\] cpuregs\[7\]\[12\] net652 VGND VGND VPWR VPWR _05475_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11014__S net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15314_ clknet_leaf_4_clk _01654_ VGND VGND VPWR VPWR cpuregs\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12526_ _02015_ _02016_ net2600 net385 VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11949__S net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15245_ clknet_leaf_14_clk _01586_ VGND VGND VPWR VPWR cpuregs\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__A1 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12457_ net1172 _05099_ net717 net865 VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_169_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output91_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11408_ cpuregs\[14\]\[29\] cpuregs\[15\]\[29\] net704 VGND VGND VPWR VPWR _06079_
+ sky130_fd_sc_hd__mux2_1
X_15176_ clknet_leaf_90_clk _01525_ VGND VGND VPWR VPWR mem_rdata_q\[27\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__08323__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12388_ net1597 net282 net363 VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__mux2_1
XANTENNA__14622__Q genblk2.pcpi_div.outsign VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14127_ clknet_leaf_92_clk _00581_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dfxtp_2
XANTENNA__12760__B2 net993 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11339_ cpuregs\[8\]\[27\] net693 VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__or2_1
XFILLER_125_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14058_ clknet_leaf_52_clk _00512_ VGND VGND VPWR VPWR cpuregs\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11315__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11684__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13009_ net538 net2394 net443 VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__mux2_1
XFILLER_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06880_ net1185 net850 VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__nand2_1
XANTENNA__09154__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08550_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__inv_2
XANTENNA__07182__B decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08993__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07501_ net1073 _03022_ _03023_ _03030_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__a31o_1
X_08481_ genblk1.genblk1.pcpi_mul.instr_mulhsu genblk1.genblk1.pcpi_mul.instr_mulh
+ _03876_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__o21a_1
XFILLER_51_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07432_ _02951_ _02956_ _02965_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_18_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07363_ genblk1.genblk1.pcpi_mul.pcpi_rd\[14\] genblk2.pcpi_div.pcpi_rd\[14\] net1110
+ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__mux2_1
XANTENNA__10329__A net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09102_ net1668 net523 net505 VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__mux2_1
X_07294_ _02821_ _02825_ _02835_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13528__A0 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09033_ net537 net2297 net512 VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09329__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold310 cpuregs\[24\]\[24\] VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 net166 VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08233__S net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold332 net51 VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold343 cpuregs\[15\]\[7\] VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14532__Q decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold354 cpuregs\[21\]\[8\] VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold365 cpuregs\[22\]\[27\] VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10762__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold376 cpuregs\[15\]\[21\] VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 cpuregs\[22\]\[17\] VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold398 cpuregs\[30\]\[8\] VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net802 VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__clkbuf_4
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09853__A net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout812 net821 VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__buf_2
X_09935_ _04445_ _04446_ _04691_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__nand3_1
Xfanout823 net826 VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout834 _03137_ VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout677_A net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout845 net846 VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__buf_2
XFILLER_58_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout856 net859 VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__clkbuf_4
Xfanout867 net869 VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__clkbuf_4
X_09866_ net984 _04643_ _04644_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__o31ai_1
Xfanout878 net882 VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__buf_2
Xhold1010 cpuregs\[12\]\[24\] VGND VGND VPWR VPWR net2324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1005_X net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1021 cpuregs\[10\]\[27\] VGND VGND VPWR VPWR net2335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09064__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout889 net890 VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1032 cpuregs\[1\]\[21\] VGND VGND VPWR VPWR net2346 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net1203 net2995 net895 _04159_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__a22o_1
Xhold1043 cpuregs\[19\]\[19\] VGND VGND VPWR VPWR net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1054 _01428_ VGND VGND VPWR VPWR net2368 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A _02702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09797_ _04582_ _04583_ net1149 VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__o21a_1
Xhold1065 cpuregs\[18\]\[18\] VGND VGND VPWR VPWR net2379 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1076 cpuregs\[19\]\[6\] VGND VGND VPWR VPWR net2390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08748_ genblk1.genblk1.pcpi_mul.rd\[41\] genblk1.genblk1.pcpi_mul.next_rs2\[42\]
+ net1091 VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__and3_1
Xhold1087 cpuregs\[5\]\[14\] VGND VGND VPWR VPWR net2401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 cpuregs\[17\]\[20\] VGND VGND VPWR VPWR net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10817__A1 net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08679_ _04035_ _04038_ _04040_ _04041_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__o211a_1
XANTENNA__10938__S net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09683__A1 net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_X net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09683__B2 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ cpuregs\[9\]\[10\] net628 net607 _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__o211a_1
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07694__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07820__B net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11690_ net1982 net540 net374 VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__mux2_1
XANTENNA__08408__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12438__B _02507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10641_ net789 _05328_ _05330_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_101_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__A decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13360_ net709 _02248_ _02270_ _02272_ net392 VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__a311o_1
XFILLER_166_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10572_ cpuregs\[26\]\[6\] net677 VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12311_ decoded_imm\[18\] net743 _06632_ _06634_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__o22a_1
XFILLER_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13291_ net708 _02190_ _02211_ net564 reg_pc\[11\] VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__a32o_1
XANTENNA__09239__S net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15030_ clknet_leaf_137_clk _01382_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_12242_ net2734 net382 net371 net2887 VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__a22o_1
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12173_ net2602 net277 net2746 VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_147_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11124_ cpuregs\[30\]\[21\] cpuregs\[31\]\[21\] net658 VGND VGND VPWR VPWR _05803_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11055_ cpuregs\[19\]\[19\] net632 net597 VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__o21a_1
XFILLER_77_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input26_X net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10006_ _04771_ _04772_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_125_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output227_A net1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10421__B net880 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14814_ clknet_leaf_78_clk _01166_ VGND VGND VPWR VPWR decoded_imm\[8\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__12258__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14745_ clknet_leaf_158_clk _01130_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11957_ net726 _06423_ net1043 VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__a21o_1
X_10908_ cpuregs\[16\]\[15\] net646 VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__or2_1
X_14676_ clknet_leaf_162_clk net2795 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11888_ _06289_ _06358_ _06287_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_15_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13627_ clknet_leaf_98_clk net945 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_ready
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08229__A2 net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10839_ net772 _05517_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__and3_1
XFILLER_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13558_ net574 net2436 net414 VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07988__A1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11679__S net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11784__A2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12509_ genblk2.pcpi_div.divisor\[48\] net870 VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__or2_1
XFILLER_146_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13489_ net2113 net583 net421 VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09149__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15228_ clknet_leaf_22_clk _01569_ VGND VGND VPWR VPWR cpuregs\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12733__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15159_ clknet_leaf_89_clk _01508_ VGND VGND VPWR VPWR mem_rdata_q\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07981_ _03274_ _03304_ _03487_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__or3_1
X_09720_ _04503_ _04505_ _04502_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__a21oi_1
X_06932_ net1126 _02515_ genblk2.pcpi_div.quotient\[2\] VGND VGND VPWR VPWR _02516_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_79_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09651_ reg_pc\[31\] net879 _04452_ net849 VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__a22o_1
X_06863_ _02457_ _02461_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__nand2_1
X_08602_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__inv_2
XANTENNA__12249__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09582_ count_instr\[61\] count_instr\[60\] _04413_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__and3_1
X_06794_ net1044 VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__inv_2
XANTENNA__09612__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08533_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__inv_2
XFILLER_70_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13134__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08464_ reg_pc\[29\] reg_pc\[28\] _03855_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__and3_1
X_07415_ _02950_ _02945_ _02943_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_34_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ net339 net2204 net528 VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__mux2_1
XFILLER_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12973__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_A net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout1167_A net266 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11224__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07346_ count_instr\[45\] net1131 net1136 count_instr\[13\] VGND VGND VPWR VPWR _02886_
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07277_ reg_pc\[9\] decoded_imm\[9\] VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nand2_1
X_09016_ net308 net1969 net517 VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__mux2_1
XFILLER_152_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout794_A net795 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold140 cpuregs\[23\]\[15\] VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 decoded_rd\[1\] VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 cpuregs\[12\]\[14\] VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 cpuregs\[26\]\[28\] VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 cpuregs\[20\]\[30\] VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 cpuregs\[31\]\[21\] VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A _02462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout620 net645 VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkbuf_2
Xfanout631 net645 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11618__A mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout642 net644 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkbuf_4
X_09918_ _04686_ _04688_ _04684_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__a21o_1
XFILLER_120_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout653 net654 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__clkbuf_2
Xfanout664 net672 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 net676 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout686 net687 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09849_ net1146 _04632_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__nand2_1
Xfanout697 net701 VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10241__B net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07364__C1 _02901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_X net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12860_ net285 net2104 net462 VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__mux2_1
XFILLER_18_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11811_ _06279_ _06280_ _06281_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07831__A net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ net1215 net2476 net2508 net906 net762 VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12449__A _02392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ clknet_leaf_73_clk _00919_ VGND VGND VPWR VPWR decoded_imm_j\[1\] sky130_fd_sc_hd__dfxtp_2
X_11742_ net1700 net1170 net729 VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__mux2_1
XANTENNA__11463__A1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14461_ clknet_leaf_65_clk _00850_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dfxtp_1
X_11673_ mem_rdata_q\[30\] _02388_ net737 _06179_ _06196_ VGND VGND VPWR VPWR _06229_
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13204__A2 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13412_ _04902_ _05025_ _04900_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__o21a_1
XANTENNA__11215__A1 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06890__A1 net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10624_ net1077 _05316_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__nand2_1
XFILLER_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06890__B2 net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14392_ clknet_leaf_86_clk _00813_ VGND VGND VPWR VPWR latched_branch sky130_fd_sc_hd__dfxtp_1
X_13343_ net1017 net396 _02252_ _02257_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__o22a_1
X_10555_ cpuregs\[2\]\[6\] cpuregs\[3\]\[6\] net674 VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__mux2_1
XFILLER_155_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12184__A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10974__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13274_ _02406_ net752 VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__nand2_1
X_10486_ net831 _05180_ _05182_ _05184_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a211o_1
XFILLER_154_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15013_ clknet_leaf_107_clk net2959 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_12225_ genblk2.pcpi_div.quotient_msk\[26\] net275 net2595 VGND VGND VPWR VPWR _06605_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12191__A2 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12156_ genblk2.pcpi_div.quotient_msk\[15\] net378 net367 net2776 VGND VGND VPWR
+ VPWR _01057_ sky130_fd_sc_hd__a22o_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06910__A net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12631__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11107_ net247 net856 _05785_ _05786_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__a22o_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12087_ net3050 _06534_ net273 VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__mux2_1
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08147__A1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07217__S net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11038_ cpuregs\[3\]\[19\] net632 net597 _05718_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__o211a_1
XFILLER_65_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06909__X _02501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07370__A2 decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12989_ net1541 net318 net448 VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__mux2_1
XANTENNA__09647__B2 net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13443__A2 net757 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14728_ clknet_leaf_170_clk _01113_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08048__S net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14659_ clknet_leaf_141_clk _01044_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_180_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_180_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07200_ _02745_ _02747_ _02748_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__a21o_1
XANTENNA__11206__A1 net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08180_ _03291_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__or2_1
X_07131_ genblk2.pcpi_div.quotient\[29\] genblk2.pcpi_div.quotient\[30\] _02671_ net1123
+ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_41_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07062_ _02623_ _02624_ _02626_ _02627_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__o22ai_1
XANTENNA__07188__A net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 net201 VGND VGND VPWR VPWR pcpi_insn[8] sky130_fd_sc_hd__buf_2
XANTENNA__15178__Q mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput212 net1015 VGND VGND VPWR VPWR pcpi_rs1[18] sky130_fd_sc_hd__buf_2
Xoutput223 net997 VGND VGND VPWR VPWR pcpi_rs1[28] sky130_fd_sc_hd__buf_2
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput234 net234 VGND VGND VPWR VPWR pcpi_rs1[9] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR pcpi_rs2[19] sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR pcpi_rs2[29] sky130_fd_sc_hd__buf_2
XANTENNA__07189__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput267 net267 VGND VGND VPWR VPWR pcpi_valid sky130_fd_sc_hd__buf_2
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13129__S net438 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14810__Q decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07635__B net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07964_ _03273_ net930 net968 VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__o21a_1
XFILLER_68_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09703_ _04496_ _04497_ _04498_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__o21a_1
X_06915_ _02494_ _02505_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__and2_1
X_07895_ net1168 net1033 VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12968__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A net376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09634_ _03837_ reg_next_pc\[23\] net926 VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__mux2_2
X_06846_ net33 net134 VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__and2_1
XANTENNA__12890__A0 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09342__S net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13372__B _05820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09565_ count_instr\[55\] count_instr\[54\] _04403_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__and3_1
X_06777_ reg_sh\[0\] VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__inv_2
XANTENNA__13434__A2 net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11445__A1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ _03902_ _03904_ _03897_ _03900_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__a211o_1
XANTENNA__10248__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ count_instr\[30\] count_instr\[29\] _04358_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__and3_1
XFILLER_169_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08447_ net301 net2247 net531 VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_171_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_171_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1072_X net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout428_X net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A _03143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08378_ _03792_ _03793_ net766 VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__mux2_1
XFILLER_165_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12716__B net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11620__B mem_rdata_q\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07329_ _02811_ _02869_ net1060 VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__o21a_1
XFILLER_165_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10340_ cpuregs\[2\]\[31\] net695 VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__or2_1
XFILLER_137_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout797_X net797 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10236__B net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10271_ _04931_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__nand2_1
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12010_ _06297_ _06346_ _06352_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12173__A2 net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07826__A net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13039__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout450 _02123_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08129__A1 net969 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout461 _02118_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08129__B2 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 _06664_ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__buf_4
X_13961_ clknet_leaf_56_clk _00415_ VGND VGND VPWR VPWR cpuregs\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout494 _04286_ VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12912_ net338 net2365 net455 VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__mux2_1
XANTENNA__12881__A0 mem_rdata_q\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13892_ clknet_leaf_40_clk _00346_ VGND VGND VPWR VPWR cpuregs\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09252__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12843_ net351 net2339 net459 VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__mux2_1
X_15631_ clknet_leaf_182_clk _01967_ VGND VGND VPWR VPWR cpuregs\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09629__B2 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15562_ clknet_leaf_29_clk _01898_ VGND VGND VPWR VPWR cpuregs\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12774_ net1220 genblk1.genblk1.pcpi_mul.next_rs1\[42\] net2504 net908 net764 VGND
+ VGND VPWR VPWR _01413_ sky130_fd_sc_hd__a221o_1
XANTENNA__12633__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14513_ clknet_leaf_79_clk _00902_ VGND VGND VPWR VPWR decoded_imm_j\[9\] sky130_fd_sc_hd__dfxtp_1
X_11725_ mem_do_wdata net982 VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__and2b_1
XFILLER_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15493_ clknet_leaf_54_clk _01829_ VGND VGND VPWR VPWR cpuregs\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_162_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_162_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13502__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14444_ clknet_leaf_90_clk _00833_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dfxtp_1
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11656_ net1405 net3 net548 VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__mux2_1
X_10607_ cpuregs\[20\]\[7\] cpuregs\[21\]\[7\] net668 VGND VGND VPWR VPWR _05300_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14375_ clknet_leaf_134_clk _00796_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dfxtp_1
XFILLER_167_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11587_ net2550 net561 _06192_ _06193_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__a22o_1
XANTENNA__11022__S net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13326_ net567 _05599_ net395 VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__o21ai_1
Xhold909 cpuregs\[5\]\[15\] VGND VGND VPWR VPWR net2223 sky130_fd_sc_hd__dlygate4sd3_1
X_10538_ cpuregs\[20\]\[5\] cpuregs\[21\]\[5\] net678 VGND VGND VPWR VPWR _05233_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13257_ _02404_ net753 VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__nand2_1
X_10469_ net987 _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__nor2_1
XANTENNA__12164__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12208_ net748 net2736 VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__nor2_1
XANTENNA__08331__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13361__B2 net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13188_ net1860 net312 net429 VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__mux2_1
X_12139_ net2663 net1223 _05094_ net749 VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__a31o_1
XFILLER_150_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1609 genblk1.genblk1.pcpi_mul.next_rs2\[22\] VGND VGND VPWR VPWR net2923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11692__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09868__B2 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12872__A0 mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07680_ _03196_ _03199_ net781 VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__a21o_1
XFILLER_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09162__S net503 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12089__A net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09350_ net1797 net326 net477 VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__mux2_1
X_08301_ net998 _03734_ net983 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__mux2_2
XFILLER_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09281_ net1573 net328 net484 VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_153_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_153_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_166_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08232_ net1056 net1169 net1162 _02690_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__a22o_1
XFILLER_21_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14805__Q decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08163_ net1145 _03293_ _03655_ _03654_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__o31a_1
XANTENNA__12028__S net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07114_ genblk2.pcpi_div.quotient\[28\] _02670_ net953 VGND VGND VPWR VPWR _02672_
+ sky130_fd_sc_hd__a21oi_1
X_08094_ _03593_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__inv_2
Xclkload60 clknet_leaf_177_clk VGND VGND VPWR VPWR clkload60/X sky130_fd_sc_hd__clkbuf_8
Xclkload71 clknet_leaf_154_clk VGND VGND VPWR VPWR clkload71/Y sky130_fd_sc_hd__inv_12
X_07045_ net950 _02611_ _02612_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__or3_1
XANTENNA__10771__S net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload82 clknet_leaf_136_clk VGND VGND VPWR VPWR clkload82/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__12552__A net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_A net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload93 clknet_leaf_144_clk VGND VGND VPWR VPWR clkload93/X sky130_fd_sc_hd__clkbuf_8
XFILLER_161_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09337__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13352__B2 net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07646__A net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout492_A net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08996_ net575 net1730 net517 VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__mux2_1
X_07947_ is_compare _02433_ net933 net928 VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__or4_4
XFILLER_130_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12863__A0 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07878_ net253 net1001 VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__and2b_1
XANTENNA__09072__S net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07334__A2 net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09617_ reg_pc\[14\] net875 _04435_ net845 VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__a22o_1
XANTENNA__11615__B mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06829_ instr_lhu instr_lh _02431_ net966 VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout924_A net925 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13407__A2 net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09548_ count_instr\[47\] count_instr\[46\] _04387_ _04394_ VGND VGND VPWR VPWR _04395_
+ sky130_fd_sc_hd__and4_1
XANTENNA__12615__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08295__A0 net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12091__A1 net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09479_ net2998 _04349_ net1239 VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10946__S net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_144_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_144_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout712_X net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11510_ net2612 mem_rdata_q\[3\] net746 VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12490_ net871 _06711_ _06712_ net386 VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__a31oi_1
XANTENNA__08416__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ cpuregs\[0\]\[30\] net691 VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__or2_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10247__A net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14160_ clknet_leaf_94_clk _00614_ VGND VGND VPWR VPWR count_instr\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11372_ cpuregs\[12\]\[28\] cpuregs\[13\]\[28\] net689 VGND VGND VPWR VPWR _06044_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13111_ net352 net2239 net435 VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10323_ _04902_ _04904_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__nor2_1
X_14091_ clknet_leaf_66_clk _00545_ VGND VGND VPWR VPWR cpuregs\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10681__S net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09247__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12146__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13042_ net1334 net95 net535 VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__mux2_1
X_10254_ _04948_ _04958_ _04959_ _04947_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__o211ai_2
XFILLER_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1201 net1204 VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__clkbuf_2
XFILLER_79_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1212 net1214 VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__buf_2
X_10185_ decoded_imm\[30\] net992 VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__and2_1
Xfanout1223 net34 VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__clkbuf_4
Xfanout1234 net1241 VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout280 _03873_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_2
X_14993_ clknet_leaf_145_clk _01345_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11106__B1 net859 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout291 _03860_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11657__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13944_ clknet_leaf_186_clk _00398_ VGND VGND VPWR VPWR cpuregs\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12401__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13875_ clknet_leaf_25_clk _00329_ VGND VGND VPWR VPWR cpuregs\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15614_ clknet_leaf_35_clk _01950_ VGND VGND VPWR VPWR cpuregs\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12826_ net291 net1923 net466 VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__mux2_1
XANTENNA__10880__A2 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12082__A1 net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15545_ clknet_leaf_42_clk _01881_ VGND VGND VPWR VPWR cpuregs\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12757_ net1214 net1578 net2575 net900 _02112_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_135_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_135_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_148_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13232__S net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10093__B1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11708_ net1925 net307 net375 VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__mux2_1
X_15476_ clknet_leaf_195_clk _01812_ VGND VGND VPWR VPWR cpuregs\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08326__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12688_ net1203 net2905 net895 net2977 net713 VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ clknet_leaf_67_clk alu_out\[27\] VGND VGND VPWR VPWR alu_out_q\[27\] sky130_fd_sc_hd__dfxtp_1
X_11639_ net1353 net741 _06222_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14358_ clknet_leaf_131_clk _00779_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
XFILLER_155_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold706 cpuregs\[31\]\[22\] VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold717 cpuregs\[5\]\[17\] VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11687__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold728 net172 VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ net567 _05527_ _02222_ net959 VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__a2bb2o_1
Xhold739 net186 VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ clknet_leaf_126_clk _00743_ VGND VGND VPWR VPWR count_cycle\[34\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12137__A2 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09157__S net503 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14360__Q net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08850_ net901 _04185_ _04187_ net2641 net1211 VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__a32o_1
XANTENNA__08996__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1406 count_cycle\[15\] VGND VGND VPWR VPWR net2720 sky130_fd_sc_hd__dlygate4sd3_1
X_07801_ net1158 net1007 VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__and2_1
Xhold1417 genblk2.pcpi_div.divisor\[21\] VGND VGND VPWR VPWR net2731 sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ genblk1.genblk1.pcpi_mul.rd\[46\] genblk1.genblk1.pcpi_mul.next_rs2\[47\]
+ net1090 VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__nand3_1
Xhold1428 genblk2.pcpi_div.divisor\[10\] VGND VGND VPWR VPWR net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 genblk2.pcpi_div.quotient\[30\] VGND VGND VPWR VPWR net2753 sky130_fd_sc_hd__dlygate4sd3_1
X_07732_ cpuregs\[25\]\[4\] net641 net614 _03250_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__o211a_1
XANTENNA__11648__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07316__A2 net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07663_ cpuregs\[24\]\[2\] net700 VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__or2_1
XFILLER_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09402_ net175 net174 _04299_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__and3_1
X_07594_ _03115_ _03116_ net1072 VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__and3b_1
XFILLER_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09620__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08277__A0 net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09333_ net1451 net582 net477 VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1302 VGND VGND VPWR VPWR picorv32_1302/HI trace_data[24] sky130_fd_sc_hd__conb_1
Xpicorv32_1313 VGND VGND VPWR VPWR picorv32_1313/HI trace_data[35] sky130_fd_sc_hd__conb_1
XANTENNA__13270__B1 net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_126_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13142__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09264_ net2322 net583 net486 VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__mux2_1
XANTENNA__08236__S net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08215_ net1050 _02384_ _02688_ net940 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__a211o_2
X_09195_ net278 net2285 net498 VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__mux2_1
XANTENNA__12981__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout505_A _04279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08146_ _03292_ net931 VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07252__A1 net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08077_ _03343_ _03577_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__nand2_1
Xclkload160 clknet_leaf_120_clk VGND VGND VPWR VPWR clkload160/Y sky130_fd_sc_hd__inv_6
Xclkload171 clknet_leaf_90_clk VGND VGND VPWR VPWR clkload171/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload182 clknet_leaf_103_clk VGND VGND VPWR VPWR clkload182/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_fanout1035_X net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09067__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09529__B1 net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07028_ genblk2.pcpi_div.dividend\[16\] net1114 _02596_ net947 VGND VGND VPWR VPWR
+ _02598_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout495_X net495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A _05082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07555__A2 net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold11 cpuregs\[0\]\[0\] VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 _01380_ VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 net36 VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ net1382 _04266_ net946 VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__mux2_1
Xhold44 cpuregs\[28\]\[24\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 cpuregs\[24\]\[10\] VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 cpuregs\[24\]\[2\] VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 cpuregs\[26\]\[18\] VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _06449_ _06450_ _06451_ net867 net271 VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__o221a_1
Xhold88 cpuregs\[28\]\[1\] VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 cpuregs\[14\]\[4\] VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__A2 decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10847__C1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10941_ cpuregs\[19\]\[16\] net621 net591 VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout927_X net927 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13660_ clknet_leaf_105_clk _00114_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ cpuregs\[17\]\[14\] net625 net607 _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__o211a_1
X_12611_ _02393_ net911 VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__nor2_1
XANTENNA__13261__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13591_ net1324 VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_117_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_169_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13052__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15330_ clknet_leaf_70_clk _01670_ VGND VGND VPWR VPWR cpuregs\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12542_ _02028_ net2581 net389 VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15261_ clknet_leaf_7_clk _01602_ VGND VGND VPWR VPWR cpuregs\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12473_ _05101_ net717 net1167 VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14212_ clknet_leaf_77_clk _00666_ VGND VGND VPWR VPWR reg_pc\[20\] sky130_fd_sc_hd__dfxtp_2
X_11424_ net837 _06090_ _06092_ _06094_ net794 VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09766__A decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15192_ clknet_leaf_5_clk _01541_ VGND VGND VPWR VPWR cpuregs\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13288__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07243__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_110_clk _00597_ VGND VGND VPWR VPWR count_instr\[14\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_89_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11355_ _06026_ _06027_ net805 VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__mux2_1
XFILLER_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12192__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11300__S net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12623__C net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10306_ _04910_ _05011_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__or2_1
X_14074_ clknet_leaf_198_clk _00528_ VGND VGND VPWR VPWR cpuregs\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11286_ cpuregs\[27\]\[25\] net642 net602 _05960_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__o211a_1
X_13025_ net313 net2371 net445 VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ _04941_ _04942_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__nand2_1
XFILLER_105_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1021 VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__clkbuf_4
Xfanout1031 net1032 VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net229 VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__clkbuf_4
X_10168_ count_cycle\[61\] _04873_ net2991 VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1053 net203 VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10550__A1 net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1064 net1065 VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1075 cpu_state\[3\] VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__buf_2
Xfanout1086 net1087 VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1097 net1100 VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__buf_1
X_10099_ net2745 _04830_ net1225 VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__o21ai_1
X_14976_ clknet_leaf_116_clk _01328_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_13927_ clknet_leaf_32_clk _00381_ VGND VGND VPWR VPWR cpuregs\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13858_ clknet_leaf_12_clk _00312_ VGND VGND VPWR VPWR cpuregs\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08259__A0 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ net357 net1914 net463 VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_108_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_8
X_13789_ clknet_leaf_7_clk _00243_ VGND VGND VPWR VPWR cpuregs\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15528_ clknet_leaf_31_clk _01864_ VGND VGND VPWR VPWR cpuregs\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15459_ clknet_leaf_56_clk _01798_ VGND VGND VPWR VPWR cpuregs\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_08000_ _03318_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__nor2_1
XANTENNA__09676__A decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold503 cpuregs\[16\]\[15\] VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13198__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07234__A1 net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11030__A2 _05710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold514 cpuregs\[4\]\[2\] VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 cpuregs\[15\]\[17\] VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold536 cpuregs\[20\]\[14\] VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold547 genblk1.genblk1.pcpi_mul.pcpi_rd\[7\] VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09951_ _04724_ _04725_ _04723_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__o21a_1
Xhold558 cpuregs\[6\]\[18\] VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 cpuregs\[13\]\[13\] VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08902_ _03980_ _03982_ _03979_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_55_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ net1127 _04442_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__nor2_1
XFILLER_112_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08833_ genblk1.genblk1.pcpi_mul.rd\[54\] genblk1.genblk1.pcpi_mul.next_rs2\[55\]
+ net1103 VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__nand3_1
Xhold1203 genblk1.genblk1.pcpi_mul.next_rs1\[46\] VGND VGND VPWR VPWR net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 _01369_ VGND VGND VPWR VPWR net2528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 genblk1.genblk1.pcpi_mul.pcpi_rd\[5\] VGND VGND VPWR VPWR net2539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13137__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1236 instr_sltiu VGND VGND VPWR VPWR net2550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 count_instr\[17\] VGND VGND VPWR VPWR net2561 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ _04113_ _04114_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__xnor2_1
Xhold1258 instr_sltu VGND VGND VPWR VPWR net2572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 _00617_ VGND VGND VPWR VPWR net2583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07715_ net807 _03231_ _03233_ net839 VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__a211o_1
XFILLER_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12976__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08695_ genblk1.genblk1.pcpi_mul.next_rs2\[34\] net1101 genblk1.genblk1.pcpi_mul.rd\[33\]
+ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout455_A net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1197_A net1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07646_ net794 _03164_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09350__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13380__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07577_ _03086_ _03089_ _03088_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout622_A net624 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10057__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09316_ net1864 net330 net479 VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__mux2_1
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09247_ net1701 net332 net488 VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__mux2_1
XANTENNA__07473__A1 net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07473__B2 net1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_X net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_X net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09178_ net346 net2385 net496 VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__mux2_1
XANTENNA__12724__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07225__A1 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08129_ net969 _03321_ _03324_ net931 _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_75_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07818__B net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11140_ net774 _05810_ _05818_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout877_X net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput45 net45 VGND VGND VPWR VPWR mem_addr[20] sky130_fd_sc_hd__buf_2
Xoutput56 net56 VGND VGND VPWR VPWR mem_addr[30] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR mem_la_addr[11] sky130_fd_sc_hd__buf_2
XFILLER_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput78 net78 VGND VGND VPWR VPWR mem_la_addr[22] sky130_fd_sc_hd__buf_2
X_11071_ cpuregs\[30\]\[20\] cpuregs\[31\]\[20\] net661 VGND VGND VPWR VPWR _05751_
+ sky130_fd_sc_hd__mux2_1
Xoutput89 net89 VGND VGND VPWR VPWR mem_la_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07528__A2 net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07834__A net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12521__A2 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10022_ _04781_ _04782_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__nor2_1
XANTENNA__09922__B1 net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13047__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14830_ clknet_leaf_187_clk _01182_ VGND VGND VPWR VPWR cpuregs\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12809__A0 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A mem_rdata[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14761_ clknet_leaf_137_clk _00046_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11973_ net865 _06328_ _06433_ _06437_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__a31o_1
XFILLER_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10924_ cpuregs\[3\]\[16\] net623 net591 _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__o211a_1
X_13712_ clknet_leaf_122_clk _00166_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10835__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07697__D1 net790 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14692_ clknet_leaf_141_clk _01077_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09260__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10855_ cpuregs\[8\]\[14\] net653 VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__or2_1
X_13643_ clknet_leaf_151_clk _00097_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13234__B1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13574_ net320 net2412 net411 VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__mux2_1
X_10786_ net822 _05469_ _05471_ _05473_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a211o_1
XANTENNA__10599__A1 net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15313_ clknet_leaf_3_clk _01653_ VGND VGND VPWR VPWR cpuregs\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12525_ net872 _02013_ _02014_ net388 VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__a31o_1
XANTENNA__11260__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13510__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12456_ _05099_ net717 net1172 VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__a21oi_1
X_15244_ clknet_leaf_41_clk _01585_ VGND VGND VPWR VPWR cpuregs\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11407_ _06075_ _06077_ net786 VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__a21o_1
X_15175_ clknet_leaf_90_clk _01524_ VGND VGND VPWR VPWR mem_rdata_q\[26\] sky130_fd_sc_hd__dfxtp_2
X_12387_ net1403 net288 net362 VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__mux2_1
XANTENNA_output84_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14126_ clknet_leaf_98_clk _00580_ VGND VGND VPWR VPWR genblk2.pcpi_div.instr_remu
+ sky130_fd_sc_hd__dfxtp_1
X_11338_ net817 _06008_ _06010_ net833 VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__o211a_1
X_14057_ clknet_leaf_50_clk _00511_ VGND VGND VPWR VPWR cpuregs\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11269_ cpuregs\[11\]\[25\] net643 net602 _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__o211a_1
XFILLER_97_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13008_ net541 net2243 net444 VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__mux2_1
XANTENNA__09913__B1 net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14959_ clknet_leaf_144_clk _01311_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_07500_ net358 _03024_ _03029_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10287__B1 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08480_ genblk1.genblk1.pcpi_mul.mul_waiting net1189 net1237 VGND VGND VPWR VPWR
+ _03876_ sky130_fd_sc_hd__and3_1
XANTENNA__09170__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07431_ reg_pc\[19\] decoded_imm\[19\] VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13225__A0 net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10039__B1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07362_ count_cycle\[14\] net971 net841 _02900_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__o211a_1
XFILLER_50_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09101_ net1501 net524 net504 VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__mux2_1
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07293_ _02821_ _02825_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__and3_1
X_09032_ net541 net2482 net513 VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__mux2_1
XFILLER_148_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07207__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14813__Q decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold300 net52 VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07207__B2 net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold311 cpuregs\[12\]\[19\] VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10345__A net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold322 cpuregs\[26\]\[1\] VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 cpuregs\[12\]\[20\] VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold344 cpuregs\[22\]\[4\] VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12751__A2 net903 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold355 net152 VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 cpuregs\[12\]\[22\] VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold377 cpuregs\[23\]\[12\] VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__X _06243_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout802 net803 VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__clkbuf_4
XFILLER_77_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold388 cpuregs\[21\]\[24\] VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 cpuregs\[29\]\[18\] VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _04446_ _04699_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__or2_1
Xfanout813 net815 VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1112_A genblk2.pcpi_div.pcpi_ready VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout824 net825 VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09345__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout835 net837 VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net852 VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__A2 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A mem_rdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout857 net858 VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__buf_2
X_09865_ _04440_ _04634_ _04647_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__o21ai_1
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1000 cpuregs\[7\]\[29\] VGND VGND VPWR VPWR net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout572_A _03761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout879 net880 VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__buf_2
Xhold1011 cpuregs\[17\]\[18\] VGND VGND VPWR VPWR net2325 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__A2 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1022 cpuregs\[7\]\[21\] VGND VGND VPWR VPWR net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 cpuregs\[7\]\[14\] VGND VGND VPWR VPWR net2347 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _04157_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__xnor2_1
Xhold1044 cpuregs\[17\]\[14\] VGND VGND VPWR VPWR net2358 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _04582_ _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__nand2_1
XFILLER_39_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1055 cpuregs\[13\]\[24\] VGND VGND VPWR VPWR net2369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A2 net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1066 cpuregs\[19\]\[14\] VGND VGND VPWR VPWR net2380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08747_ genblk1.genblk1.pcpi_mul.next_rs2\[42\] net1092 genblk1.genblk1.pcpi_mul.rd\[41\]
+ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__a21o_1
Xhold1077 cpuregs\[9\]\[21\] VGND VGND VPWR VPWR net2391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1088 cpuregs\[5\]\[9\] VGND VGND VPWR VPWR net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1099 cpuregs\[1\]\[28\] VGND VGND VPWR VPWR net2413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout458_X net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A _03137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08678_ _04040_ _04041_ _04035_ _04038_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__a211o_1
XANTENNA__08485__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07143__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09080__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__A1 net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07629_ net1080 decoded_imm_j\[18\] VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__or2_1
XFILLER_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10640_ cpuregs\[11\]\[8\] net626 net593 _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__o211a_1
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__B net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10571_ cpuregs\[25\]\[6\] net629 net609 _05264_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__o211a_1
XFILLER_166_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12310_ net1146 decoded_imm_j\[18\] net970 mem_rdata_q\[18\] VGND VGND VPWR VPWR
+ _06634_ sky130_fd_sc_hd__a22o_1
XFILLER_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13290_ net1020 net758 VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__or2_1
XFILLER_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08424__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout994_X net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12241_ net2717 net383 net372 net2734 VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_163_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12172_ net2879 net750 net368 VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06957__B1 net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11123_ net791 _05797_ _05799_ _05801_ net776 VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__o41a_1
XFILLER_96_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09255__S net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11054_ cpuregs\[17\]\[19\] net632 net610 _05734_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_178_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09371__A1 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10005_ net2857 _04770_ net1231 VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_125_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14813_ clknet_leaf_79_clk _01165_ VGND VGND VPWR VPWR decoded_imm\[9\] sky130_fd_sc_hd__dfxtp_2
XANTENNA_input19_X net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output122_A net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13505__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14744_ clknet_leaf_160_clk net2693 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11956_ net1046 net228 _02443_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__or3_2
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10907_ _05590_ _05591_ net809 VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__mux2_1
X_14675_ clknet_leaf_162_clk net2840 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11887_ _06355_ _06357_ _06291_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13626_ clknet_leaf_49_clk _00081_ VGND VGND VPWR VPWR cpuregs\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_10838_ net823 _05520_ _05522_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__a211o_1
XFILLER_158_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10769_ net1076 decoded_imm\[11\] net860 VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__o21a_1
X_13557_ net577 net2288 net411 VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__mux2_1
XFILLER_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12508_ _02395_ _05108_ net720 net866 VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__a31o_1
XFILLER_146_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13488_ net2255 net586 net422 VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__mux2_1
XFILLER_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15227_ clknet_leaf_32_clk _01568_ VGND VGND VPWR VPWR cpuregs\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12439_ net1157 _02507_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__nand2_1
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13391__C1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15158_ clknet_leaf_89_clk _01507_ VGND VGND VPWR VPWR mem_rdata_q\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06948__B1 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11695__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11941__B1 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14109_ clknet_leaf_199_clk _00563_ VGND VGND VPWR VPWR cpuregs\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15089_ clknet_leaf_19_clk _01441_ VGND VGND VPWR VPWR cpuregs\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_07980_ net968 _03309_ _03311_ net930 _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_52_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09165__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06931_ genblk2.pcpi_div.quotient\[0\] genblk2.pcpi_div.quotient\[1\] VGND VGND VPWR
+ VPWR _02515_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_26_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09650_ _03871_ reg_next_pc\[31\] net924 VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__mux2_1
X_06862_ net1089 net958 _02459_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08601_ _03969_ _03972_ _03974_ _03975_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__o211a_1
XFILLER_83_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09581_ count_instr\[60\] _04413_ count_instr\[61\] VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a21o_1
X_06793_ mem_rdata_q\[5\] VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__inv_2
X_08532_ genblk1.genblk1.pcpi_mul.rd\[8\] genblk1.genblk1.pcpi_mul.rdx\[8\] VGND VGND
+ VPWR VPWR _03918_ sky130_fd_sc_hd__nand2_1
XFILLER_24_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07413__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08463_ reg_pc\[28\] _03855_ reg_pc\[29\] VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07676__A1 net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14808__Q decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07414_ net1065 net1016 _02949_ net1079 _02948_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__a221o_1
X_08394_ _03803_ _03806_ net766 VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_34_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07428__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07345_ _02811_ _02884_ net1060 VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_63_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout320_A _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07428__B2 net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12555__A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _02357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13150__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
X_07276_ net1071 _02809_ _02810_ _02820_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__a31o_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09015_ net313 net2041 net518 VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__mux2_1
XANTENNA__07368__B decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold130 cpuregs\[12\]\[2\] VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 cpuregs\[24\]\[5\] VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _00966_ VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06939__B1 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold163 net37 VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11932__B1 net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold174 cpuregs\[8\]\[13\] VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A1 genblk2.pcpi_div.pcpi_rd\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold185 cpuregs\[12\]\[13\] VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 cpuregs\[30\]\[25\] VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net616 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09075__S net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout621 net622 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__buf_2
XANTENNA__11177__Y _05855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11618__B mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout632 net635 VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkbuf_4
X_09917_ net1127 _04445_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__xor2_1
Xfanout643 net644 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__clkbuf_2
Xfanout654 net679 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout954_A net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_8
Xfanout665 net672 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_2
Xfanout676 net679 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__clkbuf_2
X_09848_ _04630_ _04631_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__xnor2_1
Xfanout687 net696 VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__clkbuf_2
Xfanout698 net701 VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11160__A1 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout742_X net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09779_ _04545_ _04558_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11634__A net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11810_ genblk2.pcpi_div.divisor\[19\] genblk2.pcpi_div.dividend\[19\] VGND VGND
+ VPWR VPWR _06281_ sky130_fd_sc_hd__and2b_1
XANTENNA__07831__B net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ net1215 net2367 net2476 net906 net762 VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_103_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08419__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ net1462 net1171 net729 VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07667__A1 net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14460_ clknet_leaf_65_clk _00849_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11672_ is_lb_lh_lw_lbu_lhu _06228_ net547 VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__mux2_1
XFILLER_169_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10623_ _05297_ _05298_ _05315_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a21oi_2
X_13411_ net1002 net397 _02312_ _02317_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__o22a_1
X_14391_ clknet_leaf_86_clk _00812_ VGND VGND VPWR VPWR latched_stalu sky130_fd_sc_hd__dfxtp_1
XANTENNA__11215__A2 decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06890__A2 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12465__A net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13060__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13342_ net392 _02253_ _02254_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__or4_1
X_10554_ net801 _05245_ _05247_ net839 VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__a211o_1
XFILLER_139_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07278__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13273_ net1033 net752 VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10485_ cpuregs\[11\]\[1\] net633 net597 _05183_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__o211a_1
X_15012_ clknet_leaf_113_clk _01364_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_12224_ net750 _06604_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__nor2_1
XANTENNA__12715__A2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13296__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12155_ genblk2.pcpi_div.quotient_msk\[14\] net378 net367 net2785 VGND VGND VPWR
+ VPWR _01056_ sky130_fd_sc_hd__a22o_1
XANTENNA__12404__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10713__A net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11106_ net1082 _05784_ net859 VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12086_ net863 _06532_ _06533_ _06531_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__a31o_1
XFILLER_49_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_8
X_11037_ cpuregs\[2\]\[19\] net681 VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__or2_1
XFILLER_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13428__B1 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11544__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07107__B1 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08329__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09647__A2 net880 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12988_ net1425 net323 net448 VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__mux2_1
X_14727_ clknet_leaf_138_clk net2716 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11939_ net1189 _02507_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__and2_2
XANTENNA__07658__B2 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06866__C1 net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14658_ clknet_leaf_141_clk net2751 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ clknet_leaf_191_clk _00064_ VGND VGND VPWR VPWR cpuregs\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14589_ clknet_leaf_106_clk _00975_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10414__B1 _02507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07130_ genblk2.pcpi_div.dividend\[31\] _02684_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08083__A1 net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07061_ net1117 genblk2.pcpi_div.quotient\[20\] _02625_ net950 VGND VGND VPWR VPWR
+ _02627_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_41_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07188__B net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08999__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput202 net202 VGND VGND VPWR VPWR pcpi_insn[9] sky130_fd_sc_hd__buf_2
XFILLER_161_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput213 net1013 VGND VGND VPWR VPWR pcpi_rs1[19] sky130_fd_sc_hd__buf_2
Xoutput224 net995 VGND VGND VPWR VPWR pcpi_rs1[29] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR pcpi_rs2[0] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR pcpi_rs2[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_34_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput257 net257 VGND VGND VPWR VPWR pcpi_rs2[2] sky130_fd_sc_hd__buf_2
Xoutput268 net268 VGND VGND VPWR VPWR trap sky130_fd_sc_hd__buf_2
XFILLER_142_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10182__X _04888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06820__B net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07963_ net771 _03477_ _03478_ _03473_ VGND VGND VPWR VPWR alu_out\[2\] sky130_fd_sc_hd__a31o_1
XFILLER_114_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_79_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_8
X_06914_ net1084 is_sb_sh_sw _02483_ cpu_state\[6\] VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__a22o_1
X_09702_ _04496_ _04497_ _02481_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__a21oi_1
X_07894_ net1167 _02403_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__or2_1
XANTENNA__07346__B1 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06845_ mem_state\[0\] mem_state\[1\] VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__and2_1
X_09633_ reg_pc\[22\] net881 _04443_ net851 VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a22o_1
XANTENNA__12890__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13419__B1 net398 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13145__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11454__A net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09564_ _04404_ _04405_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__nor2_1
XANTENNA__08239__S net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06776_ net1053 VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__inv_2
XANTENNA__12269__B _04298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08515_ genblk1.genblk1.pcpi_mul.rd\[5\] genblk1.genblk1.pcpi_mul.next_rs2\[6\] net1096
+ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__nand3_1
XANTENNA__14538__Q is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07649__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09495_ count_instr\[29\] _04358_ count_instr\[30\] VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__a21o_1
XFILLER_24_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12984__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout535_A _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08446_ _03845_ _03848_ net769 VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__mux2_1
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08377_ reg_pc\[12\] _03788_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__xor2_1
XFILLER_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1065_X net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12716__C net1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07328_ net21 _02689_ _02694_ net4 _02812_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o221a_1
XFILLER_165_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11620__C mem_rdata_q\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10956__A1 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07259_ net1062 _02799_ _02804_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1232_X net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12572__X _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10270_ _04933_ _04975_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__or2_1
XANTENNA__10169__C1 net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10708__A1 net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout692_X net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12732__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11629__A mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07826__B net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout440 net442 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__buf_4
XANTENNA_fanout957_X net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout451 net452 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__buf_4
Xfanout462 _02118_ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_4
X_13960_ clknet_leaf_59_clk _00414_ VGND VGND VPWR VPWR cpuregs\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xfanout473 net474 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout484 _04288_ VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkbuf_8
Xfanout495 _04286_ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__buf_2
X_12911_ net341 net2139 net455 VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__mux2_1
XANTENNA__12881__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13891_ clknet_leaf_14_clk _00345_ VGND VGND VPWR VPWR cpuregs\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13055__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15630_ clknet_leaf_183_clk _01966_ VGND VGND VPWR VPWR cpuregs\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_61_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12842_ net355 net2157 net460 VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__mux2_1
XANTENNA__09629__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11436__A2 _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12633__A1 net1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15561_ clknet_leaf_19_clk _01897_ VGND VGND VPWR VPWR cpuregs\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12773_ net1220 net2540 net2573 net908 net764 VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__a221o_1
XFILLER_15_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12633__B2 net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14512_ clknet_leaf_78_clk _00901_ VGND VGND VPWR VPWR decoded_imm_j\[8\] sky130_fd_sc_hd__dfxtp_1
X_11724_ net96 net129 _06238_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__o21a_4
X_15492_ clknet_leaf_59_clk _01828_ VGND VGND VPWR VPWR cpuregs\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14443_ clknet_leaf_90_clk _00832_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ net1613 net2 net548 VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10606_ cpuregs\[22\]\[7\] cpuregs\[23\]\[7\] net668 VGND VGND VPWR VPWR _05299_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11586_ _02388_ mem_rdata_q\[13\] mem_rdata_q\[12\] VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__and3_1
X_14374_ clknet_leaf_136_clk _00795_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dfxtp_1
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13325_ net708 _02217_ _02239_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_70_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10537_ net830 _05227_ _05229_ _05231_ net790 VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_133_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13256_ net567 _05316_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__nor2_1
X_10468_ _03171_ _05142_ _05150_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a31oi_4
XFILLER_170_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11539__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12207_ genblk2.pcpi_div.quotient_msk\[17\] net269 net2735 VGND VGND VPWR VPWR _06596_
+ sky130_fd_sc_hd__a21oi_1
X_13187_ net1711 net318 net428 VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__mux2_1
X_10399_ net1165 net1166 _05102_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__or3_1
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12138_ net2989 _06577_ net274 VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__mux2_1
XFILLER_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12069_ _06518_ _06517_ _06515_ net861 VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09868__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07752__A net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12872__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10589__S net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10883__B1 net811 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08300_ reg_out\[27\] reg_next_pc\[27\] net925 VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__mux2_1
XFILLER_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09280_ net1869 net332 net484 VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__mux2_1
XFILLER_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08231_ net1056 net1170 net1162 net1055 VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__a22o_1
XANTENNA__09398__B net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10177__X _04883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08162_ _03292_ _03648_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__nor2_1
XFILLER_20_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07113_ genblk2.pcpi_div.quotient\[28\] _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__or2_1
XFILLER_107_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08093_ _03590_ _03591_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__nor2_1
XFILLER_118_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__clkinv_2
X_07044_ net1116 _02610_ genblk2.pcpi_div.quotient\[18\] VGND VGND VPWR VPWR _02612_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__09618__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload61 clknet_leaf_179_clk VGND VGND VPWR VPWR clkload61/X sky130_fd_sc_hd__clkbuf_4
Xclkload72 clknet_leaf_155_clk VGND VGND VPWR VPWR clkload72/Y sky130_fd_sc_hd__inv_8
Xclkload83 clknet_leaf_171_clk VGND VGND VPWR VPWR clkload83/X sky130_fd_sc_hd__clkbuf_8
XFILLER_115_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload94 clknet_leaf_145_clk VGND VGND VPWR VPWR clkload94/Y sky130_fd_sc_hd__clkinv_4
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11363__A1 net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12979__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08995_ net580 net1699 net518 VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_A _04288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07946_ is_compare net969 net935 net931 VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_3_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12312__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09353__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07877_ _03368_ _03394_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout273_X net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A net654 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09616_ _03800_ reg_next_pc\[14\] net920 VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__mux2_2
X_06828_ instr_or instr_ori VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__or2_1
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11615__C net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09547_ count_instr\[49\] count_instr\[48\] VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout440_X net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06759_ latched_is_lb VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__inv_2
XANTENNA__12615__B2 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_X net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09589__A net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09478_ count_instr\[24\] _04344_ _04348_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__and3_1
XFILLER_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08429_ _03833_ _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__nor2_1
XFILLER_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11440_ _06108_ _06109_ net817 VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__mux2_1
Xclkload0 clknet_4_0_0_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_22_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13040__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10929__A1 net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10247__B decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11371_ cpuregs\[14\]\[28\] cpuregs\[15\]\[28\] net689 VGND VGND VPWR VPWR _06043_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10322_ decoded_imm\[27\] net998 VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__nand2_1
X_13110_ net356 net2097 net435 VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14090_ clknet_leaf_52_clk _00544_ VGND VGND VPWR VPWR cpuregs\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08432__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13041_ net1345 net94 net535 VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__mux2_1
XFILLER_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13343__A2 net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10253_ decoded_imm\[4\] net1042 VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__or2_1
XFILLER_105_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10184_ net1188 _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__nand2b_1
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1202 net1203 VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__buf_2
Xfanout1213 net1222 VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__clkbuf_2
Xfanout1224 net34 VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1235 net1237 VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__buf_2
X_14992_ clknet_leaf_118_clk _01344_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11106__A1 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout270 net272 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout281 _03873_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_1
XANTENNA__09263__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout292 _03860_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_1
X_13943_ clknet_leaf_185_clk _00397_ VGND VGND VPWR VPWR cpuregs\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07291__B _02832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13874_ clknet_leaf_25_clk _00328_ VGND VGND VPWR VPWR cpuregs\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15613_ clknet_leaf_16_clk _01949_ VGND VGND VPWR VPWR cpuregs\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12825_ net293 net1979 net466 VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__mux2_1
XANTENNA__13513__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15544_ clknet_leaf_9_clk _01880_ VGND VGND VPWR VPWR cpuregs\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12756_ _02412_ net913 VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__nor2_1
XFILLER_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11707_ net2066 net310 net375 VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__mux2_1
X_15475_ clknet_leaf_3_clk _01811_ VGND VGND VPWR VPWR cpuregs\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12687_ net1200 genblk1.genblk1.pcpi_mul.next_rs2\[52\] net895 net2845 net712 VGND
+ VGND VPWR VPWR _01357_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14426_ clknet_leaf_67_clk alu_out\[26\] VGND VGND VPWR VPWR alu_out_q\[26\] sky130_fd_sc_hd__dfxtp_1
X_11638_ _06177_ _06198_ _06212_ _06221_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__or4_1
X_14357_ clknet_leaf_87_clk _00000_ VGND VGND VPWR VPWR decoder_trigger sky130_fd_sc_hd__dfxtp_1
X_11569_ net5 net4 _06166_ _06171_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__or4_1
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold707 cpuregs\[2\]\[10\] VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ reg_pc\[13\] net564 _02224_ net391 VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__a211o_1
Xhold718 cpuregs\[4\]\[4\] VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07747__A _02478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold729 cpuregs\[4\]\[10\] VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14288_ clknet_leaf_83_clk _00742_ VGND VGND VPWR VPWR count_cycle\[33\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10173__A net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13239_ _02403_ net753 VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__nand2_1
XFILLER_124_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08210__A1 net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12799__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07800_ _03316_ _03317_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__nor2_1
Xhold1407 genblk1.genblk1.pcpi_mul.rd\[61\] VGND VGND VPWR VPWR net2721 sky130_fd_sc_hd__dlygate4sd3_1
X_08780_ genblk1.genblk1.pcpi_mul.next_rs2\[47\] net1090 genblk1.genblk1.pcpi_mul.rd\[46\]
+ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1418 genblk2.pcpi_div.quotient_msk\[29\] VGND VGND VPWR VPWR net2732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 genblk2.pcpi_div.divisor\[27\] VGND VGND VPWR VPWR net2743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09173__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07731_ cpuregs\[24\]\[4\] net698 VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__or2_1
XFILLER_37_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07662_ _03181_ _03182_ net807 VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__mux2_1
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09401_ _04298_ net1113 net176 VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__nor3b_1
X_07593_ _03112_ _03113_ _03114_ _03100_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__a211o_1
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09332_ net1402 net585 net477 VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1303 VGND VGND VPWR VPWR picorv32_1303/HI trace_data[25] sky130_fd_sc_hd__conb_1
XFILLER_52_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpicorv32_1314 VGND VGND VPWR VPWR picorv32_1314/HI trace_valid sky130_fd_sc_hd__conb_1
XANTENNA__14816__Q decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09263_ net2191 net587 net486 VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08214_ _02383_ net1053 _02689_ net942 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__a22o_4
X_09194_ net284 net2054 net498 VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__mux2_1
X_08145_ _03464_ _03638_ _03639_ _03634_ VGND VGND VPWR VPWR alu_out\[23\] sky130_fd_sc_hd__a31o_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout400_A _04293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09348__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload150 clknet_leaf_110_clk VGND VGND VPWR VPWR clkload150/Y sky130_fd_sc_hd__inv_6
X_08076_ _03343_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__or2_1
XANTENNA__08252__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07252__A2 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload161 clknet_leaf_121_clk VGND VGND VPWR VPWR clkload161/Y sky130_fd_sc_hd__inv_8
Xclkload172 clknet_leaf_91_clk VGND VGND VPWR VPWR clkload172/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload183 clknet_leaf_105_clk VGND VGND VPWR VPWR clkload183/X sky130_fd_sc_hd__clkbuf_4
X_07027_ net1114 _02596_ genblk2.pcpi_div.dividend\[16\] VGND VGND VPWR VPWR _02597_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1028_X net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout390_X net390 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout867_A net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold12 genblk1.genblk1.pcpi_mul.next_rs1\[15\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13394__A net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold23 genblk1.genblk1.pcpi_mul.next_rs1\[18\] VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08978_ genblk1.genblk1.pcpi_mul.rd\[27\] genblk1.genblk1.pcpi_mul.rd\[59\] net956
+ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__mux2_1
Xhold34 net61 VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 cpuregs\[28\]\[4\] VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09083__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold56 genblk2.pcpi_div.instr_remu VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 cpuregs\[30\]\[24\] VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _03444_ _03446_ _03268_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__o21a_1
Xhold78 cpuregs\[22\]\[14\] VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold89 cpuregs\[26\]\[29\] VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10940_ cpuregs\[17\]\[16\] net621 net605 _05623_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__o211a_1
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ cpuregs\[16\]\[14\] net650 VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout822_X net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10957__S net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12738__A _02409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12610_ net1199 net2950 net893 net3022 _02054_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__a221o_1
X_13590_ net1321 VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13261__B2 net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12541_ genblk2.pcpi_div.divisor\[55\] _02027_ net874 VGND VGND VPWR VPWR _02028_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10258__A decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15260_ clknet_leaf_11_clk _01601_ VGND VGND VPWR VPWR cpuregs\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12472_ net1167 net715 _05101_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__or3b_1
XFILLER_138_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11024__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14211_ clknet_leaf_26_clk _00665_ VGND VGND VPWR VPWR reg_pc\[19\] sky130_fd_sc_hd__dfxtp_2
X_11423_ cpuregs\[27\]\[29\] net644 net602 _06093_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__o211a_1
XFILLER_126_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15191_ clknet_leaf_181_clk _01540_ VGND VGND VPWR VPWR cpuregs\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09258__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14142_ clknet_leaf_110_clk _00596_ VGND VGND VPWR VPWR count_instr\[13\] sky130_fd_sc_hd__dfxtp_1
X_11354_ cpuregs\[22\]\[27\] cpuregs\[23\]\[27\] net692 VGND VGND VPWR VPWR _06027_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13288__B _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10305_ _05008_ _05010_ _04911_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a21o_1
XFILLER_152_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11285_ cpuregs\[26\]\[25\] net704 VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__or2_1
X_14073_ clknet_leaf_190_clk _00527_ VGND VGND VPWR VPWR cpuregs\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10236_ decoded_imm\[6\] net1038 VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__or2_1
X_13024_ net317 net2391 net444 VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__mux2_1
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 net1011 VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 net209 VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13508__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07400__C1 _02935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10167_ count_cycle\[61\] _04873_ _04875_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__o21a_1
Xfanout1032 net234 VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12412__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1043 net229 VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__clkbuf_2
Xfanout1054 mem_wordsize\[2\] VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__buf_4
XFILLER_0_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10550__A2 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1065 net1070 VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1076 net1077 VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__clkbuf_2
Xfanout1087 cpu_state\[3\] VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14975_ clknet_leaf_116_clk _01327_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_10098_ count_cycle\[35\] count_cycle\[36\] count_cycle\[37\] _04826_ VGND VGND VPWR
+ VPWR _04831_ sky130_fd_sc_hd__and4_1
Xfanout1098 net1100 VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_145_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13926_ clknet_leaf_33_clk _00380_ VGND VGND VPWR VPWR cpuregs\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07703__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13857_ clknet_leaf_42_clk _00311_ VGND VGND VPWR VPWR cpuregs\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11552__A mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12808_ net403 net2148 net464 VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__mux2_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13252__A1 net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08337__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13788_ clknet_leaf_19_clk _00242_ VGND VGND VPWR VPWR cpuregs\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13252__B2 net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15527_ clknet_leaf_45_clk _01863_ VGND VGND VPWR VPWR cpuregs\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12739_ net1190 net1337 net2089 net883 _02103_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__a221o_1
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15458_ clknet_leaf_54_clk _01797_ VGND VGND VPWR VPWR cpuregs\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11698__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ clknet_leaf_170_clk alu_out\[9\] VGND VGND VPWR VPWR alu_out_q\[9\] sky130_fd_sc_hd__dfxtp_1
X_15389_ clknet_leaf_57_clk _01728_ VGND VGND VPWR VPWR cpuregs\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09168__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold504 cpuregs\[23\]\[27\] VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 cpuregs\[29\]\[29\] VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13198__B _05168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07234__A2 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold526 cpuregs\[21\]\[11\] VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 cpuregs\[29\]\[8\] VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14371__Q net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold548 instr_srai VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07196__B decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold559 cpuregs\[26\]\[0\] VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09950_ _04705_ _04708_ _04715_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_38_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12515__B1 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08901_ net1196 net2712 net890 _04227_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__a22o_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ net1127 _04442_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__and2_1
XFILLER_140_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11727__A net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08832_ genblk1.genblk1.pcpi_mul.next_rs2\[55\] net1103 genblk1.genblk1.pcpi_mul.rd\[54\]
+ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a21o_1
XFILLER_111_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1204 _01416_ VGND VGND VPWR VPWR net2518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 genblk2.pcpi_div.quotient_msk\[5\] VGND VGND VPWR VPWR net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 genblk1.genblk1.pcpi_mul.next_rs1\[41\] VGND VGND VPWR VPWR net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 genblk2.pcpi_div.divisor\[36\] VGND VGND VPWR VPWR net2551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _00600_ VGND VGND VPWR VPWR net2562 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ _04107_ _04110_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__nand2_1
Xhold1259 genblk1.genblk1.pcpi_mul.next_rs1\[42\] VGND VGND VPWR VPWR net2573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10829__B1 net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07714_ cpuregs\[5\]\[4\] net640 net819 _03232_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__o211a_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08694_ net899 _04053_ _04055_ net2622 net1202 VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__a32o_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07645_ cpuregs\[11\]\[2\] net640 net601 _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__o211a_1
XFILLER_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__06827__Y _02432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13153__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ reg_pc\[29\] decoded_imm\[29\] VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__and2_1
X_09315_ net1368 net332 net479 VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12992__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout615_A net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09246_ net1528 net336 net488 VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__mux2_1
XANTENNA__07473__A2 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13389__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09177_ net349 net1976 net497 VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1145_X net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11401__S net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09078__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08128_ _03319_ net932 VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__nand2_1
XANTENNA__12754__B1 net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07225__A2 _02767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08059_ _03379_ _03561_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__or2_1
Xoutput35 net35 VGND VGND VPWR VPWR mem_addr[10] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR mem_addr[21] sky130_fd_sc_hd__buf_2
Xoutput57 net57 VGND VGND VPWR VPWR mem_addr[31] sky130_fd_sc_hd__buf_2
X_11070_ net1159 net856 _05749_ _05750_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__a22o_1
Xoutput68 net68 VGND VGND VPWR VPWR mem_la_addr[12] sky130_fd_sc_hd__buf_2
Xoutput79 net79 VGND VGND VPWR VPWR mem_la_addr[23] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10517__C1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10021_ net2790 _04780_ net1223 VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11637__A mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09922__A1 net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07834__B net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11356__B net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ clknet_leaf_137_clk _00045_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11972_ net868 _06435_ _06436_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__and3_1
XFILLER_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_120_clk _00165_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10923_ cpuregs\[2\]\[16\] net659 VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__or2_1
X_14691_ clknet_leaf_141_clk _01076_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12690__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13063__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13642_ clknet_leaf_151_clk _00096_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10854_ net812 _05537_ _05539_ net823 VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__o211a_1
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09989__B2 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13573_ net324 net2494 net413 VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__mux2_1
X_10785_ cpuregs\[18\]\[12\] net552 _05472_ net779 VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__o22a_1
XFILLER_13_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15312_ clknet_leaf_194_clk _01652_ VGND VGND VPWR VPWR cpuregs\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09777__A decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12524_ genblk2.pcpi_div.divisor\[51\] net872 VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__nor2_1
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15243_ clknet_leaf_7_clk _01584_ VGND VGND VPWR VPWR cpuregs\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12455_ _06686_ net2545 net383 VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12407__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11311__S net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11406_ cpuregs\[1\]\[29\] net551 _06076_ net808 net837 VGND VGND VPWR VPWR _06077_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_169_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15174_ clknet_leaf_90_clk _01523_ VGND VGND VPWR VPWR mem_rdata_q\[25\] sky130_fd_sc_hd__dfxtp_2
X_12386_ net1487 net291 net363 VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__mux2_1
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14125_ clknet_leaf_50_clk _00579_ VGND VGND VPWR VPWR cpuregs\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_11337_ net805 _06009_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__or2_1
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output77_A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14056_ clknet_leaf_58_clk _00510_ VGND VGND VPWR VPWR cpuregs\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11268_ cpuregs\[10\]\[25\] net703 VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__or2_1
X_13007_ net572 net2220 net445 VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__mux2_1
XANTENNA__09913__A1 net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10219_ decoded_imm\[12\] net1026 net1024 decoded_imm\[13\] VGND VGND VPWR VPWR _04925_
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11199_ _05874_ _05875_ net821 VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_143_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14958_ clknet_leaf_144_clk net2951 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10287__A1 decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13909_ clknet_leaf_20_clk _00363_ VGND VGND VPWR VPWR cpuregs\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_14889_ clknet_leaf_105_clk _01241_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12681__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07152__B2 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07430_ net1074 _02956_ _02957_ _02964_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__a31o_1
XFILLER_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13225__A1 net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14366__Q net265 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11236__B1 net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07361_ net1140 count_cycle\[46\] net977 _02899_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__a211o_1
X_09100_ net1792 net539 net504 VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__mux2_1
X_07292_ reg_pc\[10\] decoded_imm\[10\] VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__xnor2_1
X_09031_ net571 net2254 net513 VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__mux2_1
XFILLER_163_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12736__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07207__A2 net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold301 cpuregs\[12\]\[15\] VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold312 genblk1.genblk1.pcpi_mul.pcpi_rd\[28\] VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 cpuregs\[22\]\[6\] VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold334 cpuregs\[29\]\[11\] VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 cpuregs\[24\]\[31\] VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 cpuregs\[12\]\[6\] VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__A2 net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold367 net40 VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 cpuregs\[28\]\[11\] VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09626__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09933_ _02480_ _04709_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__nand2_1
Xhold389 cpuregs\[23\]\[9\] VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 _03143_ VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__buf_2
XFILLER_131_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout814 net815 VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__clkbuf_4
Xfanout825 net826 VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13148__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09904__B2 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout836 net837 VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__clkbuf_4
Xfanout847 net852 VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__clkbuf_4
X_09864_ net1146 _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__nor2_1
Xfanout858 net859 VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1001 cpuregs\[18\]\[16\] VGND VGND VPWR VPWR net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 _05082_ VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1105_A net1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1012 cpuregs\[1\]\[0\] VGND VGND VPWR VPWR net2326 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _04151_ _04154_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__nand2_1
XFILLER_86_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1023 genblk1.genblk1.pcpi_mul.next_rs1\[32\] VGND VGND VPWR VPWR net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 cpuregs\[1\]\[29\] VGND VGND VPWR VPWR net2348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09795_ _04565_ _04574_ _04566_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12987__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1045 cpuregs\[17\]\[24\] VGND VGND VPWR VPWR net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 cpuregs\[18\]\[12\] VGND VGND VPWR VPWR net2370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07941__Y _03459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1067 cpuregs\[5\]\[24\] VGND VGND VPWR VPWR net2381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08746_ net887 _04097_ _04099_ net2598 net1197 VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__a32o_1
XANTENNA__12267__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1078 genblk1.genblk1.pcpi_mul.next_rs1\[23\] VGND VGND VPWR VPWR net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 cpuregs\[1\]\[15\] VGND VGND VPWR VPWR net2403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09361__S net478 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07679__C1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08677_ genblk1.genblk1.pcpi_mul.rd\[30\] genblk1.genblk1.pcpi_mul.next_rs2\[31\]
+ net1106 VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__nand3_1
XANTENNA__12672__C1 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07143__A1 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__B2 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ cpuregs\[1\]\[2\] net641 _03147_ net614 VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__o211a_1
XANTENNA__07694__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07559_ _03035_ _03046_ _03047_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_101_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10570_ cpuregs\[24\]\[6\] net677 VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__or2_1
XFILLER_166_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09229_ _03745_ _04277_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__nor2_4
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12240_ genblk2.pcpi_div.divisor\[3\] net383 net371 net2717 VGND VGND VPWR VPWR _01109_
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12171_ net2847 net380 net368 net2879 VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__a22o_1
XFILLER_150_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07845__A net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11122_ cpuregs\[11\]\[21\] net634 net591 _05800_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__o211a_1
XFILLER_123_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08440__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold890 cpuregs\[18\]\[15\] VGND VGND VPWR VPWR net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13058__S net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11053_ cpuregs\[16\]\[19\] net680 VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__or2_1
XFILLER_150_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10004_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] count_cycle\[3\] VGND
+ VGND VPWR VPWR _04771_ sky130_fd_sc_hd__and4_1
XFILLER_49_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12897__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07382__B2 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14812_ clknet_leaf_131_clk _01164_ VGND VGND VPWR VPWR decoded_imm\[10\] sky130_fd_sc_hd__dfxtp_2
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12258__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_945 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09271__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1590 instr_lw VGND VGND VPWR VPWR net2904 sky130_fd_sc_hd__dlygate4sd3_1
X_14743_ clknet_leaf_160_clk _01128_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11955_ genblk2.pcpi_div.dividend\[3\] _06422_ net277 VGND VGND VPWR VPWR _01012_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06908__B net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10906_ cpuregs\[20\]\[15\] cpuregs\[21\]\[15\] net646 VGND VGND VPWR VPWR _05591_
+ sky130_fd_sc_hd__mux2_1
X_14674_ clknet_leaf_162_clk _01059_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11886_ genblk2.pcpi_div.divisor\[14\] _02390_ _06292_ _06293_ _06356_ VGND VGND
+ VPWR VPWR _06357_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_15_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13625_ clknet_leaf_53_clk _00080_ VGND VGND VPWR VPWR cpuregs\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10837_ cpuregs\[18\]\[13\] net552 _05523_ net779 VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13521__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13556_ net581 net2212 net414 VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__mux2_1
X_10768_ net1076 _05456_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__nand2_1
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12507_ _05108_ net718 _02395_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10441__B2 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13487_ _04283_ _02127_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__nor2_1
X_10699_ cpuregs\[6\]\[10\] cpuregs\[7\]\[10\] net666 VGND VGND VPWR VPWR _05389_
+ sky130_fd_sc_hd__mux2_1
X_15226_ clknet_leaf_47_clk _01567_ VGND VGND VPWR VPWR cpuregs\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12438_ net1157 _02507_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__and2_1
XFILLER_126_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15157_ clknet_leaf_65_clk _01506_ VGND VGND VPWR VPWR mem_rdata_q\[8\] sky130_fd_sc_hd__dfxtp_1
X_12369_ net1849 net355 net360 VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__mux2_1
XANTENNA__11941__A1 net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14108_ clknet_leaf_195_clk _00562_ VGND VGND VPWR VPWR cpuregs\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07755__A net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15088_ clknet_leaf_179_clk _01440_ VGND VGND VPWR VPWR cpuregs\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14039_ clknet_leaf_184_clk _00493_ VGND VGND VPWR VPWR cpuregs\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_06930_ net953 _02510_ _02511_ _02514_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__o31ai_1
XANTENNA__11154__C1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09970__A net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06861_ _02451_ net958 mem_do_prefetch VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__and3b_1
XANTENNA__07373__A1 net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08600_ _03974_ _03975_ _03969_ _03972_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__a211o_1
X_09580_ count_instr\[60\] _04413_ _04415_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__o21a_1
X_06792_ mem_rdata_q\[2\] VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__inv_2
XANTENNA__12249__A2 net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12600__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09181__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08531_ net1195 net2883 net888 _03917_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__a22o_1
XFILLER_24_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06818__B instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08462_ reg_out\[29\] alu_out_q\[29\] net1155 VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__mux2_1
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07413_ genblk1.genblk1.pcpi_mul.pcpi_rd\[17\] genblk2.pcpi_div.pcpi_rd\[17\] net1111
+ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__mux2_1
X_08393_ _03804_ _03805_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__nor2_1
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07344_ net22 _02689_ _02694_ net5 _02812_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__o221a_1
XANTENNA__07428__A2 net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10968__C1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12555__B net716 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07275_ _02814_ _02819_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__or2_1
XANTENNA__12047__S net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1055_A mem_wordsize\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09014_ net318 net1665 net517 VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__mux2_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10790__S net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold120 cpuregs\[20\]\[3\] VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold131 cpuregs\[14\]\[21\] VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A _02378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold142 cpuregs\[20\]\[27\] VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 genblk1.genblk1.pcpi_mul.pcpi_rd\[1\] VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__S net478 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold164 cpuregs\[24\]\[6\] VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 cpuregs\[12\]\[3\] VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08260__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12290__B net739 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold186 cpuregs\[23\]\[21\] VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 cpuregs\[29\]\[21\] VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _03153_ VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkbuf_4
Xfanout611 net616 VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__clkbuf_2
Xfanout622 net624 VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__buf_2
X_09916_ net851 _04693_ _04694_ net881 net2487 VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1010_X net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout633 net635 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11618__C mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_2
XANTENNA__12488__A2 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_X net1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout655 net663 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkbuf_4
Xfanout666 net672 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkbuf_4
Xfanout677 net679 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__buf_2
X_09847_ decoded_imm_j\[17\] _04438_ _04621_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout470_X net470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout688 net691 VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout947_A net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07364__A1 net1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout699 net701 VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__buf_2
XANTENNA__07364__B2 net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_X net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09778_ _04565_ _04566_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_87_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09091__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ genblk1.genblk1.pcpi_mul.rd\[38\] genblk1.genblk1.pcpi_mul.next_rs2\[39\]
+ net1096 VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_103_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_X net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08313__B1 net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11126__S net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ net1575 net1173 net729 VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11671_ net29 net27 net28 _06226_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__nor4_1
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13410_ net394 _02313_ _02314_ _02316_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__or4_1
X_10622_ net773 _05306_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_157_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14390_ clknet_leaf_87_clk _00811_ VGND VGND VPWR VPWR latched_store sky130_fd_sc_hd__dfxtp_1
XANTENNA__08435__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10423__A1 net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13341_ net709 _02232_ _02255_ net565 reg_pc\[17\] VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__a32o_1
XFILLER_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10553_ cpuregs\[5\]\[6\] net629 net815 _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__o211a_1
XFILLER_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13272_ net567 _05386_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__nor2_1
XFILLER_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10484_ cpuregs\[10\]\[1\] net682 VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15011_ clknet_leaf_114_clk net2901 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_12223_ net2791 net273 net2820 VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09266__S net485 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13296__B _05491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12154_ net2859 net378 net366 net2863 VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__a22o_1
XANTENNA__11097__A net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11105_ net1081 decoded_imm\[20\] VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__or2_1
X_12085_ _06272_ _06521_ _06270_ _06271_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__a211o_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input31_X net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11036_ cpuregs\[1\]\[19\] net632 net610 _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__o211a_1
XANTENNA_output232_A net1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13516__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12420__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07514__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11544__B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12987_ net1567 net327 net449 VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__mux2_1
XFILLER_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14726_ clknet_leaf_138_clk _01111_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11938_ _06322_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__nor2_1
XANTENNA__07658__A2 net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10662__A1 net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14657_ clknet_leaf_143_clk net2603 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11869_ _06304_ _06339_ _06303_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_31_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13608_ clknet_leaf_195_clk _00063_ VGND VGND VPWR VPWR cpuregs\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14588_ clknet_leaf_104_clk _00974_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08345__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10414__A1 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13539_ net328 net1789 net415 VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__mux2_1
XANTENNA__10176__A net1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07060_ net1117 _02625_ net2761 VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput203 net203 VGND VGND VPWR VPWR pcpi_rs1[0] sky130_fd_sc_hd__buf_2
X_15209_ clknet_leaf_48_clk _01558_ VGND VGND VPWR VPWR cpuregs\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xoutput214 net1050 VGND VGND VPWR VPWR pcpi_rs1[1] sky130_fd_sc_hd__buf_2
Xoutput225 net225 VGND VGND VPWR VPWR pcpi_rs1[2] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VGND VGND VPWR VPWR pcpi_rs2[10] sky130_fd_sc_hd__buf_2
XANTENNA__09176__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput247 net247 VGND VGND VPWR VPWR pcpi_rs2[20] sky130_fd_sc_hd__buf_2
Xoutput258 net258 VGND VGND VPWR VPWR pcpi_rs2[30] sky130_fd_sc_hd__buf_2
XANTENNA__13116__A0 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07962_ _03278_ _03476_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__nand2_1
X_09701_ _04474_ _04484_ _04485_ _04483_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a31o_1
X_06913_ _02503_ _02504_ _02494_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__a21boi_1
XFILLER_96_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07893_ net1166 net1030 VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__and2b_1
XFILLER_55_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09632_ _03832_ reg_next_pc\[22\] net926 VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__mux2_2
X_06844_ mem_do_wdata mem_do_rdata mem_do_rinst VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__or3_1
XANTENNA__13419__B2 net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14819__Q decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09563_ net3034 _04403_ net1240 VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__o21ai_1
X_06775_ net1047 VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__inv_2
XFILLER_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08514_ genblk1.genblk1.pcpi_mul.rd\[5\] genblk1.genblk1.pcpi_mul.next_rs2\[6\] net1097
+ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_162_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09494_ net3047 _04358_ _04360_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07649__A2 decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08445_ _03846_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1172_A net1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13161__S net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout528_A _03746_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08376_ reg_out\[12\] alu_out_q\[12\] net1153 VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__mux2_1
XANTENNA__08255__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12285__B net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_177_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07327_ _02863_ _02865_ _02860_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__or3b_1
XFILLER_137_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07947__X _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10956__A2 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07258_ net1064 net1037 _02803_ net1078 _02802_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout897_A net898 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10373__X _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07189_ net26 net130 _02695_ net11 _02738_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09086__S net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11629__B mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07585__A1 genblk2.pcpi_div.pcpi_rd\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11118__C1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout430 _02129_ VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_4
XANTENNA__08003__B net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout441 net442 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_8
Xfanout452 net454 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__buf_4
Xfanout463 net464 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_X net852 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _06664_ VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_2
Xfanout485 _04288_ VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12910_ net346 net2347 net455 VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__mux2_1
Xfanout496 net497 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__buf_4
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13890_ clknet_leaf_15_clk _00344_ VGND VGND VPWR VPWR cpuregs\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12841_ net405 net2049 net460 VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__mux2_1
XFILLER_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15560_ clknet_leaf_31_clk _01896_ VGND VGND VPWR VPWR cpuregs\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12772_ net1220 net2289 net2540 net908 net764 VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__a221o_1
XANTENNA__08837__A1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14511_ clknet_leaf_80_clk _00900_ VGND VGND VPWR VPWR decoded_imm_j\[7\] sky130_fd_sc_hd__dfxtp_1
X_11723_ net1209 net268 VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__or2_1
XFILLER_159_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15491_ clknet_leaf_53_clk _01827_ VGND VGND VPWR VPWR cpuregs\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13071__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14442_ clknet_leaf_89_clk _00831_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11654_ net1406 net32 net548 VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__mux2_1
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10605_ _05285_ _05288_ _03171_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__o21a_1
X_14373_ clknet_leaf_171_clk _00794_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dfxtp_1
X_11585_ net2802 net562 _06189_ _06192_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__a22o_1
XFILLER_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13324_ net556 _02218_ _02240_ net564 reg_pc\[15\] VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__a32o_1
X_10536_ cpuregs\[27\]\[5\] net629 net595 _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__o211a_1
XFILLER_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13255_ net960 _02179_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12415__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10467_ _05165_ _05166_ net774 _05158_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__o211a_1
XFILLER_109_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12206_ net748 _06595_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__nor2_1
XANTENNA__11539__B net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13186_ net1720 net320 net428 VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__mux2_1
X_10398_ net1166 _05102_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__nor2_1
XFILLER_150_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12137_ net1189 net867 _06573_ _06576_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__a31o_1
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12068_ net1009 net722 _06516_ net861 VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__a31o_1
XANTENNA__07328__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12321__A1 decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07328__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11555__A is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11019_ net822 _05696_ _05698_ _05700_ net787 VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07752__B net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09025__A _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14709_ clknet_leaf_162_clk _01094_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_max_cap483_X net483 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07500__A1 net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08230_ net1056 net1171 net240 net942 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__a22o_2
XFILLER_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14374__Q net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08161_ _02396_ net1004 _03439_ net990 VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__a211o_1
XFILLER_118_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07112_ genblk2.pcpi_div.quotient\[27\] _02661_ net1123 VGND VGND VPWR VPWR _02670_
+ sky130_fd_sc_hd__o21a_1
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08092_ _03591_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__inv_2
X_07043_ net1116 genblk2.pcpi_div.quotient\[18\] _02610_ VGND VGND VPWR VPWR _02611_
+ sky130_fd_sc_hd__and3_1
Xclkload40 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload40/X sky130_fd_sc_hd__clkbuf_4
Xclkload51 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload51/X sky130_fd_sc_hd__clkbuf_4
Xclkload62 clknet_leaf_163_clk VGND VGND VPWR VPWR clkload62/X sky130_fd_sc_hd__clkbuf_8
Xclkload73 clknet_leaf_156_clk VGND VGND VPWR VPWR clkload73/Y sky130_fd_sc_hd__inv_8
XANTENNA__06831__B net975 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload84 clknet_leaf_173_clk VGND VGND VPWR VPWR clkload84/X sky130_fd_sc_hd__clkbuf_4
Xclkload95 clknet_leaf_146_clk VGND VGND VPWR VPWR clkload95/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_115_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07567__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11363__A2 _06034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08994_ net584 net1905 net518 VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__mux2_1
XANTENNA__10571__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_A net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09634__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07945_ instr_xor instr_xori VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout380_A net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13156__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12312__B2 mem_rdata_q\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07876_ net258 net992 VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nand2b_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09615_ reg_pc\[13\] net875 _04434_ net845 VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__a22o_1
XFILLER_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06827_ instr_or instr_ori VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__nor2_2
XANTENNA__12995__S net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10874__B2 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09546_ net1230 _04392_ _04393_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__and3_1
X_06758_ instr_bge VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__inv_2
XANTENNA__10626__A1 net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _02375_ _04347_ _04349_ net1215 VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__a211oi_1
XANTENNA_fanout812_A net821 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09589__B net1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout433_X net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_X net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08428_ reg_pc\[22\] _03829_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__and2_1
XFILLER_157_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_4_1_0_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_22_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08359_ reg_out\[9\] alu_out_q\[9\] net1153 VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout600_X net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11370_ net840 _06039_ _06041_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_115_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10321_ decoded_imm\[27\] net998 VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__and2_1
XFILLER_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13040_ net1333 net93 net535 VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12000__B1 net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10252_ _04949_ _04956_ _04957_ _04948_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__a211oi_2
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11927__X _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10183_ net1068 _02477_ _04883_ net393 VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__a31o_1
Xfanout1203 net1204 VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__buf_2
Xfanout1214 net1222 VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07853__A net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1225 net1227 VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__clkbuf_2
Xfanout1236 net1237 VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__buf_1
XANTENNA__08301__X net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14991_ clknet_leaf_118_clk net2895 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[38\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout271 net272 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13066__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11106__A2 _05784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12303__A1 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout282 net283 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_2
X_13942_ clknet_leaf_185_clk _00396_ VGND VGND VPWR VPWR cpuregs\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout293 _03857_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09180__A0 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13873_ clknet_leaf_176_clk _00327_ VGND VGND VPWR VPWR cpuregs\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15612_ clknet_leaf_45_clk _01948_ VGND VGND VPWR VPWR cpuregs\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12067__B1 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12824_ net297 net1842 net465 VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__mux2_1
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15543_ clknet_leaf_9_clk _01879_ VGND VGND VPWR VPWR cpuregs\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12755_ net1578 net899 _02111_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__a21o_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11706_ net2052 net314 net375 VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__mux2_1
X_15474_ clknet_leaf_194_clk _01810_ VGND VGND VPWR VPWR cpuregs\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12686_ net1195 net2845 net889 net3046 net712 VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__a221o_1
XFILLER_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14425_ clknet_leaf_83_clk alu_out\[25\] VGND VGND VPWR VPWR alu_out_q\[25\] sky130_fd_sc_hd__dfxtp_1
X_11637_ mem_rdata_q\[24\] mem_rdata_q\[7\] _06207_ _06220_ VGND VGND VPWR VPWR _06221_
+ sky130_fd_sc_hd__or4_1
XFILLER_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14356_ clknet_leaf_85_clk _00778_ VGND VGND VPWR VPWR mem_do_wdata sky130_fd_sc_hd__dfxtp_2
XFILLER_129_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11568_ net2994 net563 _06178_ _06185_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__a22o_1
XFILLER_156_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold708 cpuregs\[15\]\[31\] VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13307_ net556 _02204_ _02225_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__and3_1
Xhold719 cpuregs\[27\]\[11\] VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10519_ cpuregs\[1\]\[5\] net550 _05213_ net801 net829 VGND VGND VPWR VPWR _05214_
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14287_ clknet_leaf_84_clk _00741_ VGND VGND VPWR VPWR count_cycle\[32\] sky130_fd_sc_hd__dfxtp_1
X_11499_ pcpi_timeout_counter\[1\] pcpi_timeout_counter\[0\] _06160_ VGND VGND VPWR
+ VPWR _06161_ sky130_fd_sc_hd__nor3_1
XFILLER_170_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13238_ _04961_ _04968_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10173__B net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13169_ net1470 net575 net428 VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__mux2_1
XFILLER_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10553__B1 net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1408 genblk2.pcpi_div.divisor\[55\] VGND VGND VPWR VPWR net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 _01070_ VGND VGND VPWR VPWR net2733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07730_ _03247_ _03248_ net819 VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__mux2_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14369__Q net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07661_ cpuregs\[30\]\[2\] cpuregs\[31\]\[2\] net701 VGND VGND VPWR VPWR _03182_
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09400_ _04294_ _04295_ _04296_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__or4_4
XFILLER_81_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07592_ _03100_ _03114_ _03113_ _03112_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__o211a_1
X_09331_ net1537 net586 net477 VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1304 VGND VGND VPWR VPWR picorv32_1304/HI trace_data[26] sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09262_ _04277_ _04283_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__nor2_4
XFILLER_138_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08213_ _03698_ _03699_ _03693_ VGND VGND VPWR VPWR alu_out\[31\] sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_99_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09226__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09193_ net286 net2125 net499 VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__mux2_1
XFILLER_147_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07497__X _03027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08144_ _03327_ _03637_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__nand2_1
XANTENNA__06842__A net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload140 clknet_leaf_80_clk VGND VGND VPWR VPWR clkload140/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08075_ _03437_ _03576_ net989 VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__mux2_1
Xclkload151 clknet_leaf_111_clk VGND VGND VPWR VPWR clkload151/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout1135_A net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload162 clknet_leaf_122_clk VGND VGND VPWR VPWR clkload162/X sky130_fd_sc_hd__clkbuf_4
Xclkload173 clknet_leaf_92_clk VGND VGND VPWR VPWR clkload173/Y sky130_fd_sc_hd__inv_8
Xclkload184 clknet_leaf_106_clk VGND VGND VPWR VPWR clkload184/Y sky130_fd_sc_hd__inv_6
X_07026_ genblk2.pcpi_div.dividend\[15\] genblk2.pcpi_div.dividend\[14\] _02584_ VGND
+ VGND VPWR VPWR _02596_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_8_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout595_A net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07944__Y _03462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09364__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold13 _01385_ VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10370__Y _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08977_ net1629 _04265_ net945 VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__mux2_1
Xhold24 _01388_ VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold35 cpuregs\[24\]\[7\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold46 cpuregs\[22\]\[2\] VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold57 _00048_ VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _02397_ net998 _03380_ _03441_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__a221o_1
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold68 genblk1.genblk1.pcpi_mul.pcpi_rd\[27\] VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 genblk1.genblk1.pcpi_mul.pcpi_rd\[0\] VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10847__A1 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_X net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07859_ net240 net1022 VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__and2_1
X_10870_ _05554_ _05555_ net813 VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12738__B net912 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09529_ net2836 _04381_ net1227 VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout815_X net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11134__S net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12540_ net250 _02026_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10258__B net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12471_ _06698_ net2566 net386 VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__mux2_1
XFILLER_138_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14210_ clknet_leaf_27_clk _00664_ VGND VGND VPWR VPWR reg_pc\[18\] sky130_fd_sc_hd__dfxtp_2
X_11422_ cpuregs\[26\]\[29\] net707 VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__or2_1
XANTENNA__07848__A net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15190_ clknet_leaf_184_clk _01539_ VGND VGND VPWR VPWR cpuregs\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14141_ clknet_leaf_126_clk _00595_ VGND VGND VPWR VPWR count_instr\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11353_ cpuregs\[20\]\[27\] cpuregs\[21\]\[27\] net692 VGND VGND VPWR VPWR _06026_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10783__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10304_ _04912_ _04913_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_128_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14072_ clknet_leaf_186_clk _00526_ VGND VGND VPWR VPWR cpuregs\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11284_ cpuregs\[25\]\[25\] net644 net614 _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__o211a_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11327__A2 _05999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13023_ net322 net2194 net444 VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__mux2_1
X_10235_ decoded_imm\[6\] net1038 VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_167_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1000 net1001 VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09274__S net485 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1011 net215 VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__clkbuf_4
Xfanout1022 net1023 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__clkbuf_4
X_10166_ count_cycle\[61\] _04873_ net1209 VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__a21oi_1
Xfanout1033 net1034 VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__buf_2
Xfanout1044 net228 VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__buf_2
XANTENNA__07951__A1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1055 mem_wordsize\[2\] VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07951__B2 net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1066 net1070 VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1077 net1079 VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__buf_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1088 cpu_state\[2\] VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__buf_2
XFILLER_94_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14974_ clknet_leaf_118_clk _01326_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10097_ _04830_ net1225 _04829_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_128_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1099 net1100 VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_145_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10838__A1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13925_ clknet_leaf_23_clk _00379_ VGND VGND VPWR VPWR cpuregs\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkload4_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13524__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13856_ clknet_leaf_1_clk _00310_ VGND VGND VPWR VPWR cpuregs\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11552__B mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12807_ net409 net2026 net464 VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__mux2_1
XFILLER_50_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13787_ clknet_leaf_5_clk _00241_ VGND VGND VPWR VPWR cpuregs\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10999_ cpuregs\[2\]\[18\] cpuregs\[3\]\[18\] net648 VGND VGND VPWR VPWR _05681_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13252__A2 _05278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12738_ _02409_ net912 VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__nor2_1
X_15526_ clknet_leaf_39_clk _01862_ VGND VGND VPWR VPWR cpuregs\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15457_ clknet_leaf_59_clk _01796_ VGND VGND VPWR VPWR cpuregs\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07882__A_N net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12669_ net1203 net3071 net899 net2939 net713 VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__a221o_1
X_14408_ clknet_leaf_171_clk alu_out\[8\] VGND VGND VPWR VPWR alu_out_q\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07219__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07758__A net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08353__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15388_ clknet_leaf_36_clk _01727_ VGND VGND VPWR VPWR cpuregs\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_14339_ clknet_leaf_27_clk _06726_ VGND VGND VPWR VPWR reg_out\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold505 cpuregs\[2\]\[8\] VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 cpuregs\[23\]\[2\] VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold527 cpuregs\[29\]\[14\] VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 cpuregs\[20\]\[16\] VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 net202 VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08900_ _03958_ _03960_ _03957_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__a21bo_1
XFILLER_98_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12603__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ net851 _04660_ _04661_ net881 net2296 VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__a32o_1
XANTENNA__10526__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08195__A1 net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09184__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08831_ net900 _04169_ _04171_ net2884 net1203 VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__a32o_1
XFILLER_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1205 genblk1.genblk1.pcpi_mul.next_rs1\[52\] VGND VGND VPWR VPWR net2519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1216 _01046_ VGND VGND VPWR VPWR net2530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11219__S net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1227 genblk1.genblk1.pcpi_mul.next_rs1\[45\] VGND VGND VPWR VPWR net2541 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ _04111_ _04112_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nand2_1
Xhold1238 genblk2.pcpi_div.divisor\[33\] VGND VGND VPWR VPWR net2552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1249 genblk2.pcpi_div.divisor\[48\] VGND VGND VPWR VPWR net2563 sky130_fd_sc_hd__dlygate4sd3_1
X_07713_ cpuregs\[4\]\[4\] net698 VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__or2_1
XFILLER_39_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09695__A1 net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08693_ _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__inv_2
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07644_ cpuregs\[10\]\[2\] net699 VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__or2_1
XANTENNA__13228__C1 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06837__A net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07575_ reg_pc\[29\] decoded_imm\[29\] VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__nor2_1
XANTENNA__13243__A2 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09314_ net1435 net337 net479 VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__mux2_1
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09245_ net1667 net339 net488 VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__mux2_1
XANTENNA__07939__Y _03457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout510_A _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09359__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08263__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09176_ net353 net2187 net497 VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__mux2_1
XANTENNA__13389__B _05890_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12754__A1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08127_ _03464_ _03623_ _03618_ VGND VGND VPWR VPWR alu_out\[21\] sky130_fd_sc_hd__a21o_1
XANTENNA__12754__B2 net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1040_X net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1138_X net1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08058_ _03379_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout977_A net979 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput36 net36 VGND VGND VPWR VPWR mem_addr[11] sky130_fd_sc_hd__buf_2
XANTENNA_fanout598_X net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput47 net47 VGND VGND VPWR VPWR mem_addr[22] sky130_fd_sc_hd__buf_2
X_07009_ genblk2.pcpi_div.quotient\[12\] _02575_ net1118 VGND VGND VPWR VPWR _02582_
+ sky130_fd_sc_hd__o21a_1
Xoutput58 net58 VGND VGND VPWR VPWR mem_addr[3] sky130_fd_sc_hd__buf_2
Xoutput69 net69 VGND VGND VPWR VPWR mem_la_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_88_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09094__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10020_ count_cycle\[7\] count_cycle\[8\] count_cycle\[9\] _04776_ VGND VGND VPWR
+ VPWR _04781_ sky130_fd_sc_hd__and4_1
XFILLER_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11637__B mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10541__B net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1750 decoded_imm_j\[5\] VGND VGND VPWR VPWR net3064 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ net1039 net726 _06434_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout932_X net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13710_ clknet_leaf_120_clk _00164_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10922_ cpuregs\[1\]\[16\] net622 net605 _05605_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__o211a_1
X_14690_ clknet_leaf_142_clk _01075_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12690__B1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13641_ clknet_leaf_149_clk _00095_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10853_ net797 _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__or2_1
XANTENNA__13234__A2 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09989__A2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ net328 net2325 net411 VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__mux2_1
X_10784_ cpuregs\[19\]\[12\] net617 net589 VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__o21a_1
X_15311_ clknet_leaf_193_clk _01651_ VGND VGND VPWR VPWR cpuregs\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_13_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12523_ _05111_ net718 net245 VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09269__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15242_ clknet_leaf_7_clk _01583_ VGND VGND VPWR VPWR cpuregs\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12454_ _06684_ _06685_ genblk2.pcpi_div.divisor\[36\] net865 VGND VGND VPWR VPWR
+ _06686_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ cpuregs\[2\]\[29\] cpuregs\[3\]\[29\] net705 VGND VGND VPWR VPWR _06076_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15173_ clknet_leaf_91_clk _01522_ VGND VGND VPWR VPWR mem_rdata_q\[24\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_169_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12385_ net1457 net295 net363 VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__mux2_1
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14124_ clknet_leaf_54_clk _00578_ VGND VGND VPWR VPWR cpuregs\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11336_ cpuregs\[12\]\[27\] cpuregs\[13\]\[27\] net693 VGND VGND VPWR VPWR _06009_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13519__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14055_ clknet_leaf_60_clk _00509_ VGND VGND VPWR VPWR cpuregs\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11267_ cpuregs\[9\]\[25\] net643 net615 _05941_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__o211a_1
XANTENNA__12423__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10508__B1 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08177__A1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08177__B2 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13006_ net575 net2333 net444 VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__mux2_1
X_10218_ decoded_imm\[13\] net1024 VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__nand2_1
XANTENNA__11547__B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11198_ cpuregs\[4\]\[23\] cpuregs\[5\]\[23\] net675 VGND VGND VPWR VPWR _05875_
+ sky130_fd_sc_hd__mux2_1
X_10149_ count_cycle\[54\] count_cycle\[55\] _04860_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__and3_1
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_145_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14957_ clknet_leaf_121_clk _01309_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13908_ clknet_leaf_179_clk _00362_ VGND VGND VPWR VPWR cpuregs\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07688__B1 net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08348__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14888_ clknet_leaf_105_clk _01240_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07152__A2 net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13839_ clknet_leaf_45_clk _00293_ VGND VGND VPWR VPWR cpuregs\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10039__A2 _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07360_ count_instr\[46\] net1130 net1136 count_instr\[14\] VGND VGND VPWR VPWR _02899_
+ sky130_fd_sc_hd__a22o_1
X_15509_ clknet_leaf_167_clk _01845_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dfxtp_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07291_ _02834_ _02832_ _02827_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__or3b_1
XFILLER_164_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09179__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09030_ net576 net2485 net513 VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_154_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14382__Q net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12736__B2 net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10747__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold302 cpuregs\[31\]\[6\] VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09601__B2 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold313 cpuregs\[26\]\[10\] VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 cpuregs\[30\]\[29\] VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 instr_bltu VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 cpuregs\[22\]\[24\] VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 cpuregs\[13\]\[17\] VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold368 cpuregs\[10\]\[14\] VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _04705_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__xnor2_1
Xhold379 cpuregs\[14\]\[20\] VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08168__A1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout804 net806 VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08168__B2 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07427__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout815 net821 VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout826 _03137_ VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__buf_2
XFILLER_58_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _04623_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nor2_1
Xfanout837 _03137_ VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__buf_2
XANTENNA__09904__A2 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout848 net852 VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_A _03857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout859 _05134_ VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_163_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1002 cpuregs\[3\]\[5\] VGND VGND VPWR VPWR net2316 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ _04155_ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__nand2_1
XFILLER_97_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1013 cpuregs\[1\]\[1\] VGND VGND VPWR VPWR net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 _01402_ VGND VGND VPWR VPWR net2338 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09794_ _04580_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__and2_1
Xhold1035 net183 VGND VGND VPWR VPWR net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09642__S net925 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1046 cpuregs\[11\]\[23\] VGND VGND VPWR VPWR net2360 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _04098_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__inv_2
Xhold1057 cpuregs\[9\]\[22\] VGND VGND VPWR VPWR net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A _02118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1068 cpuregs\[5\]\[22\] VGND VGND VPWR VPWR net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 genblk1.genblk1.pcpi_mul.next_rs1\[51\] VGND VGND VPWR VPWR net2393 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12569__A net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13164__S net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_A _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07679__B1 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08676_ genblk1.genblk1.pcpi_mul.next_rs2\[31\] net1106 genblk1.genblk1.pcpi_mul.rd\[30\]
+ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__a21o_1
XANTENNA__08258__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12288__B net739 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07627_ net822 net796 VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_68_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout725_A _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ _03060_ _03073_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__or2_1
XFILLER_50_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout513_X net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07489_ reg_pc\[23\] decoded_imm\[23\] VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__nor2_1
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09089__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09228_ net1751 net280 net495 VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__mux2_1
XFILLER_166_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12727__B2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09159_ net1908 net291 net502 VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__mux2_1
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12170_ net2732 net380 net368 net2847 VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout882_X net882 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11121_ cpuregs\[10\]\[21\] net684 VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07845__B net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 cpuregs\[9\]\[20\] VGND VGND VPWR VPWR net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 cpuregs\[10\]\[5\] VGND VGND VPWR VPWR net2205 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08159__B2 net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11052_ _05731_ _05732_ net816 VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__mux2_1
XFILLER_89_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10003_ _04770_ net1231 _04769_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__and3b_1
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10910__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input21_A mem_rdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07382__A2 net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14811_ clknet_leaf_81_clk _01163_ VGND VGND VPWR VPWR decoded_imm\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13074__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1580 genblk1.genblk1.pcpi_mul.next_rs2\[37\] VGND VGND VPWR VPWR net2894 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_957 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14742_ clknet_leaf_160_clk _01127_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11954_ _06418_ _06419_ _06421_ net873 VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__a22o_1
Xhold1591 genblk1.genblk1.pcpi_mul.next_rs2\[53\] VGND VGND VPWR VPWR net2905 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12663__B1 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14467__Q instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10905_ cpuregs\[22\]\[15\] cpuregs\[23\]\[15\] net646 VGND VGND VPWR VPWR _05590_
+ sky130_fd_sc_hd__mux2_1
X_14673_ clknet_leaf_162_clk _01058_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11885_ _06296_ _06297_ _06351_ _06295_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_192_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_192_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output108_A net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13624_ clknet_leaf_73_clk _00079_ VGND VGND VPWR VPWR cpuregs\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_10836_ cpuregs\[19\]\[13\] net619 net590 VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_15_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13555_ net583 net2416 net413 VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__mux2_1
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10767_ net773 _05431_ _05439_ _05455_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__a31oi_4
XANTENNA__12418__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12506_ net2666 net387 _01999_ _02000_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__a22o_1
XANTENNA__10441__A2 net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13486_ net1559 net280 net425 VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__mux2_1
X_10698_ net1167 net853 _05387_ _05388_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__a22o_1
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15225_ clknet_leaf_37_clk _01566_ VGND VGND VPWR VPWR cpuregs\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12437_ _06672_ net2173 net384 VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__mux2_1
XFILLER_154_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13391__A1 net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15156_ clknet_leaf_65_clk _01505_ VGND VGND VPWR VPWR mem_rdata_q\[7\] sky130_fd_sc_hd__dfxtp_2
X_12368_ net1627 net405 net360 VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__mux2_1
XFILLER_153_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12661__B net913 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06948__A2 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14107_ clknet_leaf_195_clk _00561_ VGND VGND VPWR VPWR cpuregs\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11558__A mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11319_ _05991_ _05992_ net820 VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__mux2_1
XANTENNA__11941__A2 net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15087_ clknet_leaf_24_clk _01439_ VGND VGND VPWR VPWR cpuregs\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07755__B net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12299_ mem_rdata_q\[24\] net559 _06628_ net532 VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__a211o_1
XANTENNA__13143__A1 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14038_ clknet_leaf_185_clk _00492_ VGND VGND VPWR VPWR cpuregs\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07474__C _03005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06860_ net1060 cpu_state\[6\] VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__or2_1
XFILLER_110_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10901__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07771__A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06791_ net255 VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__inv_2
XFILLER_94_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08530_ _03915_ _03916_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07490__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14377__Q net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08461_ net289 net2531 net530 VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__mux2_1
XFILLER_24_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_183_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_183_clk sky130_fd_sc_hd__clkbuf_8
X_07412_ count_cycle\[17\] net974 net844 _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__o211a_1
XANTENNA__12406__A0 _03802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09698__A decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08392_ reg_pc\[15\] reg_pc\[14\] _03797_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_34_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07343_ _02880_ _02881_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__nand2_1
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07274_ net1064 net1034 _02818_ net1079 _02817_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__a221o_1
XANTENNA__10356__B net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09013_ net322 net2120 net517 VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__mux2_1
XFILLER_163_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12185__A2 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13382__A1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_A net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold110 genblk1.genblk1.pcpi_mul.pcpi_rd\[25\] VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold121 cpuregs\[24\]\[16\] VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold132 cpuregs\[26\]\[13\] VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11393__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold143 cpuregs\[26\]\[27\] VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 net146 VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13159__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12063__S net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold165 net159 VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 cpuregs\[22\]\[1\] VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold187 cpuregs\[21\]\[7\] VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _03153_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkbuf_4
Xhold198 net144 VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net616 VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09915_ net1184 _04444_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__or2_1
XANTENNA__12998__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout623 net624 VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkbuf_4
Xfanout634 net635 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_A net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout645 _03140_ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkbuf_4
Xfanout656 net663 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12893__A0 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout667 net672 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__clkbuf_2
X_09846_ _04628_ _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__nand2_1
XFILLER_98_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout678 net679 VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1003_X net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout689 net691 VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__buf_2
XANTENNA__09372__S net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07364__A2 net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ decoded_imm_j\[13\] _04434_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__nand2_1
X_06989_ _02563_ _02564_ net951 _02561_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout463_X net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout842_A _02702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08728_ genblk1.genblk1.pcpi_mul.next_rs2\[39\] net1096 genblk1.genblk1.pcpi_mul.rd\[38\]
+ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_87_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12645__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08659_ _04019_ _04022_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout630_X net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_174_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_174_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_120_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11670_ _06226_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__inv_2
XFILLER_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12746__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09401__A _04298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10621_ net827 _05309_ _05311_ _05313_ net789 VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__a2111o_1
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13340_ _02410_ net755 VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__nand2_1
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10552_ cpuregs\[4\]\[6\] net677 VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__or2_1
XFILLER_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13271_ _04974_ _04981_ _02193_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__a21oi_1
X_10483_ cpuregs\[9\]\[1\] net632 net610 _05181_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_118_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15010_ clknet_leaf_114_clk _01362_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_12222_ net749 net2726 VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__nor2_1
XFILLER_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07856__A net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08451__S net531 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13069__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12153_ net2803 net378 net366 net2859 VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__a22o_1
X_11104_ _05774_ _05783_ _05767_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__a21oi_4
X_12084_ _06270_ _06271_ _06272_ _06521_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__o211ai_1
XFILLER_150_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11136__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11665__X _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08001__B1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11035_ cpuregs\[0\]\[19\] net681 VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__or2_1
XANTENNA__12884__A0 mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07355__A2 decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09282__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input24_X net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output225_A net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11317__S net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12986_ net1346 net330 net447 VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__mux2_1
XANTENNA__12100__A2 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09501__B1 net1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14725_ clknet_leaf_141_clk _01110_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_165_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_165_clk sky130_fd_sc_hd__clkbuf_8
X_11937_ _06320_ _06321_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__nor2_1
XANTENNA__13532__S net416 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14656_ clknet_leaf_153_clk _01041_ VGND VGND VPWR VPWR genblk2.pcpi_div.running
+ sky130_fd_sc_hd__dfxtp_1
X_11868_ _06334_ _06338_ _06337_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__a21bo_1
X_10819_ cpuregs\[9\]\[13\] net619 net603 _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__o211a_1
X_13607_ clknet_leaf_2_clk _00062_ VGND VGND VPWR VPWR cpuregs\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14587_ clknet_leaf_114_clk net1877 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dfxtp_1
X_11799_ genblk2.pcpi_div.divisor\[23\] genblk2.pcpi_div.dividend\[23\] VGND VGND
+ VPWR VPWR _06270_ sky130_fd_sc_hd__and2b_1
XFILLER_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11052__S net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13538_ net332 net1709 net415 VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__mux2_1
XANTENNA__10176__B _02478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13469_ net1708 net345 net424 VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12167__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07766__A net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15208_ clknet_leaf_34_clk _01557_ VGND VGND VPWR VPWR cpuregs\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xoutput204 net204 VGND VGND VPWR VPWR pcpi_rs1[10] sky130_fd_sc_hd__buf_2
Xoutput215 net1011 VGND VGND VPWR VPWR pcpi_rs1[20] sky130_fd_sc_hd__buf_2
XANTENNA__08214__X net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput226 net993 VGND VGND VPWR VPWR pcpi_rs1[30] sky130_fd_sc_hd__buf_2
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11288__A net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput237 net237 VGND VGND VPWR VPWR pcpi_rs2[11] sky130_fd_sc_hd__buf_2
XANTENNA__08240__A0 net1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15139_ clknet_leaf_72_clk _01491_ VGND VGND VPWR VPWR cpuregs\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xoutput248 net248 VGND VGND VPWR VPWR pcpi_rs2[21] sky130_fd_sc_hd__buf_2
Xoutput259 net259 VGND VGND VPWR VPWR pcpi_rs2[31] sky130_fd_sc_hd__buf_2
XANTENNA__09981__A net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07961_ _03278_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__or2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09700_ _04493_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__nand2_1
X_06912_ net1088 net2671 VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__nand2_1
XANTENNA__12875__A0 mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07892_ _02394_ net1022 _03376_ _03409_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__a31o_1
XFILLER_68_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09192__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09631_ reg_pc\[21\] net881 _04442_ net851 VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a22o_1
X_06843_ _02441_ _00582_ _02446_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__or3b_1
XANTENNA__10886__C1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11227__S net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09562_ count_instr\[54\] _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__and2_1
X_06774_ net2852 VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__inv_2
XANTENNA__12627__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08513_ genblk1.genblk1.pcpi_mul.next_rs2\[6\] net1096 genblk1.genblk1.pcpi_mul.rd\[5\]
+ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__a21o_1
X_09493_ count_instr\[29\] _04358_ net1209 VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_156_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_156_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_64_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08444_ reg_pc\[25\] _03842_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08375_ net355 net2452 net529 VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout423_A net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout1165_A net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07326_ _02860_ _02864_ _02866_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__a21o_1
XFILLER_164_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10810__C1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07257_ genblk1.genblk1.pcpi_mul.pcpi_rd\[7\] genblk2.pcpi_div.pcpi_rd\[7\] net1110
+ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__mux2_1
XANTENNA__09367__S net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08271__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07188_ net1052 net1057 _02737_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout792_A net795 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08231__B1 net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11629__C mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10574__D1 net790 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout420 net422 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkbuf_4
Xfanout431 net432 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_4
XANTENNA__12866__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout442 _02125_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__buf_4
Xfanout453 net454 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__buf_4
Xfanout464 _02117_ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout475 net476 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__buf_4
Xfanout486 _04288_ VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09829_ net2569 net877 _04610_ _04614_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__a22o_1
Xfanout497 net499 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__buf_4
X_12840_ net409 net2240 net460 VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__mux2_1
XFILLER_100_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12771_ net1219 genblk1.genblk1.pcpi_mul.next_rs1\[39\] net2289 net908 net764 VGND
+ VGND VPWR VPWR _01410_ sky130_fd_sc_hd__a221o_1
XFILLER_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__B1 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_147_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_147_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11722_ net1208 net268 VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__nor2_1
X_14510_ clknet_leaf_80_clk _00899_ VGND VGND VPWR VPWR decoded_imm_j\[6\] sky130_fd_sc_hd__dfxtp_1
X_15490_ clknet_leaf_51_clk _01826_ VGND VGND VPWR VPWR cpuregs\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__06755__A net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14441_ clknet_leaf_64_clk _00830_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dfxtp_1
X_11653_ net1465 net31 net548 VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__mux2_1
X_10604_ net790 _05292_ _05294_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__or4_1
X_14372_ clknet_leaf_136_clk _00793_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dfxtp_4
X_11584_ net2281 net563 _06175_ _06192_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__a22o_1
X_13323_ net1022 net752 VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__or2_1
XFILLER_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10535_ cpuregs\[26\]\[5\] net678 VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__or2_1
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12492__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09277__S net485 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12149__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13254_ _04963_ _04965_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_133_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10466_ net834 _05161_ _05163_ net792 VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__a211o_1
X_12205_ net2776 net270 net2819 VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__a21oi_1
X_13185_ net2428 net324 net429 VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__mux2_1
XANTENNA__08222__B1 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10397_ net1167 _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__or2_1
XFILLER_124_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12136_ net864 _06574_ _06575_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__and3_1
XANTENNA__13527__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12067_ net722 _06516_ net1009 VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11018_ cpuregs\[27\]\[18\] net618 net589 _05699_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__o211a_1
XANTENNA__11555__B net1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08289__A0 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_138_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ net1785 net585 net449 VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__mux2_1
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14708_ clknet_leaf_162_clk _01093_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11290__B _05964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14639_ clknet_leaf_164_clk _01024_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08160_ _03272_ net931 _03652_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_60_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07111_ genblk2.pcpi_div.dividend\[28\] _02667_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__or2_1
X_08091_ net1161 net1018 _03344_ _03345_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__a31o_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10915__A net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11510__S net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload30 clknet_leaf_183_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__inv_8
XANTENNA__09187__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07042_ genblk2.pcpi_div.quotient\[17\] _02607_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__or2_1
Xclkload41 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload41/Y sky130_fd_sc_hd__clkinv_2
XFILLER_146_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11289__Y _05964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload52 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload52/X sky130_fd_sc_hd__clkbuf_8
Xclkload63 clknet_leaf_164_clk VGND VGND VPWR VPWR clkload63/X sky130_fd_sc_hd__clkbuf_8
Xclkload74 clknet_leaf_157_clk VGND VGND VPWR VPWR clkload74/Y sky130_fd_sc_hd__inv_12
XFILLER_115_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload85 clknet_leaf_174_clk VGND VGND VPWR VPWR clkload85/X sky130_fd_sc_hd__clkbuf_8
Xclkload96 clknet_leaf_147_clk VGND VGND VPWR VPWR clkload96/X sky130_fd_sc_hd__clkbuf_8
XFILLER_115_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07567__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12560__A2 net720 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08993_ net588 net1974 net518 VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__mux2_1
XFILLER_130_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07944_ instr_xor instr_xori VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_3_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__B1 net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07875_ net1157 net1188 VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__and2b_1
XANTENNA__11520__A0 mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_A net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06826_ instr_srl instr_srli instr_lbu instr_lb VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__or4_1
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09614_ _03795_ reg_next_pc\[13\] net920 VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__mux2_2
XANTENNA__10874__A2 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09650__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09545_ count_instr\[48\] _04391_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nand2_1
XANTENNA__12076__A1 net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06757_ instr_bgeu VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__inv_2
XFILLER_71_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_129_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_129_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_36_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13172__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11481__A net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09476_ _04344_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__and2_1
XANTENNA__10626__A2 net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08266__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08119__X alu_out\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08427_ reg_pc\[22\] _03829_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1070_X net1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_A net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1168_X net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08358_ net520 net2366 net529 VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__mux2_1
Xclkload2 clknet_4_2_0_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_22_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07309_ net991 _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__nor2_1
XFILLER_109_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08289_ net1009 _03728_ net982 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__mux2_2
XFILLER_137_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09097__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10320_ _04904_ _05024_ _04901_ _04903_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__o211a_1
XFILLER_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout795_X net795 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12000__A1 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10251_ decoded_imm\[3\] net1044 VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__nor2_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09952__B1 net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10182_ _02464_ _04882_ _04886_ _02459_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__or4bb_2
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1204 net1205 VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__clkbuf_2
Xfanout1215 net1216 VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__buf_2
Xfanout1226 net1227 VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__clkbuf_2
Xfanout1237 net1241 VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__buf_2
XANTENNA__07853__B net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10560__A net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14990_ clknet_leaf_119_clk _01342_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout272 _06403_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_2
XFILLER_115_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout283 _03870_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_2
X_13941_ clknet_leaf_188_clk _00395_ VGND VGND VPWR VPWR cpuregs\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xfanout294 _03857_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07715__C1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13872_ clknet_leaf_73_clk _00326_ VGND VGND VPWR VPWR cpuregs\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15611_ clknet_leaf_13_clk _01947_ VGND VGND VPWR VPWR cpuregs\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12823_ net301 net2086 net465 VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__mux2_1
XANTENNA__06756__Y _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12487__A net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13082__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15542_ clknet_leaf_10_clk _01878_ VGND VGND VPWR VPWR cpuregs\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12754_ net1214 genblk1.genblk1.pcpi_mul.next_rs1\[26\] net918 net999 VGND VGND VPWR
+ VPWR _02111_ sky130_fd_sc_hd__a22o_1
XFILLER_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11705_ net1906 net319 net374 VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__mux2_1
XANTENNA__07494__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15473_ clknet_leaf_192_clk _01809_ VGND VGND VPWR VPWR cpuregs\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12685_ net1197 genblk1.genblk1.pcpi_mul.next_rs2\[50\] net889 net2928 net711 VGND
+ VGND VPWR VPWR _01355_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_42_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ mem_rdata_q\[11\] mem_rdata_q\[10\] mem_rdata_q\[9\] mem_rdata_q\[8\] VGND
+ VGND VPWR VPWR _06220_ sky130_fd_sc_hd__or4_1
XFILLER_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14424_ clknet_leaf_83_clk alu_out\[24\] VGND VGND VPWR VPWR alu_out_q\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11567_ mem_rdata_q\[14\] mem_rdata_q\[13\] mem_rdata_q\[12\] VGND VGND VPWR VPWR
+ _06185_ sky130_fd_sc_hd__and3_1
X_14355_ clknet_leaf_85_clk _00777_ VGND VGND VPWR VPWR mem_do_rdata sky130_fd_sc_hd__dfxtp_2
XFILLER_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13306_ _02405_ net758 VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__nand2_1
X_10518_ cpuregs\[2\]\[5\] cpuregs\[3\]\[5\] net675 VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__mux2_1
X_14286_ clknet_leaf_97_clk _00740_ VGND VGND VPWR VPWR count_cycle\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold709 cpuregs\[5\]\[10\] VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ net2850 _06160_ _06157_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__o21bai_1
XFILLER_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13237_ net1042 net396 _02158_ _02164_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__o22a_1
X_10449_ net839 net816 _05148_ net792 VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_161_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08746__B2 net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13168_ net1526 net579 net429 VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__mux2_1
X_12119_ _06559_ _06560_ _06561_ net869 net275 VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13099_ net588 net2497 net437 VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1409 genblk1.genblk1.pcpi_mul.next_rs2\[9\] VGND VGND VPWR VPWR net2723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11285__B net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_176_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07660_ cpuregs\[28\]\[2\] cpuregs\[29\]\[2\] net701 VGND VGND VPWR VPWR _03181_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10856__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07591_ _03099_ _03101_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__and2b_1
XANTENNA__09459__C1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09330_ _04273_ _04281_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__nor2_2
XFILLER_80_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_1305 VGND VGND VPWR VPWR picorv32_1305/HI trace_data[27] sky130_fd_sc_hd__conb_1
XANTENNA__14385__Q net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09261_ net1768 net278 net490 VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__mux2_1
XANTENNA__07485__A1 genblk2.pcpi_div.pcpi_rd\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08212_ _03368_ _03697_ _03465_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_99_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09192_ net291 net1949 net498 VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08143_ _03327_ _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__or2_1
XFILLER_119_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload130 clknet_leaf_60_clk VGND VGND VPWR VPWR clkload130/Y sky130_fd_sc_hd__inv_8
X_08074_ _03374_ _03377_ _03574_ _03575_ _03375_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__o41a_1
Xclkload141 clknet_leaf_81_clk VGND VGND VPWR VPWR clkload141/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10792__A1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload152 clknet_leaf_112_clk VGND VGND VPWR VPWR clkload152/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload163 clknet_leaf_123_clk VGND VGND VPWR VPWR clkload163/Y sky130_fd_sc_hd__inv_8
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07025_ _02594_ _02595_ net950 _02592_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_77_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload174 clknet_leaf_94_clk VGND VGND VPWR VPWR clkload174/X sky130_fd_sc_hd__clkbuf_8
Xclkload185 clknet_leaf_107_clk VGND VGND VPWR VPWR clkload185/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_8_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1030_A net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1128_A decoded_imm_j\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout490_A _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10544__B2 net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout588_A _03749_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13167__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold14 genblk1.genblk1.pcpi_mul.next_rs1\[22\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ genblk1.genblk1.pcpi_mul.rd\[26\] genblk1.genblk1.pcpi_mul.rd\[58\] net957
+ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold25 genblk1.genblk1.pcpi_mul.next_rs1\[4\] VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 cpuregs\[24\]\[13\] VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold47 cpuregs\[20\]\[5\] VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _03291_ _03396_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__and2b_1
Xhold58 cpuregs\[26\]\[5\] VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12297__A1 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold69 cpuregs\[26\]\[15\] VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout755_A net757 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07858_ _03374_ _03375_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09380__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06809_ mem_do_rdata net983 VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__or2_1
X_07789_ _03303_ _03305_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout922_A net927 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09528_ count_instr\[42\] count_instr\[41\] count_instr\[40\] _04377_ VGND VGND VPWR
+ VPWR _04382_ sky130_fd_sc_hd__and4_1
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09459_ _02376_ _04335_ _04337_ net1206 VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__a211oi_1
XFILLER_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout710_X net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout808_X net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_49_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12470_ genblk2.pcpi_div.divisor\[40\] _06697_ net868 VGND VGND VPWR VPWR _06698_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11421_ cpuregs\[25\]\[29\] net644 net615 _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__o211a_1
XANTENNA__07848__B net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14140_ clknet_leaf_126_clk _00594_ VGND VGND VPWR VPWR count_instr\[11\] sky130_fd_sc_hd__dfxtp_1
X_11352_ net833 _06020_ _06022_ _06024_ net793 VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__a2111o_1
XFILLER_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10303_ _04913_ _05008_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__nand2_1
X_14071_ clknet_leaf_185_clk _00525_ VGND VGND VPWR VPWR cpuregs\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11283_ cpuregs\[24\]\[25\] net704 VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__or2_1
XFILLER_134_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13022_ net326 net2284 net445 VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__mux2_1
X_10234_ decoded_imm\[7\] net1035 VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__or2_1
XANTENNA__09925__B1 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11732__B1 _06243_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1001 net221 VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__buf_4
XANTENNA__13077__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1012 net1013 VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__buf_4
XANTENNA__07400__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10165_ _04873_ _04874_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__nor2_1
XFILLER_79_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07400__B2 net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1023 net208 VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 net233 VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__buf_2
XFILLER_0_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1045 net225 VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__buf_2
Xfanout1056 net1058 VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14973_ clknet_leaf_118_clk _01325_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_10096_ count_cycle\[35\] count_cycle\[36\] _04826_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__and3_1
Xfanout1067 net1070 VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1078 net1079 VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1089 cpu_state\[1\] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13924_ clknet_leaf_44_clk _00378_ VGND VGND VPWR VPWR cpuregs\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07703__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09290__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13855_ clknet_leaf_0_clk _00309_ VGND VGND VPWR VPWR cpuregs\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__06911__B1 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12806_ net521 net2083 net464 VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__mux2_1
XANTENNA__11552__C mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10998_ _05678_ _05679_ net809 VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__mux2_1
X_13786_ clknet_leaf_6_clk _00240_ VGND VGND VPWR VPWR cpuregs\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15525_ clknet_leaf_86_clk _01861_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07467__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12460__A1 net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12737_ net1337 net884 _02102_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__a21o_1
XANTENNA__13540__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15456_ clknet_leaf_53_clk _01795_ VGND VGND VPWR VPWR cpuregs\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12668_ net1210 net2939 net899 genblk1.genblk1.pcpi_mul.next_rs2\[32\] net713 VGND
+ VGND VPWR VPWR _01338_ sky130_fd_sc_hd__a221o_1
XFILLER_129_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14407_ clknet_leaf_136_clk alu_out\[7\] VGND VGND VPWR VPWR alu_out_q\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07219__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11619_ mem_rdata_q\[4\] mem_rdata_q\[6\] VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__nand2_1
XANTENNA__07758__B net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07219__B2 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15387_ clknet_leaf_16_clk _01726_ VGND VGND VPWR VPWR cpuregs\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11060__S net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12599_ net297 net2397 net469 VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__mux2_1
XFILLER_129_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14338_ clknet_leaf_27_clk _06725_ VGND VGND VPWR VPWR reg_out\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold506 cpuregs\[29\]\[25\] VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 genblk1.genblk1.pcpi_mul.pcpi_rd\[8\] VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold528 cpuregs\[6\]\[26\] VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold539 cpuregs\[27\]\[3\] VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ clknet_leaf_129_clk _00723_ VGND VGND VPWR VPWR count_cycle\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09916__B1 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07774__A net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__inv_2
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1206 genblk1.genblk1.pcpi_mul.next_rs1\[8\] VGND VGND VPWR VPWR net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 cpuregs\[18\]\[28\] VGND VGND VPWR VPWR net2531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08761_ genblk1.genblk1.pcpi_mul.next_rs2\[44\] net1091 genblk1.genblk1.pcpi_mul.rd\[43\]
+ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a21o_1
Xhold1228 pcpi_timeout_counter\[3\] VGND VGND VPWR VPWR net2542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 genblk2.pcpi_div.divisor\[58\] VGND VGND VPWR VPWR net2553 sky130_fd_sc_hd__dlygate4sd3_1
X_07712_ cpuregs\[6\]\[4\] cpuregs\[7\]\[4\] net698 VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__mux2_1
XANTENNA__10829__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08692_ genblk1.genblk1.pcpi_mul.next_rs2\[33\] net1101 _04050_ _04052_ VGND VGND
+ VPWR VPWR _04054_ sky130_fd_sc_hd__and4_1
XFILLER_65_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07643_ cpuregs\[9\]\[2\] net640 net614 _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__o211a_1
XANTENNA__11239__C1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07574_ net1072 _03090_ _03091_ _03098_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_24_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09313_ net1754 net339 net479 VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__mux2_1
XANTENNA__07458__A1 net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09852__C1 net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
X_09244_ net1392 net343 net489 VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1078_A net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09175_ net356 net2140 net496 VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__mux2_1
XFILLER_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08126_ _03334_ _03622_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11411__C1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08057_ _03436_ _03560_ net988 VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__mux2_1
XANTENNA__07630__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1033_X net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07008_ net947 _02579_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__or3_1
XANTENNA__09375__S net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput37 net37 VGND VGND VPWR VPWR mem_addr[12] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VGND VGND VPWR VPWR mem_addr[23] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_X net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10517__A1 net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput59 net59 VGND VGND VPWR VPWR mem_addr[4] sky130_fd_sc_hd__buf_2
XANTENNA_fanout872_A net873 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08959_ net2091 _04256_ net944 VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__mux2_1
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11934__A net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1740 count_cycle\[10\] VGND VGND VPWR VPWR net3054 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1751 count_instr\[12\] VGND VGND VPWR VPWR net3065 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ net726 _06434_ net1039 VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__a21o_1
XFILLER_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07697__A1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10921_ cpuregs\[0\]\[16\] net658 VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__or2_1
XANTENNA__13219__B1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_X net925 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11574__C_N mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10852_ cpuregs\[12\]\[14\] cpuregs\[13\]\[14\] net651 VGND VGND VPWR VPWR _05538_
+ sky130_fd_sc_hd__mux2_1
X_13640_ clknet_leaf_148_clk _00094_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13571_ net332 net2228 net411 VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__mux2_1
XANTENNA__10984__S net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10783_ cpuregs\[17\]\[12\] net617 net603 _05470_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_51_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
X_15310_ clknet_leaf_181_clk _01650_ VGND VGND VPWR VPWR cpuregs\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07859__A net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12522_ net1159 net716 _05111_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__or3b_1
XANTENNA__08307__X net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15241_ clknet_leaf_18_clk _01582_ VGND VGND VPWR VPWR cpuregs\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12453_ net1174 _05098_ net717 net865 VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__a31o_1
XFILLER_166_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12745__A2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11404_ net808 _06072_ _06074_ net839 VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__a211o_1
X_15172_ clknet_leaf_90_clk _01521_ VGND VGND VPWR VPWR mem_rdata_q\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_166_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12384_ net1571 net300 net362 VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10756__A1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14123_ clknet_leaf_66_clk _00577_ VGND VGND VPWR VPWR cpuregs\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_11335_ cpuregs\[14\]\[27\] cpuregs\[15\]\[27\] net693 VGND VGND VPWR VPWR _06008_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07621__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09285__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11266_ cpuregs\[8\]\[25\] net703 VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__or2_1
X_14054_ clknet_leaf_37_clk _00508_ VGND VGND VPWR VPWR cpuregs\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output255_A net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10732__B decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10217_ _04917_ _04920_ _04921_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__and3_1
X_13005_ net580 net2344 net445 VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__mux2_1
XANTENNA__11547__C net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12005__A net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11197_ cpuregs\[6\]\[23\] cpuregs\[7\]\[23\] net675 VGND VGND VPWR VPWR _05874_
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10148_ count_cycle\[54\] _04860_ count_cycle\[55\] VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13535__S net416 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ count_cycle\[29\] _04816_ count_cycle\[30\] VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_50_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14956_ clknet_leaf_120_clk _01308_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13907_ clknet_leaf_23_clk _00361_ VGND VGND VPWR VPWR cpuregs\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14887_ clknet_leaf_104_clk _01239_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13838_ clknet_leaf_36_clk _00292_ VGND VGND VPWR VPWR cpuregs\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11236__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13769_ clknet_leaf_52_clk _00223_ VGND VGND VPWR VPWR cpuregs\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_42_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15508_ clknet_leaf_173_clk _01844_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07769__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08364__S net529 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07290_ net1063 net1031 _02833_ net1077 _02829_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__a221o_1
XFILLER_149_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10995__A1 net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15439_ clknet_leaf_194_clk _01778_ VGND VGND VPWR VPWR cpuregs\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09984__A net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09601__A2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold303 cpuregs\[28\]\[6\] VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 cpuregs\[10\]\[15\] VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 cpuregs\[10\]\[10\] VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold336 cpuregs\[21\]\[5\] VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold347 cpuregs\[16\]\[3\] VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 cpuregs\[30\]\[27\] VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 cpuregs\[31\]\[12\] VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _04706_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__nor2_1
Xfanout805 net806 VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__buf_4
Xfanout816 net818 VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__clkbuf_4
Xfanout827 net828 VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _04439_ _04440_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nand2_1
Xfanout838 net839 VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__buf_4
Xfanout849 net850 VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__buf_2
XANTENNA__10904__D1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07376__B1 _02387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1003 cpuregs\[9\]\[9\] VGND VGND VPWR VPWR net2317 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ genblk1.genblk1.pcpi_mul.next_rs2\[52\] net1099 genblk1.genblk1.pcpi_mul.rd\[51\]
+ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__a21o_1
XANTENNA__13449__B1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09793_ decoded_imm_j\[14\] _04435_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__nand2_1
Xhold1014 cpuregs\[9\]\[0\] VGND VGND VPWR VPWR net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1025 cpuregs\[19\]\[12\] VGND VGND VPWR VPWR net2339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 cpuregs\[5\]\[1\] VGND VGND VPWR VPWR net2350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 cpuregs\[25\]\[31\] VGND VGND VPWR VPWR net2361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1058 cpuregs\[17\]\[27\] VGND VGND VPWR VPWR net2372 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ genblk1.genblk1.pcpi_mul.next_rs2\[41\] net1092 _04094_ _04096_ VGND VGND
+ VPWR VPWR _04098_ sky130_fd_sc_hd__and4_1
Xhold1069 cpuregs\[19\]\[28\] VGND VGND VPWR VPWR net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08675_ net904 _04037_ _04039_ net2789 net1217 VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__a32o_1
XANTENNA__07679__A1 net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11475__A2 _06143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_A net454 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10683__B1 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ cpuregs\[0\]\[2\] net700 VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07557_ net1072 _03074_ _03075_ _03082_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout620_A net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13180__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A net720 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08274__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07488_ net1073 _03010_ _03011_ _03018_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__a31o_1
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08127__X alu_out\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09227_ net1674 net284 net495 VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1150_X net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_X net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09158_ net2098 net295 net503 VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__mux2_1
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08109_ _03329_ _03606_ net933 _03328_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09089_ net1608 net289 net510 VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__mux2_1
XFILLER_163_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11120_ cpuregs\[9\]\[21\] net623 net606 _05798_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__o211a_1
XFILLER_150_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold870 cpuregs\[3\]\[2\] VGND VGND VPWR VPWR net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 cpuregs\[8\]\[25\] VGND VGND VPWR VPWR net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ cpuregs\[20\]\[19\] cpuregs\[21\]\[19\] net680 VGND VGND VPWR VPWR _05732_
+ sky130_fd_sc_hd__mux2_1
Xhold892 cpuregs\[18\]\[2\] VGND VGND VPWR VPWR net2206 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10002_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] VGND VGND VPWR VPWR _04770_
+ sky130_fd_sc_hd__and3_1
XFILLER_89_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ clknet_leaf_77_clk _01162_ VGND VGND VPWR VPWR decoded_imm\[12\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_125_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07119__B1 net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1570 genblk1.genblk1.pcpi_mul.rd\[53\] VGND VGND VPWR VPWR net2884 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input14_A mem_rdata[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14741_ clknet_leaf_160_clk _01126_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[20\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1581 _01343_ VGND VGND VPWR VPWR net2895 sky130_fd_sc_hd__dlygate4sd3_1
X_11953_ _02402_ _06420_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__xnor2_1
Xhold1592 count_cycle\[1\] VGND VGND VPWR VPWR net2906 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12663__B2 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10904_ net822 _05584_ _05586_ _05588_ net787 VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10674__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14672_ clknet_leaf_162_clk net2777 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11884_ _06332_ _06354_ _06343_ _06353_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__o2bb2a_1
X_13623_ clknet_leaf_46_clk _00078_ VGND VGND VPWR VPWR cpuregs\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_10835_ cpuregs\[17\]\[13\] net619 net604 _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_15_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09816__C1 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13090__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13554_ net587 net2526 net413 VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__mux2_1
X_10766_ net780 _05445_ _05454_ net777 VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__o211a_1
XFILLER_41_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12505_ net870 _01997_ _01998_ net387 VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__a31oi_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13485_ net1610 net282 net425 VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__mux2_1
X_10697_ net1076 _05386_ net853 VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__a21oi_1
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09044__A0 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13376__C1 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15224_ clknet_leaf_79_clk _01565_ VGND VGND VPWR VPWR reg_sh\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12436_ net1180 genblk2.pcpi_div.divisor\[32\] net865 VGND VGND VPWR VPWR _06672_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10729__B2 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15155_ clknet_leaf_89_clk _01504_ VGND VGND VPWR VPWR mem_rdata_q\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13391__A2 net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12367_ net1362 net409 net360 VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__mux2_1
XFILLER_141_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output82_A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14106_ clknet_leaf_196_clk _00560_ VGND VGND VPWR VPWR cpuregs\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11318_ cpuregs\[20\]\[26\] cpuregs\[21\]\[26\] net702 VGND VGND VPWR VPWR _05992_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11941__A3 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15086_ clknet_leaf_29_clk _01438_ VGND VGND VPWR VPWR cpuregs\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12298_ decoded_imm\[24\] net733 VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14037_ clknet_leaf_187_clk _00491_ VGND VGND VPWR VPWR cpuregs\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11249_ net792 _05920_ _05922_ _05924_ net778 VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__o41a_1
XANTENNA__11154__A1 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10889__S net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11574__A mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07771__B net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06790_ net256 VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__inv_2
XANTENNA__08359__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14939_ clknet_leaf_18_clk _01291_ VGND VGND VPWR VPWR cpuregs\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08460_ _03858_ _03859_ net768 VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__mux2_2
XFILLER_63_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07411_ count_instr\[17\] net1136 net977 _02946_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__a211o_1
XFILLER_90_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08391_ reg_pc\[14\] _03797_ reg_pc\[15\] VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_15_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11513__S net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07342_ _02880_ _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__or2_1
XFILLER_148_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10968__A1 net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07273_ genblk1.genblk1.pcpi_mul.pcpi_rd\[8\] genblk2.pcpi_div.pcpi_rd\[8\] net1110
+ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__mux2_1
XANTENNA__11090__B1 net811 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09012_ net326 net2275 net518 VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__mux2_1
XFILLER_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 instr_auipc VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 cpuregs\[30\]\[20\] VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__B net969 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold122 genblk1.genblk1.pcpi_mul.pcpi_rd\[2\] VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold133 net136 VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 cpuregs\[12\]\[30\] VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07438__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 cpuregs\[22\]\[9\] VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 cpuregs\[30\]\[13\] VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold177 genblk1.genblk1.pcpi_mul.next_rs1\[2\] VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07895__A_N net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold188 cpuregs\[21\]\[20\] VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold199 cpuregs\[22\]\[29\] VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 _03153_ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__buf_2
X_09914_ net984 _04689_ _04692_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__o21ai_1
Xfanout613 net616 VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1110_A net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout624 net645 VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkbuf_2
Xfanout635 net645 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1208_A net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout646 net649 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_A mem_rdata[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout657 net663 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__clkbuf_4
X_09845_ decoded_imm_j\[18\] _04439_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__or2_1
XANTENNA__12893__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout668 net672 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__buf_2
Xfanout679 _03139_ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13175__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08269__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09776_ decoded_imm_j\[13\] _04434_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__nor2_1
XFILLER_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06988_ net1120 genblk2.pcpi_div.quotient\[10\] _02562_ net951 VGND VGND VPWR VPWR
+ _02564_ sky130_fd_sc_hd__a31o_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ net892 _04081_ _04083_ net2869 net1201 VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_87_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_X net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12645__B2 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_X net1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08658_ _04023_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07609_ count_cycle\[31\] net973 net843 _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout623_X net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08589_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__inv_2
XANTENNA__09401__B net1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10620_ cpuregs\[27\]\[7\] net626 net594 _05312_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__o211a_1
XFILLER_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07202__A net1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_22_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10551_ cpuregs\[6\]\[6\] cpuregs\[7\]\[6\] net677 VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__mux2_1
X_13270_ _04974_ _04981_ net959 VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__o21ai_1
X_10482_ cpuregs\[8\]\[1\] net682 VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout992_X net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12221_ genblk2.pcpi_div.quotient_msk\[24\] net273 net2725 VGND VGND VPWR VPWR _06603_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07856__B net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09129__A _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ genblk2.pcpi_div.quotient_msk\[11\] net379 net367 net2803 VGND VGND VPWR
+ VPWR _01053_ sky130_fd_sc_hd__a22o_1
XFILLER_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11103_ net788 _05778_ _05780_ _05782_ net776 VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__o41a_1
X_12083_ _06529_ _06530_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__nor2_1
XFILLER_123_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11034_ _05713_ _05714_ net816 VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__mux2_1
XANTENNA__12884__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13085__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10895__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08179__S net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input17_X net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12985_ net1812 net333 net447 VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__mux2_1
XANTENNA_output218_A net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10647__B1 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14724_ clknet_leaf_141_clk net2718 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11936_ genblk2.pcpi_div.dividend\[0\] _06406_ net276 VGND VGND VPWR VPWR _01009_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07512__B1 net979 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11617__B_N mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14655_ clknet_leaf_150_clk _01040_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11867_ _06305_ _06306_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__nor2_1
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13606_ clknet_leaf_191_clk _00061_ VGND VGND VPWR VPWR cpuregs\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13061__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10818_ cpuregs\[8\]\[13\] net652 VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__or2_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14586_ clknet_leaf_115_clk _00972_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11798_ _06267_ _06268_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13537_ net336 net1752 net415 VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__mux2_1
X_10749_ cpuregs\[18\]\[11\] net553 _05437_ net780 VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__o22a_1
X_13468_ net1429 net348 net423 VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11569__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15207_ clknet_leaf_33_clk _01556_ VGND VGND VPWR VPWR cpuregs\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07766__B net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12419_ net293 net2039 net473 VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__mux2_1
Xoutput205 net205 VGND VGND VPWR VPWR pcpi_rs1[11] sky130_fd_sc_hd__buf_2
XFILLER_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13399_ _02412_ net756 VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__nand2_1
XFILLER_154_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput216 net1009 VGND VGND VPWR VPWR pcpi_rs1[21] sky130_fd_sc_hd__buf_2
Xoutput227 net1189 VGND VGND VPWR VPWR pcpi_rs1[31] sky130_fd_sc_hd__buf_2
Xoutput238 net238 VGND VGND VPWR VPWR pcpi_rs2[12] sky130_fd_sc_hd__buf_2
X_15138_ clknet_leaf_31_clk _01490_ VGND VGND VPWR VPWR cpuregs\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08240__A1 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput249 net249 VGND VGND VPWR VPWR pcpi_rs2[22] sky130_fd_sc_hd__buf_2
XFILLER_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10192__B net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15069_ clknet_leaf_103_clk _01421_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_07960_ _03423_ _03475_ net989 VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__mux2_1
XFILLER_142_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12324__B1 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07782__A net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06911_ net1084 is_sll_srl_sra _02477_ net1068 VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08230__X net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12875__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07891_ net1162 net1020 VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__and2b_1
XFILLER_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11508__S net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09630_ _03827_ reg_next_pc\[21\] net926 VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__mux2_2
X_06842_ net1208 _02445_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__or2_1
XANTENNA__14388__Q net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09561_ _02372_ _04401_ _04403_ net1216 VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__a211oi_1
X_06773_ net1150 VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__inv_2
XANTENNA__12627__B2 net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10638__B1 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08512_ net893 _03899_ _03901_ net2604 net1200 VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__a32o_1
X_09492_ _04358_ _04359_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07721__S net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08443_ reg_pc\[25\] _03842_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_82_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ _03786_ _03790_ net766 VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__mux2_1
XANTENNA__13052__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07325_ _02865_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__inv_2
XFILLER_149_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout1060_A net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_A _02357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09648__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07256_ count_cycle\[7\] net971 net841 _02801_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__o211a_1
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07187_ net3 net20 net1048 VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__mux2_1
XFILLER_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08231__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_A _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1113_X net1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11118__A1 net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12802__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout421 net422 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_4
XANTENNA__09383__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout432 net434 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__buf_4
XFILLER_87_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input9_X net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout443 net444 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__buf_4
Xfanout454 _02122_ VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__buf_2
XANTENNA_fanout952_A net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11418__S net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 _02117_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__buf_4
Xfanout476 _04292_ VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_4
Xfanout487 _04288_ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__buf_4
X_09828_ net1182 _04437_ _04613_ _02489_ net847 VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout498 net499 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__buf_4
XANTENNA_fanout740_X net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09759_ _04545_ _04548_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout838_X net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12770_ net1219 genblk1.genblk1.pcpi_mul.next_rs1\[38\] net2480 net908 net764 VGND
+ VGND VPWR VPWR _01409_ sky130_fd_sc_hd__a221o_1
XFILLER_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11721_ is_beq_bne_blt_bge_bltu_bgeu _06237_ net561 VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__o21a_1
XFILLER_70_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14440_ clknet_leaf_64_clk _00829_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dfxtp_1
X_11652_ net1740 net30 net548 VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__mux2_1
XFILLER_30_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13043__A1 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10603_ cpuregs\[11\]\[7\] net630 net595 _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__o211a_1
XANTENNA__11054__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14371_ clknet_leaf_167_clk _00792_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dfxtp_4
X_11583_ net1234 is_alu_reg_imm net746 VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_137_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13322_ _02409_ net754 VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__nand2_1
XANTENNA__08462__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10534_ cpuregs\[25\]\[5\] net629 net609 _05228_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__o211a_1
XANTENNA__06771__A net1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13253_ net1038 net396 _02178_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__o21ba_1
X_10465_ cpuregs\[27\]\[0\] net634 net600 _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__o211a_1
XFILLER_89_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12204_ net748 _06594_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__nor2_1
XANTENNA__08222__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13184_ net1515 net329 net427 VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__mux2_1
X_10396_ net1169 net1168 _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__or3_1
XANTENNA__08222__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12135_ _06388_ _06401_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__nand2_1
XANTENNA__09293__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12066_ net1011 _06508_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__or2_1
XFILLER_49_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11017_ cpuregs\[26\]\[18\] net648 VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__or2_1
XANTENNA__11555__C net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13543__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ net1397 net586 net449 VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08864__C net1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14707_ clknet_leaf_162_clk _01092_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_11919_ genblk2.pcpi_div.divisor\[59\] genblk2.pcpi_div.divisor\[58\] genblk2.pcpi_div.divisor\[57\]
+ genblk2.pcpi_div.divisor\[56\] VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__or4_1
X_12899_ net576 net1907 net456 VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__mux2_1
X_14638_ clknet_leaf_169_clk _01023_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__11045__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14569_ clknet_leaf_57_clk _00955_ VGND VGND VPWR VPWR cpuregs\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07110_ genblk2.pcpi_div.dividend\[28\] _02667_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__nand2_1
XFILLER_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07777__A net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08090_ _03343_ _03347_ _03576_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__and3_1
Xclkload20 clknet_leaf_194_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__10915__B decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07041_ _02608_ _02609_ _02606_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__o21ai_1
Xclkload31 clknet_leaf_184_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__inv_6
XFILLER_161_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__inv_8
Xclkload53 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload53/X sky130_fd_sc_hd__clkbuf_4
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload64 clknet_leaf_165_clk VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__clkinv_4
Xclkload75 clknet_leaf_158_clk VGND VGND VPWR VPWR clkload75/Y sky130_fd_sc_hd__inv_12
Xclkload86 clknet_leaf_175_clk VGND VGND VPWR VPWR clkload86/X sky130_fd_sc_hd__clkbuf_8
Xclkload97 clknet_leaf_148_clk VGND VGND VPWR VPWR clkload97/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10556__C1 net830 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08992_ _04272_ _04273_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__or2_1
XANTENNA__10571__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07943_ net1181 net1053 net933 _03458_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__a31o_1
XANTENNA__11238__S net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__B1 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07874_ _03389_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08120__B net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09613_ reg_pc\[12\] net875 _04433_ net845 VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__a22o_1
X_06825_ instr_sw instr_sh net970 _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__or4_1
X_09544_ count_instr\[48\] _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__or2_1
X_06756_ net1145 VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__inv_2
XFILLER_24_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11284__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11481__B net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09475_ count_instr\[23\] count_instr\[22\] VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout533_A net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08426_ reg_out\[22\] alu_out_q\[22\] net1155 VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__mux2_1
XFILLER_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11036__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08357_ _03775_ _03776_ net766 VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout700_A net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload3 clknet_4_3_0_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_8
XANTENNA_fanout419_X net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11701__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09378__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07308_ _02848_ _02849_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__xor2_1
XFILLER_149_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08282__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08288_ reg_out\[21\] reg_next_pc\[21\] net926 VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__mux2_1
XFILLER_125_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13201__B _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07239_ count_cycle\[6\] net972 net841 _02785_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10250_ _04949_ _04954_ _04955_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__nand3_1
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout788_X net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10181_ _02464_ _04882_ _04886_ _02459_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10841__A net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1205 _02378_ VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__buf_2
Xfanout1216 net1222 VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__buf_2
Xfanout1227 net1241 VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__buf_2
Xfanout1238 net1239 VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout955_X net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout273 net275 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_4
X_13940_ clknet_leaf_178_clk _00394_ VGND VGND VPWR VPWR cpuregs\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout284 _03870_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_2
Xfanout295 net296 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13871_ clknet_leaf_47_clk _00325_ VGND VGND VPWR VPWR cpuregs\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15610_ clknet_leaf_12_clk _01946_ VGND VGND VPWR VPWR cpuregs\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12822_ net306 net2058 net466 VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__mux2_1
XANTENNA__08457__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15541_ clknet_leaf_1_clk _01877_ VGND VGND VPWR VPWR cpuregs\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12753_ net1641 net899 _02110_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__a21o_1
X_11704_ net1888 net322 net374 VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__mux2_1
X_15472_ clknet_leaf_192_clk _01808_ VGND VGND VPWR VPWR cpuregs\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12684_ net1196 net2928 net888 net2948 net711 VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_42_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ clknet_leaf_76_clk alu_out\[23\] VGND VGND VPWR VPWR alu_out_q\[23\] sky130_fd_sc_hd__dfxtp_1
X_11635_ net2398 _06174_ _06176_ net731 VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06772__Y _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09288__S net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14354_ clknet_leaf_85_clk _00776_ VGND VGND VPWR VPWR mem_do_rinst sky130_fd_sc_hd__dfxtp_2
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11566_ net1649 net562 _06178_ _06184_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__a22o_1
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13305_ net1031 net752 _02223_ net708 VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__o211a_1
XFILLER_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10517_ net801 _05209_ _05211_ net838 VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__a211o_1
X_14285_ clknet_leaf_97_clk _00739_ VGND VGND VPWR VPWR count_cycle\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11497_ net2542 _06158_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__nor2_1
XANTENNA__08205__B net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12527__B1 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13236_ net959 _04960_ _02159_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__a31o_1
X_10448_ cpuregs\[8\]\[0\] cpuregs\[9\]\[0\] net686 VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__mux2_1
XANTENNA__13538__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12442__S net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13167_ net1915 net583 net429 VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__mux2_1
X_10379_ genblk2.pcpi_div.quotient_msk\[11\] genblk2.pcpi_div.quotient_msk\[10\] genblk2.pcpi_div.quotient_msk\[9\]
+ genblk2.pcpi_div.quotient_msk\[8\] VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__or4_1
XANTENNA__10553__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08859__C net1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12118_ _06266_ _06383_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__xnor2_1
X_13098_ _04272_ _04283_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__or2_1
XFILLER_2_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12049_ net1019 net1016 net1015 _06484_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__or4_1
XFILLER_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07590_ reg_pc\[30\] decoded_imm\[30\] VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__or2_1
XANTENNA__08367__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1306 VGND VGND VPWR VPWR picorv32_1306/HI trace_data[28] sky130_fd_sc_hd__conb_1
XFILLER_61_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09260_ net2002 net283 net490 VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__mux2_1
X_08211_ _03368_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__or2_1
XANTENNA__11018__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09191_ net293 net2051 net498 VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11521__S net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09198__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08142_ _03635_ _03636_ _02364_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__mux2_1
XFILLER_119_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15497__Q net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08073_ _03379_ _03559_ _03286_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__and3b_1
Xclkload120 clknet_leaf_77_clk VGND VGND VPWR VPWR clkload120/X sky130_fd_sc_hd__clkbuf_4
Xclkload131 clknet_leaf_62_clk VGND VGND VPWR VPWR clkload131/Y sky130_fd_sc_hd__inv_12
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload142 clknet_leaf_82_clk VGND VGND VPWR VPWR clkload142/Y sky130_fd_sc_hd__clkinv_2
Xclkload153 clknet_leaf_113_clk VGND VGND VPWR VPWR clkload153/Y sky130_fd_sc_hd__inv_6
X_07024_ net1116 genblk2.pcpi_div.quotient\[15\] _02593_ net950 VGND VGND VPWR VPWR
+ _02595_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_77_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload164 clknet_leaf_124_clk VGND VGND VPWR VPWR clkload164/Y sky130_fd_sc_hd__inv_8
Xclkload175 clknet_leaf_95_clk VGND VGND VPWR VPWR clkload175/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload186 clknet_leaf_108_clk VGND VGND VPWR VPWR clkload186/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08198__B1 net969 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10544__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11741__A1 net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08975_ net1424 _04264_ net946 VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__mux2_1
XFILLER_29_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold15 _01392_ VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 cpuregs\[26\]\[12\] VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold37 cpuregs\[24\]\[11\] VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07926_ _03272_ _03380_ _03439_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__and3_1
Xhold48 cpuregs\[26\]\[9\] VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold59 net50 VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout650_A net654 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07857_ net1162 net1020 VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout271_X net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout748_A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13183__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06808_ mem_do_rinst mem_do_prefetch VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__or2_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08277__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07788_ _03303_ _03305_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09527_ _04381_ net1227 _04380_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout915_A net919 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_X net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09458_ count_instr\[15\] _04330_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__and3_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11009__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08409_ net328 net2379 net528 VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__mux2_1
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09389_ net2332 net304 net402 VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__mux2_1
XFILLER_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11420_ cpuregs\[24\]\[29\] net706 VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__or2_1
XANTENNA__12221__A2 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11351_ cpuregs\[27\]\[27\] net639 net599 _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__o211a_1
XFILLER_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10302_ _05003_ _05005_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__or3_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14070_ clknet_leaf_185_clk _00524_ VGND VGND VPWR VPWR cpuregs\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11282_ _05955_ _05956_ net808 VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__mux2_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08189__B1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11667__A is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13021_ net331 net2462 net443 VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__mux2_1
XANTENNA__09925__A1 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10233_ decoded_imm\[7\] net1035 VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__nor2_1
XFILLER_79_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08312__Y _03741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10164_ net2797 _04871_ net1238 VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__o21ai_1
Xfanout1002 net1003 VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__buf_2
Xfanout1013 net213 VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__buf_4
XANTENNA__07400__A2 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1024 net1025 VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1035 net1037 VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__buf_2
Xfanout1046 net225 VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1057 net1059 VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__buf_2
X_14972_ clknet_leaf_143_clk _01324_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_10095_ count_cycle\[35\] _04826_ count_cycle\[36\] VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__a21o_1
Xfanout1068 net1070 VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 cpu_state\[3\] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13923_ clknet_leaf_16_clk _00377_ VGND VGND VPWR VPWR cpuregs\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07164__A1 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12693__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13093__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13854_ clknet_leaf_10_clk _00308_ VGND VGND VPWR VPWR cpuregs\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13237__A1 net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06911__B2 net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12805_ net527 net2242 net463 VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__mux2_1
XANTENNA__11248__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13785_ clknet_leaf_5_clk _00239_ VGND VGND VPWR VPWR cpuregs\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10997_ cpuregs\[4\]\[18\] cpuregs\[5\]\[18\] net652 VGND VGND VPWR VPWR _05679_
+ sky130_fd_sc_hd__mux2_1
X_15524_ clknet_leaf_86_clk _01860_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dfxtp_1
X_12736_ net1190 genblk1.genblk1.pcpi_mul.next_rs1\[17\] net914 net1015 VGND VGND
+ VPWR VPWR _02102_ sky130_fd_sc_hd__a22o_1
XFILLER_30_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12460__A2 net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10471__A1 net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15455_ clknet_leaf_51_clk _01794_ VGND VGND VPWR VPWR cpuregs\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12667_ genblk1.genblk1.pcpi_mul.instr_mulh _02082_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__and2_2
XFILLER_129_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12437__S net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12748__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14406_ clknet_leaf_136_clk alu_out\[6\] VGND VGND VPWR VPWR alu_out_q\[6\] sky130_fd_sc_hd__dfxtp_1
X_11618_ mem_rdata_q\[23\] mem_rdata_q\[22\] mem_rdata_q\[21\] VGND VGND VPWR VPWR
+ _06207_ sky130_fd_sc_hd__or3_1
XANTENNA__07219__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15386_ clknet_leaf_43_clk _01725_ VGND VGND VPWR VPWR cpuregs\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12598_ net301 net2179 net470 VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14337_ clknet_leaf_26_clk _06724_ VGND VGND VPWR VPWR reg_out\[17\] sky130_fd_sc_hd__dfxtp_1
X_11549_ _06165_ _06171_ _06172_ net547 VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__o31a_1
XFILLER_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold507 cpuregs\[30\]\[4\] VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 cpuregs\[12\]\[26\] VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold529 cpuregs\[25\]\[14\] VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ clknet_leaf_129_clk _00722_ VGND VGND VPWR VPWR count_cycle\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09916__A1 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13219_ net1063 net1038 net754 net557 VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a31o_1
XFILLER_124_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07774__B net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14199_ clknet_leaf_174_clk _00653_ VGND VGND VPWR VPWR reg_pc\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10526__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1207 genblk1.genblk1.pcpi_mul.next_rs1\[33\] VGND VGND VPWR VPWR net2521 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ genblk1.genblk1.pcpi_mul.rd\[43\] genblk1.genblk1.pcpi_mul.next_rs2\[44\]
+ net1091 VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__nand3_1
XANTENNA__12900__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1218 cpuregs\[3\]\[0\] VGND VGND VPWR VPWR net2532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1229 genblk2.pcpi_div.divisor\[47\] VGND VGND VPWR VPWR net2543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07790__A net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07711_ decoded_imm_j\[3\] _02701_ _03192_ _03230_ _03228_ VGND VGND VPWR VPWR _06749_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__12684__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08691_ genblk1.genblk1.pcpi_mul.next_rs2\[33\] net1101 _04050_ _04052_ VGND VGND
+ VPWR VPWR _04053_ sky130_fd_sc_hd__a22o_1
XANTENNA__07155__A1 _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11516__S net738 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07642_ cpuregs\[8\]\[2\] net700 VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__or2_1
XFILLER_54_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07573_ net359 _03092_ _03097_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_24_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09312_ net1379 net344 net479 VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__mux2_1
X_09243_ net1892 net347 net488 VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout329_A _03818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09174_ net403 net2021 net496 VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__mux2_1
X_08125_ net1144 _03328_ _03621_ _03620_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__o31a_1
XFILLER_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1140_A instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _03286_ _03559_ _03558_ _03546_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07630__A2 decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13178__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout698_A net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07007_ net1115 _02578_ genblk2.pcpi_div.dividend\[13\] VGND VGND VPWR VPWR _02580_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_150_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput38 net38 VGND VGND VPWR VPWR mem_addr[13] sky130_fd_sc_hd__buf_2
Xoutput49 net49 VGND VGND VPWR VPWR mem_addr[24] sky130_fd_sc_hd__buf_2
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1026_X net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12911__A0 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout486_X net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12810__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08958_ genblk1.genblk1.pcpi_mul.rd\[17\] genblk1.genblk1.pcpi_mul.rd\[49\] net955
+ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__mux2_1
XANTENNA__09391__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1730 decoded_imm_j\[19\] VGND VGND VPWR VPWR net3044 sky130_fd_sc_hd__dlygate4sd3_1
X_07909_ _03311_ _03426_ _03418_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__a21oi_1
Xhold1741 decoded_imm\[16\] VGND VGND VPWR VPWR net3055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1752 count_instr\[26\] VGND VGND VPWR VPWR net3066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12675__C1 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _04215_ _04218_ _04216_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__a21bo_1
XFILLER_29_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11426__S net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10686__D1 net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10920_ _05602_ _05603_ net811 VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__mux2_1
XFILLER_84_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13207__A net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10851_ cpuregs\[14\]\[14\] cpuregs\[15\]\[14\] net653 VGND VGND VPWR VPWR _05537_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout820_X net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout918_X net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_160_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13570_ net336 net2214 net411 VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__mux2_1
XFILLER_25_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10782_ cpuregs\[16\]\[12\] net646 VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__or2_1
XFILLER_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12521_ net2664 net385 _02011_ _02012_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__a22o_1
XFILLER_157_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07859__B net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15240_ clknet_leaf_7_clk _01581_ VGND VGND VPWR VPWR cpuregs\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12452_ _05098_ net717 net1174 VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_175_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11403_ cpuregs\[5\]\[29\] net644 net820 _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__o211a_1
X_15171_ clknet_leaf_66_clk _01520_ VGND VGND VPWR VPWR mem_rdata_q\[22\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_10_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12383_ net1341 net303 net362 VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14122_ clknet_leaf_52_clk _00576_ VGND VGND VPWR VPWR cpuregs\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11334_ net840 _06004_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07621__A2 decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13088__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14053_ clknet_leaf_38_clk _00507_ VGND VGND VPWR VPWR cpuregs\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11265_ net820 _05937_ _05939_ net836 VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_37_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11705__A1 net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13004_ net584 net2280 net445 VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__mux2_1
X_10216_ _04917_ _04921_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__nand2_1
X_11196_ net835 _05868_ _05870_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__a211o_1
XANTENNA_output248_A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10147_ net3045 _04860_ _04862_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__o21a_1
XFILLER_95_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ clknet_leaf_120_clk _01307_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10078_ count_cycle\[29\] _04816_ _04818_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_50_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13906_ clknet_leaf_23_clk _00360_ VGND VGND VPWR VPWR cpuregs\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10141__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07688__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14886_ clknet_leaf_49_clk _01238_ VGND VGND VPWR VPWR cpuregs\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13837_ clknet_leaf_49_clk _00291_ VGND VGND VPWR VPWR cpuregs\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13551__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10179__C _04883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13768_ clknet_leaf_57_clk _00222_ VGND VGND VPWR VPWR cpuregs\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15507_ clknet_leaf_167_clk _01843_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dfxtp_1
X_12719_ net1190 genblk1.genblk1.pcpi_mul.next_rs1\[8\] net1542 net883 _02093_ VGND
+ VGND VPWR VPWR _01379_ sky130_fd_sc_hd__a221o_1
XFILLER_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07769__B net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ clknet_leaf_112_clk _00153_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10995__A2 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15438_ clknet_leaf_193_clk _01777_ VGND VGND VPWR VPWR cpuregs\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15369_ clknet_leaf_22_clk _01708_ VGND VGND VPWR VPWR cpuregs\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11944__A1 _02443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07073__B1 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07785__A net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold304 cpuregs\[31\]\[23\] VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 genblk1.genblk1.pcpi_mul.pcpi_rd\[26\] VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08380__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold326 cpuregs\[13\]\[4\] VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 cpuregs\[23\]\[3\] VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10923__B net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold348 cpuregs\[8\]\[28\] VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ net1127 _04446_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__nor2_1
Xhold359 net156 VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout806 _03143_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__buf_2
X_09861_ _04629_ _04640_ _04642_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__and3_1
Xfanout817 net818 VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__buf_4
Xfanout828 net830 VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout839 _03136_ VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__buf_4
X_08812_ genblk1.genblk1.pcpi_mul.rd\[51\] genblk1.genblk1.pcpi_mul.next_rs2\[52\]
+ net1099 VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__nand3_1
XFILLER_58_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09792_ decoded_imm_j\[14\] _04435_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__or2_1
XFILLER_97_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1004 cpuregs\[10\]\[24\] VGND VGND VPWR VPWR net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13449__A1 net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1015 cpuregs\[1\]\[22\] VGND VGND VPWR VPWR net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 cpuregs\[7\]\[0\] VGND VGND VPWR VPWR net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1037 cpuregs\[1\]\[13\] VGND VGND VPWR VPWR net2351 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ genblk1.genblk1.pcpi_mul.next_rs2\[41\] net1091 _04094_ _04096_ VGND VGND
+ VPWR VPWR _04097_ sky130_fd_sc_hd__a22o_1
Xhold1048 instr_slli VGND VGND VPWR VPWR net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 cpuregs\[21\]\[28\] VGND VGND VPWR VPWR net2373 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__B2 net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_A _03873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08674_ _04038_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_77_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _03144_ _03145_ net819 VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13461__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07556_ net359 _03076_ _03081_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_85_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06864__A net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08408__X _03818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07487_ net358 _03012_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__o21bai_1
XFILLER_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09226_ net1829 net287 net495 VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__mux2_1
XFILLER_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13385__B1 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09157_ net2093 net299 net503 VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout401_X net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12805__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout1143_X net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11935__A1 _02384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08108_ _03328_ net931 net969 VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__o21a_1
XANTENNA__09386__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08290__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11929__B _06398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09088_ net1456 net294 net510 VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net983 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08039_ _03357_ _03362_ _03544_ _03361_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_147_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold860 _01136_ VGND VGND VPWR VPWR net2174 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11010__A net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold871 cpuregs\[3\]\[9\] VGND VGND VPWR VPWR net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 cpuregs\[3\]\[14\] VGND VGND VPWR VPWR net2196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold893 cpuregs\[11\]\[9\] VGND VGND VPWR VPWR net2207 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ cpuregs\[22\]\[19\] cpuregs\[23\]\[19\] net680 VGND VGND VPWR VPWR _05731_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout770_X net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_X net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10001_ count_cycle\[0\] count_cycle\[1\] count_cycle\[2\] VGND VGND VPWR VPWR _04769_
+ sky130_fd_sc_hd__a21o_1
XFILLER_92_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1560 _01134_ VGND VGND VPWR VPWR net2874 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1571 count_cycle\[19\] VGND VGND VPWR VPWR net2885 sky130_fd_sc_hd__dlygate4sd3_1
X_14740_ clknet_leaf_161_clk _01125_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11952_ net1046 _02443_ _06409_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__o21a_1
Xhold1582 instr_sw VGND VGND VPWR VPWR net2896 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1593 _00710_ VGND VGND VPWR VPWR net2907 sky130_fd_sc_hd__dlygate4sd3_1
X_10903_ cpuregs\[27\]\[15\] net617 net589 _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__o211a_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14671_ clknet_leaf_153_clk net2786 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11883_ _06344_ _06353_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__nor2_1
XFILLER_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13622_ clknet_leaf_49_clk _00077_ VGND VGND VPWR VPWR cpuregs\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_10834_ cpuregs\[16\]\[13\] net650 VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__or2_1
XFILLER_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08318__X _03746_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13553_ _03742_ _04275_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__or2_4
XFILLER_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10765_ net789 _05449_ _05451_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__or4_1
XFILLER_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12504_ genblk2.pcpi_div.divisor\[47\] net870 VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__or2_1
XFILLER_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13484_ net1343 net287 net425 VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__mux2_1
XFILLER_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10696_ net1076 decoded_imm\[9\] VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__or2_1
X_15223_ clknet_leaf_79_clk _01564_ VGND VGND VPWR VPWR reg_sh\[0\] sky130_fd_sc_hd__dfxtp_1
X_12435_ _06670_ _06671_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10729__A2 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15154_ clknet_leaf_89_clk _01503_ VGND VGND VPWR VPWR mem_rdata_q\[5\] sky130_fd_sc_hd__dfxtp_1
X_12366_ net1547 net522 net360 VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__mux2_1
XFILLER_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14105_ clknet_leaf_192_clk _00559_ VGND VGND VPWR VPWR cpuregs\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11317_ cpuregs\[22\]\[26\] cpuregs\[23\]\[26\] net702 VGND VGND VPWR VPWR _05991_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15085_ clknet_leaf_17_clk _01437_ VGND VGND VPWR VPWR cpuregs\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12297_ mem_rdata_q\[25\] net559 _06627_ net532 VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__a211o_1
X_14036_ clknet_leaf_179_clk _00490_ VGND VGND VPWR VPWR cpuregs\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output75_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248_ cpuregs\[11\]\[24\] net634 net597 _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__o211a_1
XFILLER_68_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07358__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07358__B2 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13546__S net418 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12450__S net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11179_ net1081 _05855_ net856 VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11574__B mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08307__A0 net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14938_ clknet_leaf_7_clk _01290_ VGND VGND VPWR VPWR cpuregs\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07530__A1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14869_ clknet_leaf_19_clk _01221_ VGND VGND VPWR VPWR cpuregs\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_07410_ count_instr\[49\] net1132 net1140 count_cycle\[49\] VGND VGND VPWR VPWR _02946_
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08375__S net529 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08390_ reg_out\[15\] alu_out_q\[15\] net1153 VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__mux2_1
XFILLER_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07341_ reg_pc\[12\] decoded_imm\[12\] _02867_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_34_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07272_ count_cycle\[8\] net971 net841 _02816_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__o211a_1
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09011_ net329 net1531 net516 VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__mux2_1
XANTENNA__13367__B1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10934__A net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 cpuregs\[14\]\[10\] VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 net135 VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__C net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold123 net148 VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 cpuregs\[12\]\[16\] VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold145 net55 VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 cpuregs\[13\]\[3\] VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 cpuregs\[22\]\[22\] VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _01372_ VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net1150 _04690_ _04691_ net1184 VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__o31a_1
Xfanout603 net606 VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkbuf_4
Xhold189 cpuregs\[24\]\[3\] VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout614 net616 VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__clkbuf_4
Xfanout625 net628 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_A net398 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12342__A1 decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13456__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout636 net639 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__clkbuf_4
Xfanout647 net649 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkbuf_4
X_09844_ decoded_imm_j\[18\] _04439_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__nand2_1
XANTENNA__12360__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout658 net663 VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06859__A net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout669 net672 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ net2675 net875 _04564_ net845 VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__a22o_1
X_06987_ net1119 _02562_ genblk2.pcpi_div.quotient\[10\] VGND VGND VPWR VPWR _02563_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08726_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11302__C1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08657_ genblk1.genblk1.pcpi_mul.next_rs2\[28\] net1105 genblk1.genblk1.pcpi_mul.rd\[27\]
+ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout730_A _06244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13191__S net430 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_929 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout828_A net830 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11704__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_X net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ count_instr\[31\] net1137 net978 _03129_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__a211o_1
XANTENNA__08285__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08588_ genblk1.genblk1.pcpi_mul.next_rs2\[17\] net1094 _03962_ _03964_ VGND VGND
+ VPWR VPWR _03966_ sky130_fd_sc_hd__and4_1
XANTENNA__10828__B net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07539_ net1069 net1000 _03065_ net1085 VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__a22o_1
XFILLER_41_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_X net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10550_ net1172 net855 _05243_ _05244_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__a22o_1
XANTENNA__07285__B1 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09209_ net1427 net350 net492 VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__mux2_1
X_10481_ _05178_ _05179_ net804 VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__mux2_1
XFILLER_148_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11369__C1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12220_ net749 net2767 VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__nor2_1
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12030__B1 net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12151_ net2798 net378 net367 net2866 VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__a22o_1
XANTENNA__10592__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11102_ cpuregs\[11\]\[20\] net622 net591 _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__o211a_1
X_12082_ net1006 net724 _06528_ net863 VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__a31o_1
Xhold690 cpuregs\[25\]\[17\] VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12333__A1 decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12333__B2 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11033_ cpuregs\[4\]\[19\] cpuregs\[5\]\[19\] net684 VGND VGND VPWR VPWR _05714_
+ sky130_fd_sc_hd__mux2_1
XFILLER_150_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06769__A net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12097__B1 net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12984_ net2127 net338 net448 VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__mux2_1
Xhold1390 genblk2.pcpi_div.divisor\[12\] VGND VGND VPWR VPWR net2704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09501__A2 _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14723_ clknet_leaf_141_clk net2899 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11935_ _02384_ net873 _06405_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06775__Y _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14654_ clknet_leaf_155_clk _01039_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_11866_ _06306_ _06336_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__and2b_1
XANTENNA__10738__B net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13605_ clknet_leaf_187_clk _00060_ VGND VGND VPWR VPWR cpuregs\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10817_ net796 _05501_ _05503_ net823 VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__o211a_1
X_14585_ clknet_leaf_104_clk _00971_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11797_ genblk2.pcpi_div.dividend\[24\] genblk2.pcpi_div.divisor\[24\] VGND VGND
+ VPWR VPWR _06268_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_31_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ net339 net1817 net415 VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__mux2_1
X_10748_ cpuregs\[19\]\[11\] net625 net593 VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__o21a_1
X_13467_ net1994 net352 net423 VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__mux2_1
X_10679_ cpuregs\[30\]\[9\] cpuregs\[31\]\[9\] net670 VGND VGND VPWR VPWR _05370_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07028__B1 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15206_ clknet_leaf_72_clk _01555_ VGND VGND VPWR VPWR cpuregs\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12418_ net297 net1516 net473 VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__mux2_1
XANTENNA__11569__B net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13398_ net569 _05926_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__nor2_1
Xoutput206 net1027 VGND VGND VPWR VPWR pcpi_rs1[12] sky130_fd_sc_hd__buf_2
XANTENNA__10473__B net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput217 net1008 VGND VGND VPWR VPWR pcpi_rs1[22] sky130_fd_sc_hd__buf_2
X_15137_ clknet_leaf_16_clk _01489_ VGND VGND VPWR VPWR cpuregs\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput228 net228 VGND VGND VPWR VPWR pcpi_rs1[3] sky130_fd_sc_hd__buf_2
X_12349_ mem_rdata_q\[8\] _06617_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__and2_1
Xoutput239 net1163 VGND VGND VPWR VPWR pcpi_rs2[13] sky130_fd_sc_hd__buf_2
XFILLER_142_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15068_ clknet_leaf_104_clk net2265 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12324__A1 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14019_ clknet_leaf_13_clk _00473_ VGND VGND VPWR VPWR cpuregs\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_06910_ net1066 _02475_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__nand2_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07782__B net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07890_ net250 _02411_ _03335_ _03401_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__o221a_1
X_06841_ mem_do_rinst reg_pc\[1\] _02444_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10886__B2 net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09560_ count_instr\[51\] count_instr\[50\] _04395_ _04402_ VGND VGND VPWR VPWR _04403_
+ sky130_fd_sc_hd__and4_1
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06772_ net1185 VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__clkinv_4
XANTENNA__06829__D net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08511_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__inv_2
XFILLER_82_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09491_ net2892 _04356_ net1239 VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11524__S net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08442_ reg_out\[25\] alu_out_q\[25\] net1155 VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08373_ _03787_ _03788_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__nor2_1
XFILLER_149_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07324_ reg_pc\[12\] decoded_imm\[12\] VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__xor2_1
XANTENNA__07267__B1 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12260__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10810__A1 net797 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07255_ net1139 count_cycle\[39\] net976 _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout311_A _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06861__B net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08216__C1 net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07186_ _02735_ net1074 _02734_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__and3b_1
XFILLER_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09964__C1 net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08231__A2 net1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout400 _04293_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout680_A net696 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout411 _02358_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_8
Xfanout422 _02356_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__buf_4
XANTENNA__13186__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_X net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout433 net434 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_8
XFILLER_58_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout444 net446 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__buf_4
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout455 net456 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_4
Xfanout466 _02117_ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ _04611_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__nor2_1
Xfanout477 _04292_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_8
Xfanout488 _04287_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout945_A _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout499 _04285_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_2
XANTENNA__07742__B2 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09758_ _04548_ _04545_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__and2b_1
XFILLER_58_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_169_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08709_ genblk1.genblk1.pcpi_mul.next_rs2\[36\] net1098 genblk1.genblk1.pcpi_mul.rd\[35\]
+ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__a21o_1
XANTENNA__11287__D1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09689_ _04474_ _04485_ _04484_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_159_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10839__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11720_ instr_sltu instr_slt instr_sltiu instr_slti VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__or4_1
XFILLER_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__06848__A3 net965 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11651_ decoded_imm_j\[20\] net25 net547 VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout900_X net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10602_ cpuregs\[10\]\[7\] net673 VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__or2_1
X_14370_ clknet_leaf_167_clk _00791_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dfxtp_4
X_11582_ net2932 net741 _06181_ is_sb_sh_sw VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12251__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13321_ net960 _02237_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__nor2_1
XFILLER_168_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10533_ cpuregs\[24\]\[5\] net678 VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__or2_1
XFILLER_167_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08315__Y _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13252_ net568 _05278_ _02172_ net960 _02177_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__o221a_1
XFILLER_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ cpuregs\[26\]\[0\] net684 VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10293__B net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ net2785 net272 net2829 VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__a21oi_1
X_13183_ net1671 net334 net427 VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__mux2_1
XFILLER_124_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10565__B1 net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10395_ net1172 net1174 net1171 _05098_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__or4_1
XANTENNA__08222__A2 net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12134_ _06388_ _06401_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__or2_1
XFILLER_97_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08331__X _03756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13096__S net442 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12306__B2 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12065_ _06277_ _06514_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11016_ cpuregs\[25\]\[18\] net618 net603 _05697_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__o211a_1
XANTENNA_output230_A net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12967_ _03745_ _04281_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nor2_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13309__A1_N net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11918_ genblk2.pcpi_div.divisor\[61\] genblk2.pcpi_div.divisor\[60\] genblk2.pcpi_div.divisor\[62\]
+ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__or3_1
X_14706_ clknet_leaf_162_clk _01091_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_12898_ net579 net2099 net457 VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__mux2_1
XANTENNA__07123__A net1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14637_ clknet_leaf_163_clk _01022_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11849_ genblk2.pcpi_div.dividend\[0\] genblk2.pcpi_div.divisor\[0\] VGND VGND VPWR
+ VPWR _06320_ sky130_fd_sc_hd__nand2b_1
XFILLER_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14568_ clknet_leaf_60_clk _00954_ VGND VGND VPWR VPWR cpuregs\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12242__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13519_ net2022 net280 net421 VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__mux2_1
XANTENNA__07777__B net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14499_ clknet_leaf_96_clk _00888_ VGND VGND VPWR VPWR instr_or sky130_fd_sc_hd__dfxtp_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload10 clknet_4_10_0_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_16
X_07040_ net1114 genblk2.pcpi_div.quotient\[17\] _02607_ net950 VGND VGND VPWR VPWR
+ _02609_ sky130_fd_sc_hd__a31o_1
Xclkload21 clknet_leaf_195_clk VGND VGND VPWR VPWR clkload21/X sky130_fd_sc_hd__clkbuf_4
Xclkload32 clknet_leaf_185_clk VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinv_2
XFILLER_127_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload43 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload54/X sky130_fd_sc_hd__clkbuf_4
Xclkload65 clknet_leaf_166_clk VGND VGND VPWR VPWR clkload65/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload76 clknet_leaf_159_clk VGND VGND VPWR VPWR clkload76/Y sky130_fd_sc_hd__inv_12
XFILLER_126_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload87 clknet_leaf_138_clk VGND VGND VPWR VPWR clkload87/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__12903__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload98 clknet_leaf_150_clk VGND VGND VPWR VPWR clkload98/Y sky130_fd_sc_hd__clkinvlp_4
X_08991_ latched_rd\[1\] latched_rd\[0\] _03743_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__or3_4
XANTENNA__11519__S net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07942_ instr_and instr_andi VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__or2_1
XANTENNA__10859__A1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07873_ _02365_ _02366_ _02413_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_3_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09612_ _03792_ reg_next_pc\[12\] net920 VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__mux2_2
XFILLER_56_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08921__B1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06824_ instr_slt instr_slti instr_bgeu instr_bge VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__or4_1
XFILLER_84_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09543_ _04391_ net1230 _04390_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__and3b_1
X_06755_ net1072 VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__inv_2
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11254__S net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09474_ net1235 _04346_ _04347_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__and3_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08425_ net316 net2146 net530 VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08356_ reg_pc\[8\] _03772_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_154_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload4 clknet_4_4_0_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_22_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07307_ reg_pc\[10\] decoded_imm\[10\] _02837_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__a21o_1
XANTENNA__10394__A net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08287_ net1010 _03727_ net981 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__mux2_2
XFILLER_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1056_X net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07238_ count_instr\[6\] net1135 net976 _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_115_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09937__C1 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08204__A2 net933 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12813__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07169_ count_instr\[34\] net1130 net1135 count_instr\[2\] VGND VGND VPWR VPWR _02720_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1223_X net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09394__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10180_ instr_sll net756 instr_slli net1068 VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__or4b_1
XANTENNA__10841__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07963__A1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1206 net1207 VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__clkbuf_4
Xfanout1217 net1218 VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__buf_2
XANTENNA__09407__B net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1228 net1230 VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__clkbuf_2
Xfanout1239 net1240 VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout850_X net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout274 net275 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_4
Xfanout285 net286 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout948_X net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07715__A1 net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout296 _03857_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13870_ clknet_leaf_38_clk _00324_ VGND VGND VPWR VPWR cpuregs\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12821_ net309 net2257 net464 VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__mux2_1
X_15540_ clknet_leaf_194_clk _01876_ VGND VGND VPWR VPWR cpuregs\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12752_ net1214 net1550 net918 net1001 VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__a22o_1
XFILLER_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11703_ net2149 net326 net375 VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__mux2_1
X_15471_ clknet_leaf_192_clk _01807_ VGND VGND VPWR VPWR cpuregs\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12683_ net1194 genblk1.genblk1.pcpi_mul.next_rs2\[48\] net886 net2915 net711 VGND
+ VGND VPWR VPWR _01353_ sky130_fd_sc_hd__a221o_1
XANTENNA__11027__A1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14422_ clknet_leaf_76_clk alu_out\[22\] VGND VGND VPWR VPWR alu_out_q\[22\] sky130_fd_sc_hd__dfxtp_1
X_11634_ net1208 _02400_ _06210_ _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_42_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08473__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14772__Q genblk2.pcpi_div.pcpi_rd\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14353_ clknet_leaf_85_clk _00775_ VGND VGND VPWR VPWR mem_do_prefetch sky130_fd_sc_hd__dfxtp_1
X_11565_ mem_rdata_q\[12\] mem_rdata_q\[13\] mem_rdata_q\[14\] VGND VGND VPWR VPWR
+ _06184_ sky130_fd_sc_hd__and3b_1
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13304_ _02408_ net754 VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__nand2_1
X_10516_ cpuregs\[5\]\[5\] net630 net815 _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__o211a_1
X_14284_ clknet_leaf_97_clk _00738_ VGND VGND VPWR VPWR count_cycle\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07651__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11496_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__inv_2
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12527__A1 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13235_ net709 _02137_ _02161_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__a31o_1
X_10447_ cpuregs\[11\]\[0\] net634 net600 _05146_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__o211a_1
X_13166_ net2059 net588 net429 VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__mux2_1
X_10378_ genblk2.pcpi_div.pcpi_wait_q genblk2.pcpi_div.pcpi_wait VGND VGND VPWR VPWR
+ _05083_ sky130_fd_sc_hd__nand2b_1
XFILLER_151_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12117_ net997 net725 _06558_ net864 VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__a31o_1
XFILLER_112_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13097_ net279 net2175 net442 VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__mux2_1
XANTENNA__12024__A net1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12048_ net3021 _06500_ net269 VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__mux2_1
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13554__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10710__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13999_ clknet_leaf_45_clk _00453_ VGND VGND VPWR VPWR cpuregs\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10198__B net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1307 VGND VGND VPWR VPWR picorv32_1307/HI trace_data[29] sky130_fd_sc_hd__conb_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08210_ net1145 _03370_ _03696_ _03695_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__o31a_1
X_09190_ net297 net1945 net498 VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__mux2_1
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08141_ _03322_ _03629_ _03319_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__a21o_1
XFILLER_119_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10777__B1 net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09631__B2 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08072_ _03379_ _03546_ _03558_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__nor3_1
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload110 clknet_leaf_45_clk VGND VGND VPWR VPWR clkload110/X sky130_fd_sc_hd__clkbuf_4
Xclkload121 clknet_leaf_50_clk VGND VGND VPWR VPWR clkload121/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload132 clknet_leaf_65_clk VGND VGND VPWR VPWR clkload132/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload143 clknet_leaf_83_clk VGND VGND VPWR VPWR clkload143/Y sky130_fd_sc_hd__bufinv_16
X_07023_ net1115 _02593_ genblk2.pcpi_div.quotient\[15\] VGND VGND VPWR VPWR _02594_
+ sky130_fd_sc_hd__a21oi_1
Xclkload154 clknet_leaf_114_clk VGND VGND VPWR VPWR clkload154/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload165 clknet_leaf_125_clk VGND VGND VPWR VPWR clkload165/Y sky130_fd_sc_hd__inv_6
Xclkload176 clknet_leaf_96_clk VGND VGND VPWR VPWR clkload176/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__10529__B1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload187 clknet_leaf_109_clk VGND VGND VPWR VPWR clkload187/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07900__A_N net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08974_ genblk1.genblk1.pcpi_mul.rd\[25\] genblk1.genblk1.pcpi_mul.rd\[57\] net956
+ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__mux2_1
XFILLER_69_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold16 reg_next_pc\[1\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 cpuregs\[26\]\[25\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _03297_ _03442_ _03396_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_90_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold38 net38 VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold49 net39 VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13464__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11773__A _06245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07856_ net1162 net1020 VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__and2_1
XFILLER_84_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06807_ genblk1.genblk1.pcpi_mul.mul_counter\[5\] VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__inv_2
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07787_ net1174 net1043 VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout643_A net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09526_ count_instr\[41\] count_instr\[40\] _04377_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09457_ count_instr\[17\] count_instr\[16\] VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout431_X net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout810_A net812 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12808__S net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout1173_X net1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11712__S net376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09389__S net402 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08408_ _03816_ _03817_ net767 VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09388_ net2018 net307 net401 VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__mux2_1
XANTENNA__08293__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12757__A1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08339_ reg_out\[5\] alu_out_q\[5\] net1154 VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__mux2_1
XANTENNA__12757__B2 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11350_ cpuregs\[26\]\[27\] net693 VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__or2_1
XFILLER_125_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10301_ _04913_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout898_X net898 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11281_ cpuregs\[30\]\[25\] cpuregs\[31\]\[25\] net704 VGND VGND VPWR VPWR _05956_
+ sky130_fd_sc_hd__mux2_1
X_13020_ net334 net2235 net443 VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__mux2_1
XFILLER_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10232_ decoded_imm\[7\] net1035 VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__nand2_1
XANTENNA__11667__B mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11193__B1 net611 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11732__A2 _06242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ count_cycle\[58\] count_cycle\[59\] count_cycle\[60\] _04868_ VGND VGND VPWR
+ VPWR _04873_ sky130_fd_sc_hd__and4_2
XFILLER_126_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1003 net220 VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__buf_4
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10940__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1014 net1015 VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1025 net207 VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__buf_2
Xfanout1036 net1037 VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__clkbuf_2
Xfanout1047 net1049 VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10998__S net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14971_ clknet_leaf_143_clk _01323_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_10094_ net3030 _04826_ _04828_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__o21a_1
Xfanout1058 net1059 VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__clkbuf_2
Xfanout1069 net1070 VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__clkbuf_2
X_13922_ clknet_leaf_15_clk _00376_ VGND VGND VPWR VPWR cpuregs\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08468__S net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13853_ clknet_leaf_199_clk _00307_ VGND VGND VPWR VPWR cpuregs\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13237__A2 net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12804_ net538 net1846 net463 VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10996_ cpuregs\[6\]\[18\] cpuregs\[7\]\[18\] net652 VGND VGND VPWR VPWR _05678_
+ sky130_fd_sc_hd__mux2_1
X_13784_ clknet_leaf_181_clk _00238_ VGND VGND VPWR VPWR cpuregs\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15523_ clknet_leaf_86_clk _01859_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dfxtp_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12735_ net1191 net2197 net2364 net884 _02101_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__a221o_1
XANTENNA__09299__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15454_ clknet_leaf_56_clk _01793_ VGND VGND VPWR VPWR cpuregs\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12666_ net1218 genblk1.genblk1.pcpi_mul.next_rs2\[32\] net905 net3023 _02082_ VGND
+ VGND VPWR VPWR _01337_ sky130_fd_sc_hd__a221o_1
XFILLER_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10471__A2 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11617_ mem_rdata_q\[27\] mem_rdata_q\[26\] _06204_ _06205_ VGND VGND VPWR VPWR _06206_
+ sky130_fd_sc_hd__and4bb_1
X_14405_ clknet_leaf_135_clk alu_out\[5\] VGND VGND VPWR VPWR alu_out_q\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12748__B2 net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15385_ clknet_leaf_15_clk _01724_ VGND VGND VPWR VPWR cpuregs\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12597_ net306 net2381 net469 VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11548_ net26 net23 VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__nand2_1
X_14336_ clknet_leaf_175_clk _06723_ VGND VGND VPWR VPWR reg_out\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08931__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold508 cpuregs\[23\]\[19\] VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13549__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold519 cpuregs\[10\]\[12\] VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14267_ clknet_leaf_122_clk _00721_ VGND VGND VPWR VPWR count_cycle\[12\] sky130_fd_sc_hd__dfxtp_1
X_11479_ net1157 net857 _06146_ _06147_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__a22o_1
X_13218_ _02474_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nand2_1
X_14198_ clknet_leaf_174_clk _00652_ VGND VGND VPWR VPWR reg_pc\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_115_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ net1448 net336 net432 VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10931__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 cpuregs\[19\]\[17\] VGND VGND VPWR VPWR net2522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 genblk2.pcpi_div.divisor\[41\] VGND VGND VPWR VPWR net2533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11593__A mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07710_ _02473_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__nand2_1
XANTENNA__07790__B net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10701__S net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08690_ genblk1.genblk1.pcpi_mul.rd\[32\] genblk1.genblk1.pcpi_mul.rdx\[32\] VGND
+ VGND VPWR VPWR _04052_ sky130_fd_sc_hd__or2_1
XANTENNA__08378__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07155__A2 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07641_ net807 _03159_ _03161_ net835 VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__o211a_1
XANTENNA__13228__A2 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06902__A2 is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12436__A0 net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09998__A net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07572_ net1068 net996 _03096_ net1085 _03095_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__a221o_1
XFILLER_80_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11239__B2 net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09311_ net1350 net348 net479 VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_15_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09242_ net1689 net350 net488 VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__mux2_1
XANTENNA__13313__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09002__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12739__B2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11104__Y _05784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09173_ net408 net1921 net496 VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__mux2_1
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08124_ _03329_ _03611_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__nor2_1
XANTENNA__11411__A1 net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13459__S net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08055_ _03287_ _03298_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__nand2_1
XANTENNA__12363__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1133_A net1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07006_ genblk2.pcpi_div.dividend\[13\] net1115 _02578_ VGND VGND VPWR VPWR _02579_
+ sky130_fd_sc_hd__and3_1
Xmax_cap761 _03883_ VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__clkbuf_1
Xoutput39 net39 VGND VGND VPWR VPWR mem_addr[14] sky130_fd_sc_hd__buf_2
XANTENNA_fanout593_A net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07918__A1 net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10922__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1019_X net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout760_A _04884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08957_ net2822 _04255_ net943 VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__mux2_1
XFILLER_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1720 count_instr\[54\] VGND VGND VPWR VPWR net3034 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13194__S net430 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout479_X net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11707__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1731 count_cycle\[54\] VGND VGND VPWR VPWR net3045 sky130_fd_sc_hd__dlygate4sd3_1
X_07908_ _03307_ _03419_ _03425_ net1043 _02393_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__a32o_1
X_08888_ net1217 net2949 net904 _04219_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__a22o_1
Xhold1742 decoded_imm\[19\] VGND VGND VPWR VPWR net3056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08288__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1753 count_cycle\[41\] VGND VGND VPWR VPWR net3067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07839_ net1166 net1029 VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__nand2_1
XANTENNA__13207__B net759 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13219__A2 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10850_ _05533_ _05535_ net781 VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__a21o_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09509_ count_instr\[35\] _04363_ _04368_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__and3_1
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10781_ _05467_ _05468_ net809 VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout813_X net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12538__S net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10989__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09843__B2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12520_ net871 _02009_ _02010_ net388 VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__a31oi_1
XANTENNA__11650__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07946__A_N is_compare VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12451_ _06683_ net2570 net383 VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__mux2_1
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11402_ cpuregs\[4\]\[29\] net706 VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__or2_1
X_15170_ clknet_leaf_65_clk _01519_ VGND VGND VPWR VPWR mem_rdata_q\[21\] sky130_fd_sc_hd__dfxtp_2
X_12382_ net1423 net307 net362 VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__mux2_1
XFILLER_165_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14121_ clknet_leaf_56_clk _00575_ VGND VGND VPWR VPWR cpuregs\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11333_ cpuregs\[1\]\[27\] net551 _06005_ net806 net833 VGND VGND VPWR VPWR _06006_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__07875__B net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14052_ clknet_leaf_44_clk _00506_ VGND VGND VPWR VPWR cpuregs\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11264_ net808 _05938_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__or2_1
XANTENNA__07594__C net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13003_ _03749_ net2328 net445 VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10215_ decoded_imm\[14\] net1022 VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__or2_1
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11195_ cpuregs\[18\]\[23\] net554 _05871_ net785 VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__o22a_1
X_10146_ count_cycle\[54\] _04860_ net1215 VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10077_ count_cycle\[29\] _04816_ net1209 VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__a21oi_1
X_14954_ clknet_leaf_34_clk _01306_ VGND VGND VPWR VPWR cpuregs\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07137__A2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09531__B1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13905_ clknet_leaf_22_clk _00359_ VGND VGND VPWR VPWR cpuregs\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14885_ clknet_leaf_48_clk _01237_ VGND VGND VPWR VPWR cpuregs\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_195_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_195_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkload2_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13836_ clknet_leaf_53_clk _00290_ VGND VGND VPWR VPWR cpuregs\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08926__S net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13767_ clknet_leaf_57_clk _00221_ VGND VGND VPWR VPWR cpuregs\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_10979_ cpuregs\[17\]\[17\] net617 net603 _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__o211a_1
X_15506_ clknet_leaf_167_clk _01842_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dfxtp_1
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12718_ _02403_ net911 VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__nor2_1
XANTENNA__11641__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13698_ clknet_leaf_116_clk _00152_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15437_ clknet_leaf_192_clk _01776_ VGND VGND VPWR VPWR cpuregs\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12649_ genblk1.genblk1.pcpi_mul.mul_waiting net1227 net250 VGND VGND VPWR VPWR _02074_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12197__A2 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15368_ clknet_leaf_30_clk _01707_ VGND VGND VPWR VPWR cpuregs\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11944__A2 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14319_ clknet_leaf_86_clk _00773_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dfxtp_1
Xhold305 cpuregs\[22\]\[25\] VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__B net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold316 cpuregs\[28\]\[20\] VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ clknet_leaf_105_clk _01640_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_finish
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold327 genblk1.genblk1.pcpi_mul.next_rs1\[26\] VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 cpuregs\[31\]\[11\] VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 cpuregs\[27\]\[14\] VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09860_ _04629_ _04642_ _04640_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__a21oi_1
Xfanout807 _03143_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__buf_4
XANTENNA__12911__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout818 net821 VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 net830 VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09770__B1 net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08811_ net892 _04152_ _04154_ net2652 net1195 VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__a32o_1
X_09791_ net2741 net875 _04576_ _04579_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__a22o_1
XFILLER_98_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1005 cpuregs\[5\]\[2\] VGND VGND VPWR VPWR net2319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13449__A2 net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1016 cpuregs\[9\]\[25\] VGND VGND VPWR VPWR net2330 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ genblk1.genblk1.pcpi_mul.rd\[40\] genblk1.genblk1.pcpi_mul.rdx\[40\] VGND
+ VGND VPWR VPWR _04096_ sky130_fd_sc_hd__or2_1
Xhold1027 cpuregs\[2\]\[4\] VGND VGND VPWR VPWR net2341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 cpuregs\[5\]\[31\] VGND VGND VPWR VPWR net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 cpuregs\[4\]\[24\] VGND VGND VPWR VPWR net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08673_ _04029_ _04032_ _04034_ _04036_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_186_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_186_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_132_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07624_ cpuregs\[4\]\[2\] cpuregs\[5\]\[2\] net700 VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ net1069 net999 _03080_ net1085 _03079_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout341_A _03807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12358__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout439_A net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11632__A1 net1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11093__C1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07486_ net1067 net1007 _03016_ net1082 _03015_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__a221o_1
XFILLER_139_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09225_ net1772 net292 net494 VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__mux2_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout606_A _03148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09156_ net1935 net303 net503 VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__mux2_1
XANTENNA__06880__A net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08424__X _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13189__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08107_ _03336_ net928 _03599_ _03605_ VGND VGND VPWR VPWR alu_out\[19\] sky130_fd_sc_hd__a211o_1
XANTENNA__11935__A2 net873 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08261__A0 net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09087_ net1719 net298 net511 VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__mux2_1
XANTENNA__12093__S net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1136_X net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07187__S net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08038_ _03360_ _03364_ _03528_ _03349_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__or4bb_1
Xhold850 cpuregs\[3\]\[23\] VGND VGND VPWR VPWR net2164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold861 cpuregs\[10\]\[31\] VGND VGND VPWR VPWR net2175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout596_X net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold872 cpuregs\[16\]\[31\] VGND VGND VPWR VPWR net2186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold883 genblk1.genblk1.pcpi_mul.next_rs1\[16\] VGND VGND VPWR VPWR net2197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12821__S net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold894 cpuregs\[2\]\[6\] VGND VGND VPWR VPWR net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06879__X _02478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ net2605 net2906 _04768_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__a21oi_1
X_09989_ net2607 net879 _04760_ net849 VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__a22o_1
XANTENNA__13218__A _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1550 instr_ori VGND VGND VPWR VPWR net2864 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_150_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1561 net190 VGND VGND VPWR VPWR net2875 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1572 genblk2.pcpi_div.quotient_msk\[23\] VGND VGND VPWR VPWR net2886 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_177_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_177_clk sky130_fd_sc_hd__clkbuf_8
X_11951_ net873 _06325_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout930_X net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1583 genblk1.genblk1.pcpi_mul.rd\[23\] VGND VGND VPWR VPWR net2897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1594 genblk2.pcpi_div.quotient\[2\] VGND VGND VPWR VPWR net2908 sky130_fd_sc_hd__dlygate4sd3_1
X_10902_ cpuregs\[26\]\[15\] net646 VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__or2_1
XFILLER_123_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11882_ _06299_ _06351_ _06352_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__or3_1
X_14670_ clknet_leaf_153_clk _01055_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10674__A2 net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13621_ clknet_leaf_71_clk _00076_ VGND VGND VPWR VPWR cpuregs\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_10833_ _05518_ _05519_ net797 VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__mux2_1
XFILLER_26_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09816__A1 net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09816__B2 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13552_ net278 net2186 net417 VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__mux2_1
X_10764_ cpuregs\[11\]\[11\] net625 net593 _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__o211a_1
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12503_ _05107_ net718 net241 VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__a21bo_1
XFILLER_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13483_ net1407 net290 net425 VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__mux2_1
X_10695_ net773 _05377_ _05385_ _05369_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__a31oi_4
XANTENNA__12179__A2 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13376__A1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12434_ net2811 _06669_ net917 VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__a21oi_1
X_15222_ clknet_leaf_87_clk _00011_ VGND VGND VPWR VPWR cpu_state\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__06790__A net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11387__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14780__Q genblk2.pcpi_div.pcpi_rd\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13099__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15153_ clknet_leaf_89_clk _01502_ VGND VGND VPWR VPWR mem_rdata_q\[4\] sky130_fd_sc_hd__dfxtp_1
X_12365_ net1522 net525 net360 VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__mux2_1
XANTENNA__07055__B2 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13400__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_101_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_91_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11316_ net836 _05985_ _05987_ _05989_ net794 VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__a2111o_1
X_14104_ clknet_leaf_186_clk _00558_ VGND VGND VPWR VPWR cpuregs\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15084_ clknet_leaf_32_clk _01436_ VGND VGND VPWR VPWR cpuregs\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12296_ decoded_imm\[25\] net733 VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__and2_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14035_ clknet_leaf_25_clk _00489_ VGND VGND VPWR VPWR cpuregs\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12887__A0 mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11247_ cpuregs\[10\]\[24\] net686 VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12351__A2 net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output68_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11178_ net1081 decoded_imm\[22\] VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__or2_1
XANTENNA__11347__S net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10129_ net2701 _04848_ _04850_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12639__B1 net919 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14937_ clknet_leaf_19_clk _01289_ VGND VGND VPWR VPWR cpuregs\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08858__A2 net1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13562__S net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06869__B2 net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14868_ clknet_leaf_6_clk _01220_ VGND VGND VPWR VPWR cpuregs\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13819_ clknet_leaf_196_clk _00273_ VGND VGND VPWR VPWR cpuregs\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14799_ clknet_leaf_81_clk _01151_ VGND VGND VPWR VPWR decoded_imm\[23\] sky130_fd_sc_hd__dfxtp_2
XFILLER_32_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07340_ _02877_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07271_ net1139 count_cycle\[40\] net976 _02815_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__a211o_1
XANTENNA__12906__S net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11090__A2 net624 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09010_ net334 net1741 net516 VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__mux2_1
XANTENNA__13367__A1 net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11378__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold102 cpuregs\[20\]\[25\] VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 cpuregs\[29\]\[12\] VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__D net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold124 cpuregs\[28\]\[21\] VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold135 cpuregs\[24\]\[4\] VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 genblk1.genblk1.pcpi_mul.pcpi_rd\[23\] VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 cpuregs\[20\]\[18\] VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 net139 VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 cpuregs\[12\]\[18\] VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _04443_ _04444_ _04672_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__and3_1
XANTENNA__12878__A0 mem_rdata_q\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout604 net606 VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__clkbuf_2
Xfanout615 net616 VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout626 net627 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12342__A2 net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout637 net639 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__buf_2
X_09843_ _04626_ _04627_ net2667 net877 VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__a2bb2o_1
Xfanout648 net649 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout291_A _03860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout659 net663 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout389_A net390 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06986_ genblk2.pcpi_div.quotient\[9\] _02556_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__or2_1
X_09774_ _04433_ _04563_ net1183 VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__mux2_1
XFILLER_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08725_ _04073_ _04076_ _04078_ _04080_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_159_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_159_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_174_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13472__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08656_ genblk1.genblk1.pcpi_mul.rd\[27\] genblk1.genblk1.pcpi_mul.next_rs2\[28\]
+ net1105 VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__nand3_1
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07607_ count_instr\[63\] net1133 net1141 count_cycle\[63\] VGND VGND VPWR VPWR _03129_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ genblk1.genblk1.pcpi_mul.next_rs2\[17\] net1094 _03962_ _03964_ VGND VGND
+ VPWR VPWR _03965_ sky130_fd_sc_hd__a22o_1
XANTENNA__10397__A net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_X net1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07538_ genblk1.genblk1.pcpi_mul.pcpi_rd\[26\] genblk2.pcpi_div.pcpi_rd\[26\] net1113
+ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_189_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07469_ count_instr\[53\] net1134 net1142 count_cycle\[53\] VGND VGND VPWR VPWR _03001_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout511_X net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06881__Y _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12816__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout609_X net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09208_ net1648 net354 net493 VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__mux2_1
XFILLER_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10480_ cpuregs\[14\]\[1\] cpuregs\[15\]\[1\] net683 VGND VGND VPWR VPWR _05179_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09139_ net1600 net523 net500 VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__mux2_1
XANTENNA__08234__A0 net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12150_ net2756 net378 net367 net2798 VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__a22o_1
XFILLER_136_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout880_X net880 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_X net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11101_ cpuregs\[10\]\[20\] net657 VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__or2_1
XFILLER_78_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12869__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12081_ net724 _06528_ net1006 VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__a21oi_1
Xhold680 cpuregs\[14\]\[12\] VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold691 cpuregs\[7\]\[10\] VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ cpuregs\[6\]\[19\] cpuregs\[7\]\[19\] net684 VGND VGND VPWR VPWR _05713_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12333__A2 net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12983_ net1518 net340 net447 VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__mux2_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1380 genblk2.pcpi_div.quotient\[3\] VGND VGND VPWR VPWR net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1391 _01117_ VGND VGND VPWR VPWR net2705 sky130_fd_sc_hd__dlygate4sd3_1
X_14722_ clknet_leaf_142_clk net2965 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11934_ net866 _06320_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__and3_1
XFILLER_72_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06785__A net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14775__Q genblk2.pcpi_div.pcpi_rd\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14653_ clknet_leaf_153_clk _01038_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11865_ genblk2.pcpi_div.divisor\[8\] _06305_ genblk2.pcpi_div.dividend\[8\] VGND
+ VGND VPWR VPWR _06336_ sky130_fd_sc_hd__or3b_1
XANTENNA_output106_A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13604_ clknet_leaf_184_clk _00059_ VGND VGND VPWR VPWR cpuregs\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_10816_ net809 _05502_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__or2_1
XFILLER_158_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11796_ genblk2.pcpi_div.divisor\[24\] genblk2.pcpi_div.dividend\[24\] VGND VGND
+ VPWR VPWR _06267_ sky130_fd_sc_hd__and2b_1
X_14584_ clknet_leaf_117_clk _00970_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07276__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13535_ net344 net1433 net416 VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__mux2_1
XFILLER_41_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10747_ cpuregs\[17\]\[11\] net625 net607 _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__o211a_1
XFILLER_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13466_ net2080 net356 net424 VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__mux2_1
X_10678_ net780 _05359_ _05368_ net777 VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__o211a_1
XANTENNA__09100__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15205_ clknet_leaf_33_clk _01554_ VGND VGND VPWR VPWR cpuregs\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08225__B1 net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12021__A1 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12417_ net301 net1939 net474 VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__mux2_1
XFILLER_127_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13397_ _05021_ _05023_ _02304_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__a21oi_1
XFILLER_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput207 net1025 VGND VGND VPWR VPWR pcpi_rs1[13] sky130_fd_sc_hd__buf_2
Xoutput218 net1006 VGND VGND VPWR VPWR pcpi_rs1[23] sky130_fd_sc_hd__buf_2
X_15136_ clknet_leaf_43_clk _01488_ VGND VGND VPWR VPWR cpuregs\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xoutput229 net229 VGND VGND VPWR VPWR pcpi_rs1[4] sky130_fd_sc_hd__buf_2
X_12348_ net3019 net745 _06654_ _06655_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__o22a_1
XFILLER_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13557__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15067_ clknet_leaf_104_clk net2470 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_12279_ net174 _04299_ net175 VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__and3b_1
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12324__A2 _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14018_ clknet_leaf_12_clk _00472_ VGND VGND VPWR VPWR cpuregs\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11532__A0 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06840_ mem_do_wdata mem_do_rdata _02442_ _02443_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__o211a_1
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10886__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06771_ net1087 VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__inv_2
XANTENNA__13285__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08510_ genblk1.genblk1.pcpi_mul.next_rs2\[5\] net1098 _03896_ _03898_ VGND VGND
+ VPWR VPWR _03900_ sky130_fd_sc_hd__and4_1
X_09490_ count_instr\[28\] count_instr\[27\] count_instr\[26\] _04352_ VGND VGND VPWR
+ VPWR _04358_ sky130_fd_sc_hd__and4_1
XANTENNA__10638__A2 net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08386__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08239__X net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08161__C1 net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08441_ net306 net2331 net531 VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__mux2_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07303__B _02843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08372_ reg_pc\[11\] reg_pc\[10\] _03780_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07323_ _02863_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__inv_2
XANTENNA__09661__C1 _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13321__A net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07254_ count_instr\[39\] net1130 net1135 count_instr\[7\] VGND VGND VPWR VPWR _02800_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09010__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07185_ _02731_ _02732_ _02733_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout304_A _03849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_A net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10023__B1 net1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10574__A1 net830 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13467__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12371__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1213_A net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout401 _04293_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__buf_4
Xfanout412 _02358_ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_2
Xfanout423 net426 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11523__A0 mem_rdata_q\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout434 _02128_ VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__buf_4
Xfanout445 net446 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout673_A net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07727__C1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 _02119_ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__buf_4
Xfanout467 net468 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_4
X_09826_ _04437_ _04600_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__nor2_1
Xfanout478 _04292_ VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1001_X net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout489 _04287_ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07742__A2 net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09757_ _04527_ _04546_ _04535_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout840_A _03136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06969_ _02542_ _02543_ _02547_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout938_A net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06950__B1 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11715__S net376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08708_ genblk1.genblk1.pcpi_mul.rd\[35\] genblk1.genblk1.pcpi_mul.next_rs2\[36\]
+ net1098 VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__nand3_1
XANTENNA__08296__S net925 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09688_ _04463_ _04467_ _04476_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_159_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08639_ genblk1.genblk1.pcpi_mul.next_rs2\[25\] net1103 _04006_ _04008_ VGND VGND
+ VPWR VPWR _04009_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout726_X net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07213__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11039__C1 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11650_ net3044 net11 net546 VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__mux2_1
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10601_ cpuregs\[9\]\[7\] net630 net609 _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__o211a_1
XANTENNA__07258__A1 net1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11581_ net2912 net740 _06176_ is_sb_sh_sw VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__a22o_1
XFILLER_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07258__B2 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11054__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12546__S net390 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13320_ _04920_ _02236_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__xnor2_1
X_10532_ _05225_ _05226_ net802 VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__mux2_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13251_ reg_pc\[6\] net565 _02174_ _02176_ net392 VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__a2111oi_1
X_10463_ cpuregs\[25\]\[0\] net634 net611 _05162_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_40_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12202_ net749 _06593_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__nor2_1
X_13182_ net1777 net337 net428 VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__mux2_1
XFILLER_136_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10394_ net1174 _05098_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__or2_1
XFILLER_124_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12133_ net993 _06567_ _02507_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07430__A1 net1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13503__A1 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12064_ _02359_ genblk2.pcpi_div.dividend\[20\] _06363_ VGND VGND VPWR VPWR _06514_
+ sky130_fd_sc_hd__a21bo_1
XANTENNA__11514__A0 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11015_ cpuregs\[24\]\[18\] net648 VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__or2_1
XANTENNA__07194__B1 _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10722__D1 net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input22_X net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout990 _02364_ VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09590__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13267__B1 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output223_A net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13406__A net570 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12966_ net279 net2525 net453 VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__mux2_1
XFILLER_46_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ clknet_leaf_162_clk _01090_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11917_ genblk2.pcpi_div.divisor\[30\] _02389_ _06387_ VGND VGND VPWR VPWR _06388_
+ sky130_fd_sc_hd__o21ai_1
X_12897_ net585 net2444 net457 VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_61_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14636_ clknet_leaf_169_clk _01021_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_11848_ genblk2.pcpi_div.divisor\[1\] genblk2.pcpi_div.dividend\[1\] VGND VGND VPWR
+ VPWR _06319_ sky130_fd_sc_hd__and2b_1
XANTENNA__08934__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11045__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10765__A net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14567_ clknet_leaf_31_clk _00953_ VGND VGND VPWR VPWR cpuregs\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11779_ net33 net268 net1234 VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__and3b_1
XFILLER_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13518_ net1621 net282 net421 VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__mux2_1
X_14498_ clknet_leaf_93_clk _00887_ VGND VGND VPWR VPWR instr_sra sky130_fd_sc_hd__dfxtp_1
Xclkload11 clknet_4_11_0_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinv_8
Xclkload22 clknet_leaf_196_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__bufinv_16
X_13449_ net994 net756 net558 _02328_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__o211a_1
Xclkload33 clknet_leaf_186_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__inv_8
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload44 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__clkinv_2
XFILLER_133_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload55 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__10005__B1 net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12545__A2 net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload66 clknet_leaf_167_clk VGND VGND VPWR VPWR clkload66/Y sky130_fd_sc_hd__bufinv_16
Xclkload77 clknet_leaf_160_clk VGND VGND VPWR VPWR clkload77/Y sky130_fd_sc_hd__inv_12
XANTENNA__10556__B2 net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload88 clknet_leaf_139_clk VGND VGND VPWR VPWR clkload88/Y sky130_fd_sc_hd__inv_6
XANTENNA__11596__A mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload99 clknet_leaf_34_clk VGND VGND VPWR VPWR clkload99/Y sky130_fd_sc_hd__inv_8
X_15119_ clknet_leaf_24_clk _01471_ VGND VGND VPWR VPWR cpuregs\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_08990_ latched_rd\[2\] latched_rd\[4\] latched_rd\[3\] VGND VGND VPWR VPWR _04272_
+ sky130_fd_sc_hd__or3b_1
XFILLER_134_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07972__A2 net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07941_ instr_and instr_andi VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__nor2_2
X_07872_ instr_bne is_slti_blt_slt VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09611_ reg_pc\[11\] net875 _04432_ net845 VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__a22o_1
XFILLER_68_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06823_ instr_auipc instr_lui VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__or2_1
XFILLER_84_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09542_ count_instr\[47\] count_instr\[46\] _04387_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__and3_1
X_06754_ genblk2.pcpi_div.running VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__inv_2
XANTENNA__12220__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09005__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07488__A1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09473_ count_instr\[22\] _04344_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_1
XANTENNA__11284__A2 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08424_ _03827_ _03830_ net768 VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__mux2_1
XANTENNA__10492__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07601__X _03124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08355_ reg_out\[8\] alu_out_q\[8\] net1153 VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__mux2_1
XANTENNA__11036__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12366__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout421_A net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13430__B1 net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06872__B net975 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07306_ _02846_ _02847_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__nand2_1
Xclkload5 clknet_4_5_0_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_8
XFILLER_20_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ reg_out\[20\] reg_next_pc\[20\] net926 VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__mux2_1
XANTENNA__11992__B1 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07237_ count_instr\[38\] net1130 net1139 count_cycle\[38\] VGND VGND VPWR VPWR _02784_
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1049_X net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07168_ net23 net130 _02695_ net10 _02718_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout790_A net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13197__S net430 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07099_ genblk2.pcpi_div.dividend\[26\] net1122 _02657_ net948 VGND VGND VPWR VPWR
+ _02659_ sky130_fd_sc_hd__a31oi_1
XFILLER_121_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1207 _02378_ VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__clkbuf_2
Xfanout1218 net1222 VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__clkbuf_2
Xfanout1229 net1230 VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout676_X net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07176__B1 net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout275 _06403_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout286 net288 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout297 _03852_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
X_09809_ _04573_ _04595_ _04594_ _04580_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12820_ net315 net2016 net465 VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__mux2_1
XANTENNA__09423__B net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12751_ net1550 net903 _02109_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__a21o_1
XFILLER_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_81_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_8
X_11702_ net1909 net330 net373 VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__mux2_1
XANTENNA__10483__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15470_ clknet_leaf_20_clk _01806_ VGND VGND VPWR VPWR cpuregs\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12682_ net1194 net2915 net885 net2978 net711 VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__a221o_1
X_14421_ clknet_leaf_76_clk alu_out\[21\] VGND VGND VPWR VPWR alu_out_q\[21\] sky130_fd_sc_hd__dfxtp_1
X_11633_ mem_rdata_q\[4\] mem_rdata_q\[5\] mem_rdata_q\[6\] mem_rdata_q\[3\] VGND
+ VGND VPWR VPWR _06218_ sky130_fd_sc_hd__or4b_1
XANTENNA__07878__B net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14352_ clknet_leaf_109_clk _00774_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_11564_ net2778 net561 _06178_ _06183_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__a22o_1
XANTENNA__10786__A1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11983__B1 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13303_ _04927_ _02221_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__xnor2_1
X_10515_ cpuregs\[4\]\[5\] net676 VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__or2_1
X_11495_ pcpi_timeout_counter\[2\] pcpi_timeout_counter\[1\] pcpi_timeout_counter\[0\]
+ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__or3_1
X_14283_ clknet_leaf_96_clk _00737_ VGND VGND VPWR VPWR count_cycle\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07894__A net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13234_ reg_pc\[4\] net565 net557 _02160_ net392 VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__a221o_1
X_10446_ cpuregs\[10\]\[0\] net684 VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__or2_1
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10377_ genblk2.pcpi_div.pcpi_wait_q genblk2.pcpi_div.pcpi_wait VGND VGND VPWR VPWR
+ _05082_ sky130_fd_sc_hd__and2b_2
X_13165_ _04275_ _02127_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__nor2_1
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12116_ net725 _06558_ net997 VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__a21oi_1
X_13096_ net283 net1917 net442 VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__mux2_1
XFILLER_105_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12024__B net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12047_ _06497_ _06499_ net861 VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__mux2_1
XANTENNA__08929__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11355__S net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13998_ clknet_leaf_36_clk _00452_ VGND VGND VPWR VPWR cpuregs\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07134__A net1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12949_ net346 net2196 net451 VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13570__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10474__B1 net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpicorv32_1308 VGND VGND VPWR VPWR picorv32_1308/HI trace_data[30] sky130_fd_sc_hd__conb_1
XFILLER_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14619_ clknet_leaf_107_clk _01005_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07890__A1 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15599_ clknet_leaf_182_clk _01935_ VGND VGND VPWR VPWR cpuregs\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__Y _02693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08140_ _03323_ _03630_ _03405_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_99_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09631__A2 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08071_ _03341_ net932 net928 _03343_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__a221o_1
Xclkload100 clknet_leaf_35_clk VGND VGND VPWR VPWR clkload100/Y sky130_fd_sc_hd__clkinv_4
XFILLER_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload111 clknet_leaf_46_clk VGND VGND VPWR VPWR clkload111/Y sky130_fd_sc_hd__inv_6
Xclkload122 clknet_leaf_51_clk VGND VGND VPWR VPWR clkload122/Y sky130_fd_sc_hd__inv_8
XFILLER_128_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12914__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload133 clknet_leaf_66_clk VGND VGND VPWR VPWR clkload133/Y sky130_fd_sc_hd__clkinv_4
X_07022_ genblk2.pcpi_div.quotient\[14\] _02587_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__or2_1
XANTENNA__12518__A2 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload144 clknet_leaf_127_clk VGND VGND VPWR VPWR clkload144/X sky130_fd_sc_hd__clkbuf_8
Xclkload155 clknet_leaf_115_clk VGND VGND VPWR VPWR clkload155/Y sky130_fd_sc_hd__clkinv_4
Xclkload166 clknet_leaf_84_clk VGND VGND VPWR VPWR clkload166/Y sky130_fd_sc_hd__inv_6
XANTENNA__10529__A1 net790 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload177 clknet_leaf_97_clk VGND VGND VPWR VPWR clkload177/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08198__A2 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07309__A net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08973_ net1389 _04263_ net945 VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__mux2_1
Xhold17 genblk1.genblk1.pcpi_mul.next_rs1\[14\] VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _03272_ _03439_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__a21oi_1
Xhold28 cpuregs\[26\]\[20\] VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 instr_ecall_ebreak VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07855_ _03369_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__and2_1
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout371_A net372 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout469_A net470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06806_ net2515 VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__inv_2
X_07786_ net1174 net1042 VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__nor2_1
XFILLER_43_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09525_ count_instr\[40\] _04377_ count_instr\[41\] VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a21o_1
XFILLER_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12454__B2 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13480__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10465__B1 net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09456_ net1228 _04334_ _04335_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__and3_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07330__B1 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08407_ reg_pc\[18\] _03813_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout424_X net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A _03143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09387_ net2017 net311 net401 VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__mux2_1
XANTENNA__13403__B1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout1166_X net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08338_ net573 net2440 net531 VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__mux2_1
XFILLER_165_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08269_ net1028 _03718_ net980 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__mux2_1
XANTENNA__12824__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10300_ decoded_imm\[20\] net1010 VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__or2_1
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11280_ cpuregs\[28\]\[25\] cpuregs\[29\]\[25\] net706 VGND VGND VPWR VPWR _05955_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout793_X net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10231_ decoded_imm\[7\] net1035 VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__and2_1
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11667__C net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10162_ _04871_ _04872_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_167_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_X net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1004 net1005 VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__buf_2
XANTENNA__07875__A_N net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09138__A1 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1015 net212 VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__buf_4
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1026 net1027 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1037 net232 VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__buf_2
X_14970_ clknet_leaf_146_clk _01322_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10093_ count_cycle\[35\] _04826_ net1206 VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1048 net1049 VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__clkbuf_4
Xfanout1059 mem_wordsize\[1\] VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__buf_4
XANTENNA__12142__B1 net372 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07653__S net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13921_ clknet_leaf_14_clk _00375_ VGND VGND VPWR VPWR cpuregs\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13852_ clknet_leaf_197_clk _00306_ VGND VGND VPWR VPWR cpuregs\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12803_ net543 net2064 net464 VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__mux2_1
XFILLER_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11248__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13783_ clknet_leaf_181_clk _00237_ VGND VGND VPWR VPWR cpuregs\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_54_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
X_10995_ net1160 net855 _05676_ _05677_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__a22o_1
X_15522_ clknet_leaf_86_clk _01858_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dfxtp_1
XANTENNA__10456__B1 net611 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12734_ _02408_ net911 VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__nor2_1
XANTENNA__08337__X _03761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14783__Q genblk2.pcpi_div.pcpi_rd\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15453_ clknet_leaf_59_clk _01792_ VGND VGND VPWR VPWR cpuregs\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12665_ genblk1.genblk1.pcpi_mul.mul_waiting net1237 net1157 VGND VGND VPWR VPWR
+ _02082_ sky130_fd_sc_hd__and3_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14404_ clknet_leaf_134_clk alu_out\[4\] VGND VGND VPWR VPWR alu_out_q\[4\] sky130_fd_sc_hd__dfxtp_1
X_11616_ mem_rdata_q\[25\] mem_rdata_q\[24\] VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__nor2_1
X_15384_ clknet_leaf_12_clk _01723_ VGND VGND VPWR VPWR cpuregs\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12596_ net309 net2027 net468 VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14335_ clknet_leaf_176_clk _06722_ VGND VGND VPWR VPWR reg_out\[15\] sky130_fd_sc_hd__dfxtp_1
X_11547_ net27 net28 net29 VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__nand3b_1
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold509 cpuregs\[25\]\[7\] VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14266_ clknet_leaf_122_clk _00720_ VGND VGND VPWR VPWR count_cycle\[11\] sky130_fd_sc_hd__dfxtp_1
X_11478_ net1084 _05076_ net857 VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13217_ _02383_ _02402_ net755 VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__mux2_1
X_10429_ is_beq_bne_blt_bge_bltu_bgeu _03457_ _04881_ _05124_ _05131_ VGND VGND VPWR
+ VPWR _00776_ sky130_fd_sc_hd__a41o_1
X_14197_ clknet_leaf_133_clk _00651_ VGND VGND VPWR VPWR reg_pc\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13148_ net1615 net341 net431 VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13565__S net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13079_ net349 net1733 net439 VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__mux2_1
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12133__B1 _02507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1209 cpuregs\[18\]\[1\] VGND VGND VPWR VPWR net2523 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__B mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07640_ net819 _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__or2_1
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07571_ genblk1.genblk1.pcpi_mul.pcpi_rd\[28\] genblk2.pcpi_div.pcpi_rd\[28\] net1112
+ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__mux2_1
XANTENNA__11239__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12909__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
X_09310_ net1505 net350 net479 VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__mux2_1
XANTENNA__10447__B1 net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07799__A net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08394__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09241_ net1548 net354 net489 VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__mux2_1
XANTENNA__13313__B _05563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09172_ net521 net1819 net496 VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__mux2_1
X_08123_ _03402_ _03619_ net1144 VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07615__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ _03288_ _03301_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__nand2_1
XANTENNA__07738__S net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07005_ genblk2.pcpi_div.dividend\[12\] _02572_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1126_A genblk2.pcpi_div.outsign VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11175__B2 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13475__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08591__A2 net1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08956_ genblk1.genblk1.pcpi_mul.rd\[16\] genblk1.genblk1.pcpi_mul.rd\[48\] net954
+ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__mux2_1
XANTENNA__06878__A _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1710 instr_xori VGND VGND VPWR VPWR net3024 sky130_fd_sc_hd__dlygate4sd3_1
X_07907_ _02392_ net228 _03278_ _03423_ _03420_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a221o_1
Xhold1721 genblk1.genblk1.pcpi_mul.next_rs2\[38\] VGND VGND VPWR VPWR net3035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11478__A2 _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1732 genblk1.genblk1.pcpi_mul.next_rs2\[50\] VGND VGND VPWR VPWR net3046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1743 instr_rdcycle VGND VGND VPWR VPWR net3057 sky130_fd_sc_hd__dlygate4sd3_1
X_08887_ _04217_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout374_X net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1754 genblk1.genblk1.pcpi_mul.next_rs1\[24\] VGND VGND VPWR VPWR net3068 sky130_fd_sc_hd__dlygate4sd3_1
X_07838_ _03351_ _03354_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__or2_1
XFILLER_84_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11008__B net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_A net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07769_ net1163 net1024 VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__nand2_1
XANTENNA__09828__C1 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12819__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_X net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_123_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09508_ _02374_ _04367_ _04369_ net1206 VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_140_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10780_ cpuregs\[20\]\[12\] cpuregs\[21\]\[12\] net646 VGND VGND VPWR VPWR _05468_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09439_ count_instr\[11\] _04323_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout806_X net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08317__B _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12450_ genblk2.pcpi_div.divisor\[35\] _06682_ net868 VGND VGND VPWR VPWR _06683_
+ sky130_fd_sc_hd__mux2_1
X_11401_ cpuregs\[6\]\[29\] cpuregs\[7\]\[29\] net706 VGND VGND VPWR VPWR _06072_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07606__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12554__S net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ net1432 net310 net362 VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14120_ clknet_leaf_58_clk _00574_ VGND VGND VPWR VPWR cpuregs\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10610__B1 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11332_ cpuregs\[2\]\[27\] cpuregs\[3\]\[27\] net692 VGND VGND VPWR VPWR _06005_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14051_ clknet_leaf_13_clk _00505_ VGND VGND VPWR VPWR cpuregs\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11263_ cpuregs\[12\]\[25\] cpuregs\[13\]\[25\] net703 VGND VGND VPWR VPWR _05938_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13002_ _04272_ _04275_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__or2_1
XFILLER_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10214_ _04916_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__nor2_1
XANTENNA__08031__A1 net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11194_ cpuregs\[19\]\[23\] net630 net595 VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__o21a_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10145_ _04860_ _04861_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__nor2_1
XANTENNA__07891__B net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06788__A net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07236__X _02783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14778__Q genblk2.pcpi_div.pcpi_rd\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10076_ _04816_ _04817_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__nor2_1
X_14953_ clknet_leaf_48_clk _01305_ VGND VGND VPWR VPWR cpuregs\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ clknet_leaf_32_clk _00358_ VGND VGND VPWR VPWR cpuregs\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14884_ clknet_leaf_72_clk _01236_ VGND VGND VPWR VPWR cpuregs\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13835_ clknet_leaf_68_clk _00289_ VGND VGND VPWR VPWR cpuregs\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_27_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_44_950 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13414__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13766_ clknet_leaf_35_clk _00220_ VGND VGND VPWR VPWR cpuregs\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_10978_ cpuregs\[16\]\[17\] net647 VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__or2_1
XANTENNA__09103__S net505 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15505_ clknet_leaf_172_clk _01841_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dfxtp_1
X_12717_ net1192 net1354 net2520 net883 _02092_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__a221o_1
X_13697_ clknet_leaf_146_clk _00151_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_15436_ clknet_leaf_192_clk _01775_ VGND VGND VPWR VPWR cpuregs\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08942__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ net2923 net899 _02073_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__a21o_1
X_15367_ clknet_leaf_17_clk _01706_ VGND VGND VPWR VPWR cpuregs\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12579_ net538 net2304 net468 VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__mux2_1
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14318_ clknet_leaf_93_clk _00772_ VGND VGND VPWR VPWR count_cycle\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10601__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15298_ clknet_leaf_99_clk _01639_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.instr_mul
+ sky130_fd_sc_hd__dfxtp_1
Xhold306 cpuregs\[31\]\[3\] VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 cpuregs\[10\]\[9\] VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 net137 VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold339 cpuregs\[21\]\[21\] VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ clknet_leaf_68_clk _00703_ VGND VGND VPWR VPWR reg_next_pc\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout808 _03143_ VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__buf_2
XANTENNA__10904__A1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout819 net821 VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__buf_4
X_08810_ _04153_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__inv_2
XANTENNA__08389__S net529 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09790_ net1183 _04434_ _04578_ _02489_ net846 VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__o221a_1
Xhold1006 cpuregs\[2\]\[1\] VGND VGND VPWR VPWR net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 cpuregs\[18\]\[24\] VGND VGND VPWR VPWR net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _04094_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__inv_2
Xhold1028 cpuregs\[9\]\[30\] VGND VGND VPWR VPWR net2342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1039 cpuregs\[5\]\[27\] VGND VGND VPWR VPWR net2353 sky130_fd_sc_hd__dlygate4sd3_1
X_08672_ _04034_ _04036_ _04029_ _04032_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__a211o_1
XFILLER_39_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07623_ cpuregs\[6\]\[2\] cpuregs\[7\]\[2\] net700 VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07554_ genblk1.genblk1.pcpi_mul.pcpi_rd\[27\] genblk2.pcpi_div.pcpi_rd\[27\] net1113
+ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_81_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09013__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07485_ genblk1.genblk1.pcpi_mul.pcpi_rd\[22\] genblk2.pcpi_div.pcpi_rd\[22\] net1112
+ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout334_A _03815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09224_ net1654 net295 net494 VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__mux2_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12374__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09155_ net1523 net307 net502 VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout501_A net503 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06880__B net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11396__A1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08106_ _03465_ _03604_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__nor2_1
XFILLER_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09086_ net1416 net302 net511 VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__mux2_1
X_08037_ _03351_ _03522_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__nand2_1
XFILLER_162_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1031_X net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold840 cpuregs\[13\]\[25\] VGND VGND VPWR VPWR net2154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1129_X net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold851 cpuregs\[15\]\[9\] VGND VGND VPWR VPWR net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 cpuregs\[19\]\[15\] VGND VGND VPWR VPWR net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 cpuregs\[2\]\[12\] VGND VGND VPWR VPWR net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 cpuregs\[9\]\[13\] VGND VGND VPWR VPWR net2198 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08440__X _03844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout491_X net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold895 cpuregs\[3\]\[24\] VGND VGND VPWR VPWR net2209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout589_X net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A _02432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09988_ _04756_ _04759_ net1186 _04451_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08299__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08939_ net1861 _04246_ net943 VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1540 genblk2.pcpi_div.quotient\[27\] VGND VGND VPWR VPWR net2854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 count_instr\[62\] VGND VGND VPWR VPWR net2865 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1562 genblk2.pcpi_div.divisor\[23\] VGND VGND VPWR VPWR net2876 sky130_fd_sc_hd__dlygate4sd3_1
X_11950_ _06315_ _06324_ _06323_ _06316_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_142_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1573 genblk2.pcpi_div.divisor\[6\] VGND VGND VPWR VPWR net2887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1584 genblk2.pcpi_div.divisor\[3\] VGND VGND VPWR VPWR net2898 sky130_fd_sc_hd__dlygate4sd3_1
X_10901_ cpuregs\[25\]\[15\] net617 net603 _05585_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__o211a_1
Xhold1595 genblk2.pcpi_div.quotient_msk\[7\] VGND VGND VPWR VPWR net2909 sky130_fd_sc_hd__dlygate4sd3_1
X_11881_ _06295_ _06296_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__nand2b_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12549__S net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13620_ clknet_leaf_72_clk _00075_ VGND VGND VPWR VPWR cpuregs\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_10832_ cpuregs\[22\]\[13\] cpuregs\[23\]\[13\] net651 VGND VGND VPWR VPWR _05519_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11084__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13551_ net283 net2045 net417 VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__mux2_1
X_10763_ cpuregs\[10\]\[11\] net653 VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__or2_1
XFILLER_160_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12502_ net1162 net715 _05107_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__or3b_1
X_13482_ net1473 net295 net425 VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__mux2_1
XFILLER_157_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10694_ net827 _05380_ _05382_ _05384_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__a211o_1
XFILLER_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15221_ clknet_leaf_85_clk _00010_ VGND VGND VPWR VPWR cpu_state\[6\] sky130_fd_sc_hd__dfxtp_1
X_12433_ genblk1.genblk1.pcpi_mul.mul_counter\[4\] _06669_ VGND VGND VPWR VPWR _06670_
+ sky130_fd_sc_hd__or2_1
XFILLER_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12584__A0 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15152_ clknet_leaf_89_clk _01501_ VGND VGND VPWR VPWR mem_rdata_q\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12364_ net1411 net540 net361 VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__mux2_1
XFILLER_165_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10595__C1 net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14103_ clknet_leaf_185_clk _00557_ VGND VGND VPWR VPWR cpuregs\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11315_ cpuregs\[27\]\[26\] net642 net601 _05988_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__o211a_1
XFILLER_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15083_ clknet_leaf_48_clk _01435_ VGND VGND VPWR VPWR cpuregs\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12295_ mem_rdata_q\[26\] net559 _06626_ net532 VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__a211o_1
XANTENNA__11139__A1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08004__A1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14034_ clknet_leaf_23_clk _00488_ VGND VGND VPWR VPWR cpuregs\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08004__B2 net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11246_ cpuregs\[9\]\[24\] net634 net611 _05921_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__o211a_1
XANTENNA__12887__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output253_A net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06789__Y _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10532__S net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11177_ net774 _05846_ _05854_ _05838_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__a31oi_4
X_10128_ net2701 _04848_ net1228 VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12639__B2 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10059_ count_cycle\[23\] _04804_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__and2_1
X_14936_ clknet_leaf_5_clk _01288_ VGND VGND VPWR VPWR cpuregs\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08937__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14867_ clknet_leaf_6_clk _01219_ VGND VGND VPWR VPWR cpuregs\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12459__S net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13818_ clknet_leaf_198_clk _00272_ VGND VGND VPWR VPWR cpuregs\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13064__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14798_ clknet_leaf_81_clk _01150_ VGND VGND VPWR VPWR decoded_imm\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11075__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13749_ clknet_leaf_19_clk _00203_ VGND VGND VPWR VPWR cpuregs\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10822__B1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07270_ count_instr\[40\] net1131 net1136 count_instr\[8\] VGND VGND VPWR VPWR _02815_
+ sky130_fd_sc_hd__a22o_1
X_15419_ clknet_leaf_16_clk _01758_ VGND VGND VPWR VPWR cpuregs\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13367__A2 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08243__A1 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold103 cpuregs\[28\]\[28\] VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 cpuregs\[30\]\[30\] VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 net56 VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 genblk1.genblk1.pcpi_mul.next_rs1\[29\] VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12922__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold147 net46 VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold158 cpuregs\[12\]\[8\] VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _04443_ _04672_ _04444_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__a21oi_1
Xhold169 cpuregs\[15\]\[11\] VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 net606 VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__clkbuf_4
Xfanout616 _03148_ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout627 net628 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__buf_2
X_09842_ net1182 _04438_ net847 VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout638 net639 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_2
XFILLER_58_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout649 net654 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11550__A1 net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09008__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09773_ net984 _04561_ _04562_ _04559_ _04560_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a32o_1
X_06985_ genblk2.pcpi_div.dividend\[10\] _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout284_A _03870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08724_ _04078_ _04080_ _04073_ _04076_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__a211o_1
XFILLER_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11302__A1 net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_clk_X clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ net902 _04020_ _04022_ net2683 net1212 VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__a32o_1
XANTENNA__12369__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11273__S net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_A net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout549_A net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07606_ net25 net939 net937 VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13055__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08586_ genblk1.genblk1.pcpi_mul.rd\[16\] genblk1.genblk1.pcpi_mul.rdx\[16\] VGND
+ VGND VPWR VPWR _03964_ sky130_fd_sc_hd__or2_1
X_07537_ net359 _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__nor2_1
XFILLER_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10813__B1 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1079_X net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07468_ net358 _02999_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__nor2_1
XFILLER_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09207_ net1430 net405 net493 VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__mux2_1
XFILLER_22_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout504_X net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07399_ genblk1.genblk1.pcpi_mul.pcpi_rd\[16\] genblk2.pcpi_div.pcpi_rd\[16\] net1111
+ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__mux2_1
XANTENNA__11369__B2 net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09138_ net1603 net524 net500 VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__mux2_1
XANTENNA__08234__A1 net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ net1607 net523 net509 VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__mux2_1
XFILLER_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12832__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10592__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12318__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11100_ cpuregs\[9\]\[20\] net622 net605 _05779_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__o211a_1
XFILLER_151_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09707__A decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12080_ net1008 _06523_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__or2_1
XANTENNA__11956__B net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold670 cpuregs\[9\]\[11\] VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold681 cpuregs\[20\]\[31\] VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 cpuregs\[7\]\[12\] VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net244 net855 _05711_ _05712_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__a22o_1
XFILLER_150_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11972__A net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12982_ net1632 net343 net447 VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__mux2_1
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1370 net189 VGND VGND VPWR VPWR net2684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07661__S net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input12_A mem_rdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1381 _06582_ VGND VGND VPWR VPWR net2695 sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ clknet_leaf_142_clk net2580 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11933_ genblk2.pcpi_div.divisor\[0\] genblk2.pcpi_div.dividend\[0\] VGND VGND VPWR
+ VPWR _06404_ sky130_fd_sc_hd__nand2b_1
Xhold1392 genblk1.genblk1.pcpi_mul.rdx\[24\] VGND VGND VPWR VPWR net2706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11183__S net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14652_ clknet_leaf_155_clk _01037_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13046__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11864_ _02361_ genblk2.pcpi_div.dividend\[8\] _06334_ VGND VGND VPWR VPWR _06335_
+ sky130_fd_sc_hd__a21o_1
X_13603_ clknet_leaf_183_clk _00058_ VGND VGND VPWR VPWR cpuregs\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10815_ cpuregs\[14\]\[13\] cpuregs\[15\]\[13\] net652 VGND VGND VPWR VPWR _05502_
+ sky130_fd_sc_hd__mux2_1
X_14583_ clknet_leaf_69_clk _00969_ VGND VGND VPWR VPWR latched_rd\[4\] sky130_fd_sc_hd__dfxtp_2
X_11795_ _06264_ _06265_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__or2_1
XFILLER_41_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ net348 net2070 net415 VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10746_ cpuregs\[16\]\[11\] net665 VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__or2_1
XFILLER_159_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13465_ net1415 net404 net424 VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__mux2_1
XFILLER_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10677_ net789 _05363_ _05365_ _05367_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__or4_1
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15204_ clknet_leaf_22_clk _01553_ VGND VGND VPWR VPWR cpuregs\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12416_ net306 net2363 net473 VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__mux2_1
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13396_ _05021_ _05023_ net959 VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__o21ai_1
Xoutput208 net1023 VGND VGND VPWR VPWR pcpi_rs1[14] sky130_fd_sc_hd__buf_2
X_15135_ clknet_leaf_13_clk _01487_ VGND VGND VPWR VPWR cpuregs\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12347_ net1151 decoded_imm_j\[2\] _06617_ mem_rdata_q\[9\] net733 VGND VGND VPWR
+ VPWR _06655_ sky130_fd_sc_hd__a221o_1
Xoutput219 net1005 VGND VGND VPWR VPWR pcpi_rs1[24] sky130_fd_sc_hd__buf_2
XFILLER_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output80_A net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07984__B1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15066_ clknet_leaf_104_clk _01418_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_12278_ net175 net174 _04299_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__and3b_1
XFILLER_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09725__A1 net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14017_ clknet_leaf_42_clk _00471_ VGND VGND VPWR VPWR cpuregs\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11229_ cpuregs\[17\]\[24\] net640 net614 _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__o211a_1
XFILLER_68_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13573__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06770_ net1227 VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__inv_2
XANTENNA__07571__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14919_ clknet_leaf_113_clk _01271_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08440_ _03840_ _03843_ net768 VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__mux2_2
XANTENNA__13037__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08371_ reg_pc\[11\] reg_pc\[10\] _03780_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__and3_1
XANTENNA__12917__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07322_ reg_pc\[10\] decoded_imm\[10\] _02847_ _02862_ VGND VGND VPWR VPWR _02863_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12260__A2 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08255__X net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07253_ net30 net130 _02695_ net16 _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__a221o_1
XANTENNA__10437__S net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07184_ _02732_ _02733_ _02731_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__a21o_1
XANTENNA__08216__A1 net1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1039_A net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout402 _04293_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_4
Xfanout413 _02358_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_4
XANTENNA__09716__B2 net852 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout424 net426 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_4
Xfanout435 net436 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1206_A net1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout446 _02124_ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12720__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A mem_rdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09825_ _04437_ _04600_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__and2_1
Xfanout457 _02119_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__buf_4
Xfanout468 _02051_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__buf_4
XFILLER_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout666_A net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout479 net483 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout287_X net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13483__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09756_ _04535_ _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__nand2_1
X_06968_ net951 _02545_ _02546_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__or3_1
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08707_ net894 _04064_ _04066_ net2703 net1202 VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__a32o_1
X_09687_ _04482_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__nor2_1
X_06899_ is_slli_srli_srai _02471_ _02493_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout454_X net454 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__D1 net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08638_ genblk1.genblk1.pcpi_mul.rd\[24\] genblk1.genblk1.pcpi_mul.rdx\[24\] VGND
+ VGND VPWR VPWR _04008_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_159_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10201__A decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08569_ _03941_ _03944_ _03946_ _03948_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__o211a_1
XANTENNA__12827__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06892__Y _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_X net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10600_ cpuregs\[8\]\[7\] net673 VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__or2_1
XFILLER_23_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07258__A2 net1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11580_ net2849 net740 _06183_ _06191_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__a22o_1
XFILLER_120_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12251__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09201__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10531_ cpuregs\[30\]\[5\] cpuregs\[31\]\[5\] net678 VGND VGND VPWR VPWR _05226_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12539__B1 net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13250_ net1045 net754 _02175_ net709 VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__o211a_1
X_10462_ cpuregs\[24\]\[0\] net684 VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__or2_1
XANTENNA__13200__A1 net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout990_X net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ net2863 net274 net2944 VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13181_ net1574 net341 net427 VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__mux2_1
X_10393_ net1180 net1178 net1176 net1177 VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__or4_2
XANTENNA__10565__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12132_ genblk2.pcpi_div.dividend\[30\] net275 _06572_ VGND VGND VPWR VPWR _01039_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12063_ genblk2.pcpi_div.dividend\[20\] _06513_ net269 VGND VGND VPWR VPWR _01029_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07718__B1 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11014_ _05694_ _05695_ net809 VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__mux2_1
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07194__A1 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07194__B2 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout980 net981 VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__buf_4
Xfanout991 _02363_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__buf_4
XANTENNA__06796__A net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input15_X net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12965_ net284 net2456 net453 VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__mux2_1
XANTENNA__13406__B _05964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output216_A net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14704_ clknet_leaf_153_clk _01089_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_11916_ _06263_ _06384_ _06260_ _06262_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_47_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07404__B decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12896_ net588 net2340 net457 VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__mux2_1
X_14635_ clknet_leaf_169_clk _01020_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11847_ genblk2.pcpi_div.dividend\[2\] genblk2.pcpi_div.divisor\[2\] VGND VGND VPWR
+ VPWR _06318_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11641__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13422__A net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14566_ clknet_leaf_37_clk _00952_ VGND VGND VPWR VPWR cpuregs\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11778_ _02417_ _06239_ _06250_ _06251_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__o31ai_1
XANTENNA__12242__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09111__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13517_ net1586 net287 net421 VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__mux2_1
XANTENNA__11213__Y _05890_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10729_ cpuregs\[18\]\[10\] net553 _05418_ net780 VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__o22a_1
XFILLER_119_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14497_ clknet_leaf_95_clk _00886_ VGND VGND VPWR VPWR instr_srl sky130_fd_sc_hd__dfxtp_1
XANTENNA__12038__A net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13448_ net1000 net757 _02336_ _02501_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__o211a_1
Xclkload12 clknet_4_12_0_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_8
XFILLER_139_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload23 clknet_leaf_197_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_6
XANTENNA__08950__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload34 clknet_leaf_187_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__inv_6
XANTENNA__13568__S net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_173_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload45 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__bufinv_16
Xclkload56 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload56/Y sky130_fd_sc_hd__inv_6
Xclkload67 clknet_leaf_169_clk VGND VGND VPWR VPWR clkload67/Y sky130_fd_sc_hd__clkinv_4
X_13379_ _02410_ net760 VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__nand2_1
Xclkload78 clknet_leaf_161_clk VGND VGND VPWR VPWR clkload78/Y sky130_fd_sc_hd__clkinv_8
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11753__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10556__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07957__B1 net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload89 clknet_leaf_140_clk VGND VGND VPWR VPWR clkload89/Y sky130_fd_sc_hd__clkinvlp_4
X_15118_ clknet_leaf_27_clk _01470_ VGND VGND VPWR VPWR cpuregs\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15049_ clknet_leaf_105_clk _01401_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07940_ _02377_ _02384_ net969 VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_188_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07871_ _03382_ _03386_ _03387_ _03388_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_3_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ _03786_ reg_next_pc\[11\] net920 VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__mux2_2
X_06822_ _02423_ _02424_ _02425_ _02426_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13258__A1 net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11269__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09541_ count_instr\[46\] _04387_ count_instr\[47\] VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a21o_1
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06753_ genblk2.pcpi_div.divisor\[8\] VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__inv_2
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11117__A net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09472_ count_instr\[22\] _04344_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__or2_1
X_08423_ _03828_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__nor2_1
XFILLER_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13332__A net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08354_ net524 net2309 net529 VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__mux2_1
XANTENNA__12233__A2 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__S net519 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07305_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload6 clknet_4_6_0_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_16
X_08285_ net1012 _03726_ net981 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__mux2_2
XANTENNA_fanout414_A _02358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09956__S net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07236_ net29 net130 _02695_ net15 _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__a221o_1
XFILLER_165_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13478__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09937__A1 net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11787__A net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12382__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07167_ _02383_ net19 _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_132_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07329__X _02870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07098_ net1122 _02657_ genblk2.pcpi_div.dividend\[26\] VGND VGND VPWR VPWR _02658_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout783_A net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1208 net1209 VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1111_X net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1219 net1221 VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1209_X net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input7_X net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_A net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11726__S net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout276 net277 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_4
Xfanout287 net288 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_2
X_09808_ _04567_ _04582_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__nand2_1
Xfanout298 _03852_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_1
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09739_ net1149 _04526_ _04528_ _04531_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout836_X net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12750_ net1214 net3068 net918 net1003 VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__a22o_1
XFILLER_55_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11701_ net1988 net332 net373 VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__mux2_1
XFILLER_70_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12681_ net1194 net3070 net885 genblk1.genblk1.pcpi_mul.next_rs2\[45\] net711 VGND
+ VGND VPWR VPWR _01351_ sky130_fd_sc_hd__a221o_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14420_ clknet_leaf_77_clk alu_out\[20\] VGND VGND VPWR VPWR alu_out_q\[20\] sky130_fd_sc_hd__dfxtp_1
X_11632_ net1134 net737 _06215_ _06217_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10585__B _05278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14351_ clknet_leaf_87_clk _06740_ VGND VGND VPWR VPWR reg_out\[31\] sky130_fd_sc_hd__dfxtp_1
X_11563_ _02388_ _06179_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__nor2_2
XFILLER_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13302_ decoded_imm\[12\] net1026 _04983_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__a21o_1
X_10514_ cpuregs\[6\]\[5\] cpuregs\[7\]\[5\] net676 VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__mux2_1
X_14282_ clknet_leaf_100_clk _00736_ VGND VGND VPWR VPWR count_cycle\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11494_ genblk2.pcpi_div.pcpi_wait genblk1.genblk1.pcpi_mul.pcpi_wait net267 net1237
+ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__or4bb_1
XFILLER_137_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13233_ net1033 net758 VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__or2_1
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10445_ _05143_ _05144_ net804 VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__mux2_1
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11735__A1 net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12932__B1 decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13164_ net1594 net281 net434 VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__mux2_1
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10376_ _04889_ _05039_ _05077_ _05081_ _04890_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__o41a_1
X_12115_ net1001 net999 _06549_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__or3_2
X_13095_ net286 net2386 net441 VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_15_0_clk_X clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12046_ _06285_ _06359_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07167__A1 _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10540__S net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10171__B1 net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10710__A2 net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09106__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07415__A _02950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13997_ clknet_leaf_50_clk _00451_ VGND VGND VPWR VPWR cpuregs\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07134__B net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12948_ net349 net2024 net452 VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__mux2_1
XANTENNA__08945__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ mem_rdata_q\[16\] net8 net962 VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__mux2_1
XANTENNA__12467__S net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1309 VGND VGND VPWR VPWR picorv32_1309/HI trace_data[31] sky130_fd_sc_hd__conb_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14618_ clknet_leaf_117_clk _01004_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dfxtp_1
XANTENNA__12215__A2 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15598_ clknet_leaf_183_clk _01934_ VGND VGND VPWR VPWR cpuregs\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13384__A2_N _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07150__A net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11423__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14549_ clknet_leaf_179_clk _00935_ VGND VGND VPWR VPWR cpuregs\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10777__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08070_ net968 _03342_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__nor2_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload101 clknet_leaf_36_clk VGND VGND VPWR VPWR clkload101/Y sky130_fd_sc_hd__clkinv_2
Xclkload112 clknet_leaf_47_clk VGND VGND VPWR VPWR clkload112/Y sky130_fd_sc_hd__inv_8
Xclkload123 clknet_leaf_52_clk VGND VGND VPWR VPWR clkload123/Y sky130_fd_sc_hd__clkinv_4
Xclkload134 clknet_leaf_67_clk VGND VGND VPWR VPWR clkload134/X sky130_fd_sc_hd__clkbuf_8
X_07021_ genblk2.pcpi_div.dividend\[15\] _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload145 clknet_leaf_128_clk VGND VGND VPWR VPWR clkload145/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_127_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload156 clknet_leaf_116_clk VGND VGND VPWR VPWR clkload156/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload167 clknet_leaf_85_clk VGND VGND VPWR VPWR clkload167/Y sky130_fd_sc_hd__bufinv_16
Xclkload178 clknet_leaf_98_clk VGND VGND VPWR VPWR clkload178/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__07149__X _02702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08972_ genblk1.genblk1.pcpi_mul.rd\[24\] genblk1.genblk1.pcpi_mul.rd\[56\] net956
+ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__mux2_1
XFILLER_142_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07923_ _02396_ net1004 _03272_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__a31o_1
Xhold18 _01384_ VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 cpuregs\[14\]\[29\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12687__C1 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07854_ _03370_ _03371_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__or2_1
XFILLER_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09016__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06805_ is_sltiu_bltu_sltu VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__inv_2
X_07785_ net1174 net1042 VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__nand2_1
XFILLER_25_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09524_ count_instr\[40\] _04377_ _04379_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__o21a_1
XFILLER_24_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11111__C1 net840 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11662__A0 decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09455_ count_instr\[16\] _04332_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout531_A _03746_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07979__B net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12377__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11281__S net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08406_ reg_out\[18\] alu_out_q\[18\] net1154 VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__mux2_1
X_09386_ net2085 net314 net401 VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__mux2_1
XANTENNA__13403__B2 net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08337_ _03757_ _03760_ net767 VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__mux2_2
XFILLER_165_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout417_X net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_X net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08268_ reg_out\[11\] reg_next_pc\[11\] net920 VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout998_A net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07219_ net28 net130 _02695_ net14 _02766_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__a221o_1
X_08199_ _03371_ _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__nor2_1
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10230_ decoded_imm\[8\] net1033 VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__nand2_2
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout786_X net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10925__C1 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11193__A2 net624 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10161_ net2968 _04869_ net1238 VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__o21ai_1
XFILLER_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12840__S net460 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11544__C_N net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1005 net219 VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__buf_4
XFILLER_0_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1016 net211 VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__buf_4
Xfanout1027 net206 VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__buf_2
XANTENNA__12678__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1038 net231 VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout953_X net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10092_ _04826_ _04827_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__nor2_1
XFILLER_75_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1049 net1050 VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__buf_2
X_13920_ clknet_leaf_8_clk _00374_ VGND VGND VPWR VPWR cpuregs\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13851_ clknet_leaf_196_clk _00305_ VGND VGND VPWR VPWR cpuregs\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11028__Y _05710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12802_ net571 net1881 net465 VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__mux2_1
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13782_ clknet_leaf_180_clk _00236_ VGND VGND VPWR VPWR cpuregs\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10994_ net1078 decoded_imm\[17\] net860 VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__o21a_1
XFILLER_90_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15521_ clknet_leaf_75_clk _01857_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dfxtp_1
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12733_ net1191 net1326 net2197 net884 _02100_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__S net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15452_ clknet_leaf_35_clk _01791_ VGND VGND VPWR VPWR cpuregs\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12664_ net3027 net905 _02081_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__a21o_1
XFILLER_124_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14403_ clknet_leaf_134_clk alu_out\[3\] VGND VGND VPWR VPWR alu_out_q\[3\] sky130_fd_sc_hd__dfxtp_1
X_11615_ mem_rdata_q\[31\] mem_rdata_q\[30\] net746 _06194_ VGND VGND VPWR VPWR _06204_
+ sky130_fd_sc_hd__and4_1
XFILLER_89_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15383_ clknet_leaf_41_clk _01722_ VGND VGND VPWR VPWR cpuregs\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12595_ net314 net2382 net469 VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__mux2_1
XFILLER_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14334_ clknet_leaf_177_clk _06721_ VGND VGND VPWR VPWR reg_out\[14\] sky130_fd_sc_hd__dfxtp_1
X_11546_ net1414 _06170_ net547 VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__mux2_1
XFILLER_51_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08353__X _03774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14265_ clknet_leaf_122_clk _00719_ VGND VGND VPWR VPWR count_cycle\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11477_ net1084 decoded_imm\[31\] VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_94_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13216_ net959 _04956_ _02145_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__and3_1
X_10428_ _05130_ mem_do_rinst _05127_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14196_ clknet_leaf_132_clk _00650_ VGND VGND VPWR VPWR reg_pc\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13147_ net1476 net345 net432 VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__mux2_1
X_10359_ cpuregs\[18\]\[31\] net554 _05064_ net783 VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_55_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ net352 net1833 net439 VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12669__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12133__A1 net993 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11366__S net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12029_ net1021 _06480_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__or2_1
XANTENNA__11593__C mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10144__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10695__A1 net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13581__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07570_ count_cycle\[28\] net973 net843 _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__o211a_1
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09837__B1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09240_ net1749 net405 net489 VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_1_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09171_ net526 net2387 net496 VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__mux2_1
XANTENNA__12925__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08122_ _03330_ _03613_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__nor2_1
XANTENNA__08263__X net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07615__A2 decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08053_ _03379_ net930 _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10445__S net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12226__A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07004_ _02573_ _02574_ _02576_ _02577_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__o22ai_1
XFILLER_134_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11175__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08955_ net2568 _04254_ net943 VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout481_A _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1700 genblk1.genblk1.pcpi_mul.next_rs2\[26\] VGND VGND VPWR VPWR net3014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout579_A _03753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1711 genblk2.pcpi_div.dividend\[12\] VGND VGND VPWR VPWR net3025 sky130_fd_sc_hd__dlygate4sd3_1
X_07906_ _03278_ _03423_ _03420_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__a21oi_1
Xhold1722 instr_lb VGND VGND VPWR VPWR net3036 sky130_fd_sc_hd__dlygate4sd3_1
X_08886_ _04211_ _04214_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__nand2_1
XFILLER_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1733 count_instr\[29\] VGND VGND VPWR VPWR net3047 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1744 genblk2.pcpi_div.dividend\[4\] VGND VGND VPWR VPWR net3058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1755 genblk2.pcpi_div.divisor\[16\] VGND VGND VPWR VPWR net3069 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07000__B1 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10686__A1 net830 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07837_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__inv_2
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout746_A net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13491__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07768_ net1163 net1024 VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__or2_1
XFILLER_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09507_ _04363_ _04368_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__and2_1
XFILLER_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout534_X net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07699_ cpuregs\[22\]\[3\] cpuregs\[23\]\[3\] net674 VGND VGND VPWR VPWR _03219_
+ sky130_fd_sc_hd__mux2_1
XFILLER_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09438_ _04323_ net1226 _04322_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__and3b_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09369_ net1778 net542 net400 VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout701_X net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12835__S net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11400_ net255 net857 _06070_ _06071_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__a22o_1
XANTENNA__07606__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12380_ net2122 net313 net362 VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__mux2_1
XFILLER_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11331_ _06002_ _06003_ net817 VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10355__S net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14050_ clknet_leaf_11_clk _00504_ VGND VGND VPWR VPWR cpuregs\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11262_ cpuregs\[14\]\[25\] cpuregs\[15\]\[25\] net703 VGND VGND VPWR VPWR _05937_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13001_ net2515 net907 VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__and2_1
XFILLER_140_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13560__A0 net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10213_ decoded_imm\[15\] net1020 VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__and2_1
XANTENNA__12570__S net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11193_ cpuregs\[17\]\[23\] net624 net611 _05869_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__o211a_1
X_10144_ net2862 _04858_ net1235 VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__o21ai_1
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10075_ net2747 _04814_ net1236 VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__o21ai_1
X_14952_ clknet_leaf_72_clk _01304_ VGND VGND VPWR VPWR cpuregs\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12666__A2 genblk1.genblk1.pcpi_mul.next_rs2\[32\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ clknet_leaf_47_clk _00357_ VGND VGND VPWR VPWR cpuregs\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14883_ clknet_leaf_47_clk _01235_ VGND VGND VPWR VPWR cpuregs\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_13834_ clknet_leaf_46_clk _00288_ VGND VGND VPWR VPWR cpuregs\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10429__A1 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13414__B _05999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13765_ clknet_leaf_16_clk _00219_ VGND VGND VPWR VPWR cpuregs\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_10977_ _05658_ _05659_ net809 VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__mux2_1
XANTENNA__08098__A2 net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15504_ clknet_leaf_167_clk _01840_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dfxtp_1
X_12716_ genblk1.genblk1.pcpi_mul.mul_waiting net1223 net1034 VGND VGND VPWR VPWR
+ _02092_ sky130_fd_sc_hd__and3_1
X_13696_ clknet_leaf_151_clk _00150_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15435_ clknet_leaf_20_clk _01774_ VGND VGND VPWR VPWR cpuregs\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12647_ net1210 genblk1.genblk1.pcpi_mul.next_rs2\[23\] net918 net249 VGND VGND VPWR
+ VPWR _02073_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07058__B1 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12051__B1 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15366_ clknet_leaf_31_clk _01705_ VGND VGND VPWR VPWR cpuregs\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12578_ net541 net2211 net468 VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__mux2_1
XFILLER_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11529_ mem_rdata_q\[22\] net2423 net742 VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__mux2_1
X_14317_ clknet_leaf_94_clk _00771_ VGND VGND VPWR VPWR count_cycle\[62\] sky130_fd_sc_hd__dfxtp_1
X_15297_ clknet_leaf_56_clk _01638_ VGND VGND VPWR VPWR cpuregs\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold307 cpuregs\[15\]\[30\] VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold318 cpuregs\[30\]\[14\] VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14248_ clknet_leaf_75_clk _00702_ VGND VGND VPWR VPWR reg_next_pc\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold329 cpuregs\[23\]\[6\] VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13576__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14179_ clknet_leaf_109_clk _00633_ VGND VGND VPWR VPWR count_instr\[50\] sky130_fd_sc_hd__dfxtp_1
Xfanout809 net812 VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__buf_4
XFILLER_140_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12106__A1 net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1007 cpuregs\[16\]\[28\] VGND VGND VPWR VPWR net2321 sky130_fd_sc_hd__dlygate4sd3_1
X_08740_ genblk1.genblk1.pcpi_mul.rd\[40\] genblk1.genblk1.pcpi_mul.rdx\[40\] VGND
+ VGND VPWR VPWR _04094_ sky130_fd_sc_hd__nand2_1
Xhold1018 cpuregs\[25\]\[25\] VGND VGND VPWR VPWR net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 cpuregs\[11\]\[22\] VGND VGND VPWR VPWR net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__B1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10668__A1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08671_ genblk1.genblk1.pcpi_mul.rd\[29\] genblk1.genblk1.pcpi_mul.next_rs2\[30\]
+ net1106 VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__nand3_1
XFILLER_94_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07622_ net986 decoded_imm_j\[1\] _03141_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__o21a_2
XFILLER_66_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07553_ count_cycle\[27\] net973 net843 _03078_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__o211a_1
XANTENNA__11078__D1 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07297__B1 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07484_ count_cycle\[22\] net973 net843 _03014_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_17_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11093__B2 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09223_ net1932 net299 net495 VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__mux2_1
XFILLER_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A _03823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_A net1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13340__A _02410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09154_ net1618 net310 net502 VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__mux2_1
XFILLER_147_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3_0_clk_X clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08105_ _03336_ _03603_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__xor2_1
X_09085_ net1666 net305 net511 VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1236_A net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08036_ _03302_ net930 _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__o21ai_1
Xhold830 cpuregs\[17\]\[12\] VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 cpuregs\[3\]\[16\] VGND VGND VPWR VPWR net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__A1 decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap560 _06229_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13486__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold852 cpuregs\[4\]\[22\] VGND VGND VPWR VPWR net2166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net707 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold863 cpuregs\[23\]\[22\] VGND VGND VPWR VPWR net2177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold874 cpuregs\[15\]\[6\] VGND VGND VPWR VPWR net2188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06889__A net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_X net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold885 cpuregs\[29\]\[1\] VGND VGND VPWR VPWR net2199 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold896 cpuregs\[18\]\[13\] VGND VGND VPWR VPWR net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ net1152 _04757_ _04758_ net1186 VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout863_A net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_X net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08938_ genblk1.genblk1.pcpi_mul.rd\[7\] genblk1.genblk1.pcpi_mul.rd\[39\] net954
+ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__mux2_1
Xhold1530 _01069_ VGND VGND VPWR VPWR net2844 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10659__A1 net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1541 count_instr\[59\] VGND VGND VPWR VPWR net2855 sky130_fd_sc_hd__dlygate4sd3_1
X_08869_ net1213 net2917 net901 _04203_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__a22o_1
Xhold1552 genblk2.pcpi_div.quotient_msk\[11\] VGND VGND VPWR VPWR net2866 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1563 genblk2.pcpi_div.quotient\[9\] VGND VGND VPWR VPWR net2877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout749_X net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1574 genblk1.genblk1.pcpi_mul.rd\[19\] VGND VGND VPWR VPWR net2888 sky130_fd_sc_hd__dlygate4sd3_1
X_10900_ cpuregs\[24\]\[15\] net649 VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__or2_1
Xhold1585 _01108_ VGND VGND VPWR VPWR net2899 sky130_fd_sc_hd__dlygate4sd3_1
X_11880_ _06294_ _06350_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__or2_1
Xhold1596 reg_next_pc\[24\] VGND VGND VPWR VPWR net2910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09204__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10831_ cpuregs\[20\]\[13\] cpuregs\[21\]\[13\] net651 VGND VGND VPWR VPWR _05518_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_64_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout916_X net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13550_ net286 net2620 net418 VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__mux2_1
XANTENNA__15730__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10762_ cpuregs\[9\]\[11\] net628 net607 _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__o211a_1
XFILLER_25_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12501_ _01995_ _01996_ net2623 net386 VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13481_ net1554 net299 net425 VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__mux2_1
X_10693_ cpuregs\[18\]\[9\] net553 _05383_ net780 VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__o22a_1
X_15220_ clknet_leaf_88_clk _00009_ VGND VGND VPWR VPWR cpu_state\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12432_ net917 _06668_ _06669_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__or3b_1
XFILLER_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15151_ clknet_leaf_90_clk _01500_ VGND VGND VPWR VPWR mem_rdata_q\[2\] sky130_fd_sc_hd__dfxtp_1
X_12363_ net1372 net543 net361 VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__mux2_1
XFILLER_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14102_ clknet_leaf_185_clk _00556_ VGND VGND VPWR VPWR cpuregs\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11314_ cpuregs\[26\]\[26\] net703 VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__or2_1
XFILLER_126_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15082_ clknet_leaf_37_clk _01434_ VGND VGND VPWR VPWR cpuregs\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12294_ decoded_imm\[26\] net733 VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__and2_1
XFILLER_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14033_ clknet_leaf_179_clk _00487_ VGND VGND VPWR VPWR cpuregs\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11245_ cpuregs\[8\]\[24\] net686 VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06799__A net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11176_ net831 _05849_ _05851_ _05853_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__a211o_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10127_ _04848_ _04849_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__nor2_1
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10058_ _04804_ _04805_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__nor2_1
X_14935_ clknet_leaf_6_clk _01287_ VGND VGND VPWR VPWR cpuregs\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07515__A1 net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11644__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07515__B2 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14866_ clknet_leaf_20_clk _01218_ VGND VGND VPWR VPWR cpuregs\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10768__B _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09114__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13817_ clknet_leaf_191_clk _00271_ VGND VGND VPWR VPWR cpuregs\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14797_ clknet_leaf_75_clk _01149_ VGND VGND VPWR VPWR decoded_imm\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_21_clk _00202_ VGND VGND VPWR VPWR cpuregs\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10822__A1 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ clknet_leaf_146_clk _00133_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_15418_ clknet_leaf_43_clk _01757_ VGND VGND VPWR VPWR cpuregs\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09976__C1 net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15349_ clknet_leaf_42_clk _01689_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_1
XANTENNA__10586__B1 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold104 cpuregs\[26\]\[31\] VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold115 cpuregs\[14\]\[13\] VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 cpuregs\[22\]\[19\] VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 cpuregs\[28\]\[2\] VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 net163 VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 cpuregs\[14\]\[27\] VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _04686_ _04688_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout606 _03148_ VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07203__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout617 net620 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__buf_2
X_09841_ _04621_ _04622_ _04625_ net1182 VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__o211a_1
Xfanout628 net631 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload14_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout639 net645 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_2
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07317__B _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09772_ _04433_ _04551_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__nand2b_1
X_06984_ genblk2.pcpi_div.dividend\[9\] _02553_ net1119 VGND VGND VPWR VPWR _02560_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_67_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08723_ genblk1.genblk1.pcpi_mul.rd\[37\] genblk1.genblk1.pcpi_mul.next_rs2\[38\]
+ net1099 VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__nand3_1
XFILLER_27_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__inv_2
XFILLER_26_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10510__B1 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09024__S net519 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07605_ _03125_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout444_A net446 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_A net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07536_ net19 net938 net937 VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12263__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12385__S net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11471__D1 net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07987__B net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07467_ net14 net938 net936 VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout611_A net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout709_A _02501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09206_ net1766 net409 net492 VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__mux2_1
XFILLER_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07398_ count_cycle\[16\] net974 net844 _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__o211a_1
XANTENNA__13212__C1 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11369__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09137_ net1616 net539 net500 VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__mux2_1
XANTENNA__10041__A2 _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09068_ net1507 net524 net508 VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__mux2_1
XFILLER_162_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout980_A net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08019_ net968 _03358_ _03360_ net930 _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__o221a_1
XANTENNA__12318__B2 mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11956__C _02443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold660 cpuregs\[8\]\[0\] VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 cpuregs\[10\]\[26\] VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold682 cpuregs\[6\]\[13\] VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net1075 _05710_ net855 VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold693 cpuregs\[29\]\[2\] VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout866_X net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07227__B decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12981_ net1480 net347 net447 VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__mux2_1
Xhold1360 genblk1.genblk1.pcpi_mul.rdx\[4\] VGND VGND VPWR VPWR net2674 sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ clknet_leaf_155_clk _01105_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[31\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1371 genblk2.pcpi_div.quotient\[6\] VGND VGND VPWR VPWR net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1382 genblk1.genblk1.pcpi_mul.rd\[30\] VGND VGND VPWR VPWR net2696 sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ _06258_ _06402_ net384 VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__a21oi_2
XFILLER_91_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1393 genblk1.genblk1.pcpi_mul.rd\[58\] VGND VGND VPWR VPWR net2707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10501__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08170__A1 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14651_ clknet_leaf_157_clk _01036_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11863_ _06332_ _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__and2_1
XFILLER_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10814_ cpuregs\[12\]\[13\] cpuregs\[13\]\[13\] net651 VGND VGND VPWR VPWR _05501_
+ sky130_fd_sc_hd__mux2_1
X_13602_ clknet_leaf_192_clk _00057_ VGND VGND VPWR VPWR cpuregs\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11057__A1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12254__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14582_ clknet_leaf_69_clk _00968_ VGND VGND VPWR VPWR latched_rd\[3\] sky130_fd_sc_hd__dfxtp_2
X_11794_ genblk2.pcpi_div.dividend\[28\] genblk2.pcpi_div.divisor\[28\] VGND VGND
+ VPWR VPWR _06265_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_31_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ net350 net1816 net415 VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__mux2_1
X_10745_ _05432_ _05433_ net813 VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__mux2_1
XFILLER_41_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12006__B1 net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13464_ net1544 net407 net424 VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__mux2_1
X_10676_ cpuregs\[11\]\[9\] net628 net593 _05366_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_62_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__C1 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12415_ net309 net1986 net472 VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__mux2_1
X_15203_ clknet_leaf_36_clk _01552_ VGND VGND VPWR VPWR cpuregs\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08225__A2 net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13395_ net2764 net397 _02297_ _02303_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__o22a_1
XFILLER_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15134_ clknet_leaf_12_clk _01486_ VGND VGND VPWR VPWR cpuregs\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12346_ mem_rdata_q\[22\] _06223_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__and2_1
Xoutput209 net1021 VGND VGND VPWR VPWR pcpi_rs1[15] sky130_fd_sc_hd__buf_2
XFILLER_142_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15065_ clknet_leaf_104_clk net2234 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12277_ _06616_ net2960 _06613_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__mux2_1
X_14016_ clknet_leaf_1_clk _00470_ VGND VGND VPWR VPWR cpuregs\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09109__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output73_A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11228_ cpuregs\[16\]\[24\] net699 VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__or2_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11159_ net792 _05832_ _05834_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__or4_1
XANTENNA__08948__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14918_ clknet_leaf_111_clk _01270_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08161__A1 _02396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14849_ clknet_leaf_57_clk _01201_ VGND VGND VPWR VPWR cpuregs\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12245__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08370_ reg_pc\[10\] _03780_ reg_pc\[11\] VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__a21oi_1
XFILLER_90_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07321_ _02835_ _02848_ _02861_ _02846_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__o31ai_1
XFILLER_149_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07252_ net1048 net7 _02797_ net1052 net1057 VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__o2111a_1
XFILLER_31_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07183_ reg_pc\[3\] decoded_imm\[3\] VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__or2_1
XANTENNA__08216__A2 net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08271__X net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07903__A_N net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10453__S net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12234__A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09527__B net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09019__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout403 net404 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09716__A2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout414 _02358_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout425 net426 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__buf_4
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07727__A1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout394_A _04888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout436 net438 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_4
XFILLER_87_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout447 net448 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__buf_4
XANTENNA__12720__B2 net1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09824_ _02481_ _04608_ _04609_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__or3_1
Xfanout458 _02119_ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__buf_2
Xfanout469 net470 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_4
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06967_ net1120 _02544_ genblk2.pcpi_div.quotient\[7\] VGND VGND VPWR VPWR _02546_
+ sky130_fd_sc_hd__a21oi_1
X_09755_ _04524_ _04534_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout659_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11287__A1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08706_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__inv_2
X_09686_ decoded_imm_j\[5\] _04426_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__and2_1
X_06898_ net1232 _02445_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__and2_1
XFILLER_82_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08637_ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_159_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_X net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A _03137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1189_X net1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11039__A1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07998__A net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08568_ _03946_ _03948_ _03941_ _03944_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a211o_1
XANTENNA__13433__C1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08446__X _03849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10695__Y _05386_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07519_ reg_pc\[25\] decoded_imm\[25\] VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__nand2_1
XFILLER_167_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08499_ net894 _03888_ _03890_ net2624 net1199 VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout614_X net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13004__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ cpuregs\[28\]\[5\] cpuregs\[29\]\[5\] net678 VGND VGND VPWR VPWR _05225_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12539__A1 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10461_ _05159_ _05160_ net804 VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__mux2_1
XANTENNA__09404__A1 net1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12843__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13200__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12200_ net748 net2835 VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13180_ net1857 net345 net428 VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10392_ net1223 _05096_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__nand2_1
XFILLER_108_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout983_X net983 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10871__B net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12131_ _06568_ _06569_ _06570_ _06571_ net274 VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__o221a_1
XANTENNA__10363__S net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10970__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12062_ net863 _06363_ _06512_ _06511_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__a31o_1
Xhold490 cpuregs\[23\]\[10\] VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ cpuregs\[28\]\[18\] cpuregs\[29\]\[18\] net648 VGND VGND VPWR VPWR _05695_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout970 _02428_ VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout981 net983 VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__buf_4
Xfanout992 net993 VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__clkbuf_4
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11278__B2 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12964_ net286 net2453 net453 VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__mux2_1
XFILLER_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1190 genblk1.genblk1.pcpi_mul.next_rs1\[43\] VGND VGND VPWR VPWR net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_14703_ clknet_leaf_153_clk _01088_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_11915_ _06263_ _06384_ _06262_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__a21o_1
XFILLER_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output111_A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _04283_ _06663_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__or2_2
XANTENNA_output209_A net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14634_ clknet_leaf_170_clk _01019_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11846_ genblk2.pcpi_div.divisor\[2\] genblk2.pcpi_div.dividend\[2\] VGND VGND VPWR
+ VPWR _06317_ sky130_fd_sc_hd__nand2b_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11_0_clk_X clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13422__B net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11777_ _02418_ _02448_ net964 _06239_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__or4_1
X_14565_ clknet_leaf_43_clk _00951_ VGND VGND VPWR VPWR cpuregs\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09643__B2 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13516_ net1787 net290 net421 VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__mux2_1
X_10728_ cpuregs\[19\]\[10\] net626 net593 VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_60_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14496_ clknet_leaf_95_clk _00885_ VGND VGND VPWR VPWR instr_xor sky130_fd_sc_hd__dfxtp_1
XFILLER_146_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13447_ net961 _05034_ _02348_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__nor3_1
X_10659_ net773 _05342_ _05350_ _05334_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__a31oi_4
Xclkload13 clknet_4_14_0_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_8
Xclkload24 clknet_leaf_198_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__clkinv_2
Xclkload35 clknet_leaf_188_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__inv_8
XANTENNA__11202__A1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload46/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13378_ _04910_ _05011_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__nand2_1
Xclkload57 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__inv_8
Xclkload68 clknet_leaf_172_clk VGND VGND VPWR VPWR clkload68/Y sky130_fd_sc_hd__inv_6
XANTENNA__07957__A1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload79 clknet_leaf_162_clk VGND VGND VPWR VPWR clkload79/Y sky130_fd_sc_hd__bufinv_16
X_15117_ clknet_leaf_21_clk _01469_ VGND VGND VPWR VPWR cpuregs\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12329_ decoded_imm\[10\] net735 _06643_ mem_rdata_q\[30\] _06644_ VGND VGND VPWR
+ VPWR _01164_ sky130_fd_sc_hd__a221o_1
XFILLER_170_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10961__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07148__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15048_ clknet_leaf_108_clk _01400_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13584__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07870_ _03335_ _03348_ _03356_ _03365_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__or4_1
X_06821_ instr_fence instr_and instr_sra instr_xor VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09540_ count_instr\[46\] _04387_ _04389_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__o21a_1
X_06752_ genblk2.pcpi_div.divisor\[16\] VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__inv_2
XFILLER_36_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10477__C1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09471_ _04344_ _04345_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__nor2_1
X_08422_ reg_pc\[21\] reg_pc\[20\] _03821_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__and3_1
XFILLER_51_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09302__S net482 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08353_ _03770_ _03773_ net766 VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__mux2_4
XFILLER_149_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07304_ reg_pc\[11\] decoded_imm\[11\] VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_154_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08284_ reg_out\[19\] reg_next_pc\[19\] net922 VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__mux2_1
XANTENNA__07645__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload7 clknet_4_7_0_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_8
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07235_ _02383_ net24 _02781_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__o21a_1
XFILLER_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1149_A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07166_ net1048 net2 net1057 net1052 VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_132_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07948__A1 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07097_ genblk2.pcpi_div.dividend\[25\] genblk2.pcpi_div.dividend\[24\] _02647_ VGND
+ VGND VPWR VPWR _02657_ sky130_fd_sc_hd__or3_1
XANTENNA__10036__X _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1209 _02378_ VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_X net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13494__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout776_A net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07345__X _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout277 _06403_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_2
X_09807_ _04566_ _04581_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__nand2_1
Xfanout288 _03865_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout299 _03852_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_2
X_07999_ net1143 _03428_ _03429_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout943_A _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_X net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12457__B1 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09738_ net984 _04529_ _04530_ _02380_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__a31o_1
XFILLER_43_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12838__S net460 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09669_ _04465_ _04466_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout829_X net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11742__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11700_ net1991 net337 net374 VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__mux2_1
X_12680_ net1193 genblk1.genblk1.pcpi_mul.next_rs2\[45\] net886 net2826 net711 VGND
+ VGND VPWR VPWR _01350_ sky130_fd_sc_hd__a221o_1
XANTENNA__10483__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09212__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11631_ net3029 net737 _06206_ _06217_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__a22o_1
XFILLER_70_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09625__B2 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ net2609 net561 _06178_ _06182_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14350_ clknet_leaf_67_clk _06739_ VGND VGND VPWR VPWR reg_out\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11432__A1 net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14127__Q net267 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13301_ _02215_ _02216_ _02220_ net395 net1027 VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__o32a_1
X_10513_ net1175 net860 _05208_ _03264_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__o22a_1
XFILLER_155_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14281_ clknet_leaf_100_clk _00735_ VGND VGND VPWR VPWR count_cycle\[26\] sky130_fd_sc_hd__dfxtp_1
X_11493_ net3036 _02455_ _06156_ latched_is_lb VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__a22o_1
XANTENNA__12573__S net470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13232_ net1044 net1040 net755 VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__mux2_1
X_10444_ cpuregs\[14\]\[0\] cpuregs\[15\]\[0\] net685 VGND VGND VPWR VPWR _05144_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12932__A1 net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13163_ net1458 _03870_ net434 VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__mux2_1
X_10375_ net1068 net760 _05078_ net566 reg_pc\[31\] VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__a32o_1
XFILLER_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12114_ genblk2.pcpi_div.dividend\[27\] _06557_ net275 VGND VGND VPWR VPWR _01036_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13094_ net290 net2130 net441 VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__mux2_1
XFILLER_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12045_ _06285_ _06359_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__nand2b_1
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07167__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12160__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06914__A2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07415__B _02945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13996_ clknet_leaf_53_clk _00450_ VGND VGND VPWR VPWR cpuregs\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12947_ net353 net2231 net452 VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__mux2_1
XANTENNA__11120__B1 net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11652__S net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08086__X alu_out\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12878_ mem_rdata_q\[15\] net7 net962 VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__mux2_1
XANTENNA__09122__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10776__B net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14617_ clknet_leaf_93_clk _01003_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dfxtp_1
X_11829_ genblk2.pcpi_div.divisor\[11\] genblk2.pcpi_div.dividend\[11\] VGND VGND
+ VPWR VPWR _06300_ sky130_fd_sc_hd__and2b_1
XFILLER_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15597_ clknet_leaf_192_clk _01933_ VGND VGND VPWR VPWR cpuregs\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12049__A net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14548_ clknet_leaf_24_clk _00934_ VGND VGND VPWR VPWR cpuregs\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08961__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13579__S net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10631__C1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14479_ clknet_leaf_96_clk _00868_ VGND VGND VPWR VPWR instr_lhu sky130_fd_sc_hd__dfxtp_1
Xclkload102 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload102/Y sky130_fd_sc_hd__inv_8
Xclkload113 clknet_leaf_48_clk VGND VGND VPWR VPWR clkload113/Y sky130_fd_sc_hd__clkinv_4
X_07020_ genblk2.pcpi_div.dividend\[14\] _02584_ net1115 VGND VGND VPWR VPWR _02591_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__13176__A1 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload124 clknet_leaf_53_clk VGND VGND VPWR VPWR clkload124/Y sky130_fd_sc_hd__bufinv_16
Xclkload135 clknet_leaf_68_clk VGND VGND VPWR VPWR clkload135/Y sky130_fd_sc_hd__inv_6
XFILLER_162_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload146 clknet_leaf_129_clk VGND VGND VPWR VPWR clkload146/Y sky130_fd_sc_hd__clkinv_2
XFILLER_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11187__B1 net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload157 clknet_leaf_117_clk VGND VGND VPWR VPWR clkload157/Y sky130_fd_sc_hd__inv_6
Xclkload168 clknet_leaf_86_clk VGND VGND VPWR VPWR clkload168/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload179 clknet_leaf_99_clk VGND VGND VPWR VPWR clkload179/Y sky130_fd_sc_hd__clkinv_8
XFILLER_170_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08971_ net1460 _04262_ net945 VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__mux2_1
XFILLER_115_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07922_ net252 net1002 VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__and2b_1
Xhold19 net62 VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07853_ net258 net992 VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__nor2_1
XFILLER_69_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08201__S net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06804_ net996 VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__inv_2
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07784_ _03298_ _03300_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09523_ count_instr\[40\] _04377_ net1214 VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10967__A net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09454_ count_instr\[16\] _04332_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1099_A net1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10465__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11662__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09032__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08405_ net332 net2131 net528 VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__mux2_1
X_09385_ net1837 net316 net399 VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout524_A _03774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08336_ _03758_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__nor2_1
XANTENNA__08291__A0 net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13489__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08267_ net1029 _03717_ net981 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__mux2_1
XANTENNA__07995__B net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12393__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_140_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1054_X net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07218_ net1052 net1057 _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__and3_1
X_08198_ _03370_ net931 net969 VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout893_A net898 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07149_ net991 _02387_ _02701_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__and3_2
XANTENNA__07397__A2 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10160_ count_cycle\[58\] count_cycle\[59\] _04868_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout779_X net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1006 net218 VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11737__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1017 net211 VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__dlymetal6s2s_1
X_10091_ net2940 _04825_ net1228 VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__o21ai_1
XFILLER_126_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1028 net205 VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__buf_2
Xfanout1039 net231 VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09207__S net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12142__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15506__Q net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15733__A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13850_ clknet_leaf_198_clk _00304_ VGND VGND VPWR VPWR cpuregs\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_145_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12801_ net575 net2311 net464 VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__mux2_1
XANTENNA__09731__A decoded_imm_j\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_172_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13781_ clknet_leaf_20_clk _00235_ VGND VGND VPWR VPWR cpuregs\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_10993_ net1078 _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__nand2_1
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11102__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15520_ clknet_leaf_81_clk _01856_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11653__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12732_ _02407_ net911 VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__nor2_1
XANTENNA__10456__A2 net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07251__A _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15451_ clknet_leaf_17_clk _01790_ VGND VGND VPWR VPWR cpuregs\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12663_ net1218 genblk1.genblk1.pcpi_mul.next_rs2\[31\] net917 net258 VGND VGND VPWR
+ VPWR _02081_ sky130_fd_sc_hd__a22o_1
X_14402_ clknet_leaf_130_clk alu_out\[2\] VGND VGND VPWR VPWR alu_out_q\[2\] sky130_fd_sc_hd__dfxtp_1
X_11614_ net1862 net741 _06203_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_187_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15382_ clknet_leaf_8_clk _01721_ VGND VGND VPWR VPWR cpuregs\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12594_ net317 net2356 net470 VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__mux2_1
XFILLER_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14333_ clknet_leaf_177_clk _06720_ VGND VGND VPWR VPWR reg_out\[13\] sky130_fd_sc_hd__dfxtp_1
X_11545_ _06166_ _06169_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__nor2_1
XFILLER_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_131_clk sky130_fd_sc_hd__clkbuf_8
X_11476_ net258 net857 _06144_ _06145_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__a22o_1
X_14264_ clknet_leaf_122_clk _00718_ VGND VGND VPWR VPWR count_cycle\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10427_ _02489_ _05125_ _05129_ _05121_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__o211a_1
X_13215_ _04949_ _04955_ _04954_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__a21o_1
XANTENNA__11220__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14195_ clknet_leaf_132_clk _00649_ VGND VGND VPWR VPWR reg_pc\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10358_ cpuregs\[19\]\[31\] net638 net599 VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__o21a_1
X_13146_ net1499 net348 net431 VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__mux2_1
XFILLER_151_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11647__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13077_ net356 net1893 net439 VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _04987_ _04989_ _04990_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12028_ genblk2.pcpi_div.dividend\[15\] _06483_ net269 VGND VGND VPWR VPWR _01024_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09117__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_198_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_198_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11593__D mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08956__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13979_ clknet_leaf_196_clk _00433_ VGND VGND VPWR VPWR cpuregs\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10447__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11644__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15649_ clknet_leaf_49_clk _01985_ VGND VGND VPWR VPWR cpuregs\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09170_ net537 net2208 net496 VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__mux2_1
XFILLER_159_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08121_ net966 _03331_ _03333_ net929 _03617_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__a221o_1
XANTENNA__08273__A0 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07076__B2 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_122_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_147_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13102__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08052_ _03377_ net932 _03378_ net968 VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07003_ net1118 genblk2.pcpi_div.quotient\[12\] _02575_ net950 VGND VGND VPWR VPWR
+ _02577_ sky130_fd_sc_hd__a31o_1
XANTENNA__08025__B1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12941__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10368__D1 net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07379__A2 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13338__A net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10461__S net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08954_ genblk1.genblk1.pcpi_mul.rd\[15\] genblk1.genblk1.pcpi_mul.rd\[47\] net954
+ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__mux2_1
XANTENNA__09535__B net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_A net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09027__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1701 mem_rdata_q\[5\] VGND VGND VPWR VPWR net3015 sky130_fd_sc_hd__dlygate4sd3_1
X_07905_ _03285_ _03422_ _03421_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__o21ai_1
Xhold1712 latched_is_lh VGND VGND VPWR VPWR net3026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08885_ _04215_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_189_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_189_clk sky130_fd_sc_hd__clkbuf_8
Xhold1723 reg_pc\[19\] VGND VGND VPWR VPWR net3037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 mem_rdata_q\[2\] VGND VGND VPWR VPWR net3048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout474_A _06664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1745 reg_pc\[23\] VGND VGND VPWR VPWR net3059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1756 genblk1.genblk1.pcpi_mul.next_rs2\[46\] VGND VGND VPWR VPWR net3070 sky130_fd_sc_hd__dlygate4sd3_1
X_07836_ _03352_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__and2_1
XFILLER_38_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12388__S net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09828__A1 net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07767_ net1047 net1178 VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout641_A net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09828__B2 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09506_ count_instr\[34\] count_instr\[33\] count_instr\[32\] VGND VGND VPWR VPWR
+ _04368_ sky130_fd_sc_hd__and3_1
XFILLER_72_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07698_ cpuregs\[20\]\[3\] cpuregs\[21\]\[3\] net674 VGND VGND VPWR VPWR _03218_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09437_ count_instr\[10\] count_instr\[9\] _04318_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1171_X net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ net1941 net573 net402 VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__mux2_1
X_08319_ latched_branch _02368_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_113_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_8
X_09299_ net1746 net584 net481 VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__mux2_1
XANTENNA__13012__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ cpuregs\[4\]\[27\] cpuregs\[5\]\[27\] net695 VGND VGND VPWR VPWR _06003_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_169_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11261_ net836 _05931_ _05935_ net786 VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__a211o_1
XANTENNA__15728__A net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12851__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13000_ _06255_ _06611_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__and2_1
XFILLER_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10212_ _04916_ _04917_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__nor2_1
XFILLER_122_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09726__A net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11192_ cpuregs\[16\]\[23\] net685 VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__or2_1
XFILLER_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10143_ count_cycle\[51\] count_cycle\[52\] count_cycle\[53\] _04854_ VGND VGND VPWR
+ VPWR _04860_ sky130_fd_sc_hd__and4_2
XPHY_EDGE_ROW_120_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10074_ count_cycle\[26\] count_cycle\[27\] count_cycle\[28\] _04811_ VGND VGND VPWR
+ VPWR _04816_ sky130_fd_sc_hd__and4_1
X_14951_ clknet_leaf_47_clk _01303_ VGND VGND VPWR VPWR cpuregs\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13902_ clknet_leaf_37_clk _00356_ VGND VGND VPWR VPWR cpuregs\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14882_ clknet_leaf_34_clk _01234_ VGND VGND VPWR VPWR cpuregs\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13833_ clknet_leaf_48_clk _00287_ VGND VGND VPWR VPWR cpuregs\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10429__A2 _03457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10400__A net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13764_ clknet_leaf_40_clk _00218_ VGND VGND VPWR VPWR cpuregs\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10976_ cpuregs\[20\]\[17\] cpuregs\[21\]\[17\] net646 VGND VGND VPWR VPWR _05659_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15503_ clknet_leaf_171_clk _01839_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dfxtp_1
X_12715_ net1354 net883 _02091_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__a21o_1
X_13695_ clknet_leaf_147_clk _00149_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15434_ clknet_leaf_181_clk _01773_ VGND VGND VPWR VPWR cpuregs\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12646_ net2823 net895 _02072_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_96_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08255__A0 net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_104_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_8
X_15365_ clknet_leaf_45_clk _01704_ VGND VGND VPWR VPWR cpuregs\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12577_ net571 net2268 net468 VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__mux2_1
XFILLER_157_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14316_ clknet_leaf_93_clk _00770_ VGND VGND VPWR VPWR count_cycle\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11528_ mem_rdata_q\[21\] net1896 net742 VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__mux2_1
XFILLER_129_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10601__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15296_ clknet_leaf_54_clk _01637_ VGND VGND VPWR VPWR cpuregs\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold308 cpuregs\[30\]\[10\] VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold319 genblk1.genblk1.pcpi_mul.pcpi_rd\[3\] VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14247_ clknet_leaf_75_clk _00701_ VGND VGND VPWR VPWR reg_next_pc\[24\] sky130_fd_sc_hd__dfxtp_1
X_11459_ cpuregs\[16\]\[30\] net688 VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__or2_1
XANTENNA__11011__C1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14178_ clknet_leaf_109_clk net2585 VGND VGND VPWR VPWR count_instr\[49\] sky130_fd_sc_hd__dfxtp_1
X_13129_ net282 net2486 net438 VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__mux2_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1008 cpuregs\[23\]\[1\] VGND VGND VPWR VPWR net2322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_140_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1019 cpuregs\[9\]\[3\] VGND VGND VPWR VPWR net2333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08670_ genblk1.genblk1.pcpi_mul.rd\[29\] genblk1.genblk1.pcpi_mul.next_rs2\[30\]
+ net1106 VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__and3_1
XFILLER_94_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14985__Q genblk1.genblk1.pcpi_mul.next_rs2\[32\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07621_ net986 decoded_imm_j\[1\] _03141_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ count_instr\[27\] net1138 net978 _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07483_ count_instr\[22\] net1137 net978 _03013_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__a211o_1
XFILLER_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11093__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12936__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09222_ net1820 net303 net495 VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__mux2_1
XFILLER_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09310__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09153_ net2020 net314 net502 VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__mux2_1
XANTENNA__13340__B net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11779__C net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08104_ net1144 _03600_ _03601_ _03602_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__a22o_1
X_09084_ net1538 net311 net510 VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__mux2_1
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08035_ net968 _03299_ net934 _03298_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__o22a_1
XFILLER_162_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold820 cpuregs\[9\]\[10\] VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 cpuregs\[25\]\[29\] VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 cpuregs\[18\]\[10\] VGND VGND VPWR VPWR net2156 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__B1 _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07618__X _03139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12345__A2 net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold853 cpuregs\[1\]\[25\] VGND VGND VPWR VPWR net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold864 cpuregs\[3\]\[17\] VGND VGND VPWR VPWR net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 cpuregs\[6\]\[16\] VGND VGND VPWR VPWR net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06889__B is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold886 cpuregs\[6\]\[14\] VGND VGND VPWR VPWR net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 cpuregs\[5\]\[5\] VGND VGND VPWR VPWR net2211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09986_ _04450_ _04451_ _04736_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__and3_1
XFILLER_131_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08937_ net2837 _04245_ net944 VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout477_X net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A net859 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1520 genblk2.pcpi_div.quotient\[13\] VGND VGND VPWR VPWR net2834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1531 genblk1.genblk1.pcpi_mul.next_rs2\[51\] VGND VGND VPWR VPWR net2845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 genblk2.pcpi_div.quotient_msk\[17\] VGND VGND VPWR VPWR net2856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08868_ _04201_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__xnor2_1
Xhold1553 genblk2.pcpi_div.quotient_msk\[24\] VGND VGND VPWR VPWR net2867 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12700__A _02384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1564 genblk1.genblk1.pcpi_mul.rd\[57\] VGND VGND VPWR VPWR net2878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1575 count_instr\[56\] VGND VGND VPWR VPWR net2889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07819_ net244 net1014 VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__and2_1
Xhold1586 genblk1.genblk1.pcpi_mul.next_rs2\[57\] VGND VGND VPWR VPWR net2900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 genblk1.genblk1.pcpi_mul.rd\[11\] VGND VGND VPWR VPWR net2911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout644_X net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08799_ genblk1.genblk1.pcpi_mul.next_rs2\[50\] net1096 genblk1.genblk1.pcpi_mul.rd\[49\]
+ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__a21o_1
XFILLER_72_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13007__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10830_ net823 _05512_ _05514_ _05516_ net787 VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10220__A decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12846__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10761_ cpuregs\[8\]\[11\] net666 VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout811_X net811 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12500_ net871 _01993_ _01994_ net387 VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__a31o_1
X_13480_ net1560 net303 net425 VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__mux2_1
X_10692_ cpuregs\[19\]\[9\] net627 net594 VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__o21a_1
XFILLER_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09220__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08237__A0 net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12431_ genblk1.genblk1.pcpi_mul.mul_counter\[3\] genblk1.genblk1.pcpi_mul.mul_counter\[2\]
+ _06666_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__or3_1
XFILLER_139_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15150_ clknet_leaf_91_clk _01499_ VGND VGND VPWR VPWR mem_rdata_q\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12362_ net1377 net573 net361 VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__mux2_1
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10595__A1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14101_ clknet_leaf_186_clk _00555_ VGND VGND VPWR VPWR cpuregs\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11313_ cpuregs\[25\]\[26\] net643 net615 _05986_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_91_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15081_ clknet_leaf_105_clk _01433_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12293_ mem_rdata_q\[27\] net559 _06625_ net532 VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__a211o_1
XANTENNA__10890__A net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12581__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14032_ clknet_leaf_32_clk _00486_ VGND VGND VPWR VPWR cpuregs\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11244_ net818 _05917_ _05919_ net834 VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__o211a_1
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11175_ cpuregs\[18\]\[22\] net554 _05852_ net783 VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__o22a_1
X_10126_ count_cycle\[47\] _04846_ net1228 VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__o21ai_1
XANTENNA_output239_A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10057_ net2851 _04802_ net1235 VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__o21ai_1
X_14934_ clknet_leaf_20_clk _01286_ VGND VGND VPWR VPWR cpuregs\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07515__A2 net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14865_ clknet_leaf_181_clk _01217_ VGND VGND VPWR VPWR cpuregs\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload0_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13816_ clknet_leaf_187_clk _00270_ VGND VGND VPWR VPWR cpuregs\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_14796_ clknet_leaf_67_clk _01148_ VGND VGND VPWR VPWR decoded_imm\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12272__A1 net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13747_ clknet_leaf_21_clk _00201_ VGND VGND VPWR VPWR cpuregs\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10959_ _05640_ _05641_ net811 VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__mux2_1
XANTENNA__11660__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13441__A net570 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13678_ clknet_leaf_146_clk _00132_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15417_ clknet_leaf_16_clk _01756_ VGND VGND VPWR VPWR cpuregs\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12629_ net1192 genblk1.genblk1.pcpi_mul.next_rs2\[14\] net915 net1163 VGND VGND
+ VPWR VPWR _02064_ sky130_fd_sc_hd__a22o_1
XANTENNA__08228__B1 net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12057__A net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13221__B1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15348_ clknet_leaf_13_clk _01688_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_1
Xhold105 net35 VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 cpuregs\[29\]\[10\] VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ clknet_leaf_196_clk _01620_ VGND VGND VPWR VPWR cpuregs\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold127 cpuregs\[26\]\[14\] VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07585__S net1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold138 cpuregs\[26\]\[16\] VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_137_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold149 cpuregs\[12\]\[7\] VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11535__A0 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout607 net609 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkbuf_4
X_09840_ net984 _04623_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__nand3_1
XFILLER_99_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14422__D alu_out\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout618 net620 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__buf_2
Xfanout629 net631 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_2
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09771_ _04551_ _04433_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__nand2b_1
X_06983_ net948 _02554_ _02555_ _02559_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__o31ai_1
XFILLER_101_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08722_ genblk1.genblk1.pcpi_mul.rd\[37\] genblk1.genblk1.pcpi_mul.next_rs2\[38\]
+ net1099 VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__and3_1
XANTENNA__08269__X net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09305__S net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07614__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08653_ _04013_ _04016_ _04018_ _04019_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__o211a_1
XFILLER_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07604_ reg_pc\[31\] decoded_imm\[31\] VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__xnor2_1
X_08584_ genblk1.genblk1.pcpi_mul.rd\[16\] genblk1.genblk1.pcpi_mul.rdx\[16\] VGND
+ VGND VPWR VPWR _03962_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_120_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07535_ _03047_ _03049_ _03060_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__nand3_1
XFILLER_169_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1081_A net1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_A net438 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07466_ _02994_ _02996_ _02997_ net1073 VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__o211a_1
XFILLER_168_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09040__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09205_ net1851 net522 net492 VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__mux2_1
XANTENNA__12015__A1 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08219__B1 net266 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07397_ count_instr\[16\] net1136 net977 _02933_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout604_A net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09967__B1 net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09136_ net1750 net542 net501 VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__mux2_1
XFILLER_108_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13497__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09067_ net2129 net539 net508 VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__mux2_1
XFILLER_118_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1134_X net1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07348__X _02888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08018_ _03357_ net934 VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__or2_1
XFILLER_104_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11526__A0 mem_rdata_q\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold650 cpuregs\[8\]\[6\] VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 cpuregs\[15\]\[12\] VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold672 cpuregs\[4\]\[23\] VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14332__D _06719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold683 cpuregs\[29\]\[24\] VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 cpuregs\[10\]\[3\] VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10215__A decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09969_ net1129 _04450_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout859_X net859 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11745__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12980_ net1344 net350 net447 VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__mux2_1
XFILLER_94_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1350 genblk2.pcpi_div.divisor\[49\] VGND VGND VPWR VPWR net2664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09215__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1361 reg_next_pc\[12\] VGND VGND VPWR VPWR net2675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11931_ _06259_ _06388_ _06400_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__o21ai_1
Xhold1372 _06585_ VGND VGND VPWR VPWR net2686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1383 genblk1.genblk1.pcpi_mul.rd\[46\] VGND VGND VPWR VPWR net2697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 genblk1.genblk1.pcpi_mul.rdx\[52\] VGND VGND VPWR VPWR net2708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08170__A2 net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14650_ clknet_leaf_157_clk _01035_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11862_ genblk2.pcpi_div.divisor\[8\] genblk2.pcpi_div.dividend\[8\] VGND VGND VPWR
+ VPWR _06333_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13601_ clknet_leaf_178_clk _00056_ VGND VGND VPWR VPWR cpuregs\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10813_ _05497_ _05499_ net779 VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__a21o_1
X_14581_ clknet_leaf_69_clk _00967_ VGND VGND VPWR VPWR latched_rd\[2\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__12576__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13451__B1 _06143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11793_ genblk2.pcpi_div.divisor\[28\] genblk2.pcpi_div.dividend\[28\] VGND VGND
+ VPWR VPWR _06264_ sky130_fd_sc_hd__and2b_1
XFILLER_41_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13532_ net354 net1983 net416 VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__mux2_1
XFILLER_159_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10744_ cpuregs\[20\]\[11\] cpuregs\[21\]\[11\] net665 VGND VGND VPWR VPWR _05433_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12006__A1 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13463_ net1634 net520 net424 VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__mux2_1
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10675_ cpuregs\[10\]\[9\] net667 VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1290 VGND VGND VPWR VPWR picorv32_1290/HI trace_data[12] sky130_fd_sc_hd__conb_1
X_15202_ clknet_leaf_38_clk _01551_ VGND VGND VPWR VPWR cpuregs\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12414_ net314 net2166 net473 VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__mux2_1
X_13394_ net393 _02298_ _02300_ _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__or4_1
XFILLER_127_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15133_ clknet_leaf_41_clk _01485_ VGND VGND VPWR VPWR cpuregs\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12345_ decoded_imm\[3\] net745 _06652_ _06653_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__o22a_1
XFILLER_154_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15064_ clknet_leaf_104_clk net2518 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11517__A0 mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12276_ _06239_ _06614_ net730 VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__o21bai_1
XFILLER_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14015_ clknet_leaf_0_clk _00469_ VGND VGND VPWR VPWR cpuregs\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11227_ _05901_ _05902_ net818 VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__mux2_1
XFILLER_96_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output66_A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11158_ cpuregs\[11\]\[22\] net633 net597 _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__o211a_1
XFILLER_96_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11655__S net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10109_ count_cycle\[41\] _04836_ net1204 VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__a21oi_1
X_11089_ cpuregs\[4\]\[20\] net661 VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__or2_1
XANTENNA__12340__A mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09125__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14917_ clknet_leaf_111_clk _01269_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08161__A2 net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14848_ clknet_leaf_60_clk _01200_ VGND VGND VPWR VPWR cpuregs\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08964__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10795__A net797 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14779_ clknet_leaf_154_clk _00034_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07320_ _02807_ _02822_ _02821_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__o21a_1
XFILLER_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07251_ _02383_ net25 VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__or2_1
XANTENNA__14417__D alu_out\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07672__A1 decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09949__B1 net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07182_ reg_pc\[3\] decoded_imm\[3\] VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nand2_1
XANTENNA__10019__B net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13110__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14503__Q instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout404 _03785_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout415 _02357_ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_8
Xfanout426 _02355_ VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__buf_4
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout437 net438 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_8
X_09823_ _04606_ _04607_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__and2b_1
Xfanout448 net450 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_8
Xfanout459 _02118_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10731__A1 net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13346__A net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09754_ _04543_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__nor2_1
XANTENNA__07615__Y _03136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06966_ net1120 genblk2.pcpi_div.quotient\[7\] _02544_ VGND VGND VPWR VPWR _02545_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09035__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08705_ _04057_ _04060_ _04062_ _04063_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__o211a_1
XFILLER_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09685_ decoded_imm_j\[5\] _04426_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__nor2_1
X_06897_ _02491_ _02492_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout554_A _03156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08636_ genblk1.genblk1.pcpi_mul.rd\[24\] genblk1.genblk1.pcpi_mul.rdx\[24\] VGND
+ VGND VPWR VPWR _04006_ sky130_fd_sc_hd__nand2_1
XFILLER_54_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07360__B1 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07631__X _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08567_ genblk1.genblk1.pcpi_mul.rd\[13\] genblk1.genblk1.pcpi_mul.next_rs2\[14\]
+ net1093 VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__nand3_1
XANTENNA__12396__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09101__A1 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A net821 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07518_ reg_pc\[25\] decoded_imm\[25\] VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__nor2_1
XFILLER_23_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08498_ _03889_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__inv_2
XFILLER_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ _02930_ _02941_ _02953_ _02965_ _02981_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__o41a_1
XANTENNA_fanout607_X net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10460_ cpuregs\[30\]\[0\] cpuregs\[31\]\[0\] net684 VGND VGND VPWR VPWR _05160_
+ sky130_fd_sc_hd__mux2_1
XFILLER_148_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09119_ net1801 net302 net507 VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10391_ net864 _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__nand2_1
XANTENNA__13020__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12130_ net864 _06387_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__nand2_1
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07878__A_N net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12061_ _06278_ _06362_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__or2_1
Xhold480 cpuregs\[15\]\[20\] VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 cpuregs\[28\]\[8\] VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__B1 _02729_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11012_ cpuregs\[30\]\[18\] cpuregs\[31\]\[18\] net648 VGND VGND VPWR VPWR _05694_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10722__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13256__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout960 _02462_ VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout971 net972 VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__buf_2
Xfanout982 net983 VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 net226 VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__buf_4
XFILLER_18_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11278__A2 net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12475__A1 net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12963_ net291 net2495 net453 VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__mux2_1
XFILLER_45_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_84_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_8
Xhold1180 cpuregs\[17\]\[19\] VGND VGND VPWR VPWR net2494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _01413_ VGND VGND VPWR VPWR net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_14702_ clknet_leaf_153_clk _01087_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11914_ _06261_ _06263_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ mem_rdata_q\[31\] net25 net962 VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__mux2_1
XFILLER_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07351__B1 _02888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14633_ clknet_leaf_170_clk _01018_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ genblk2.pcpi_div.divisor\[2\] genblk2.pcpi_div.dividend\[2\] VGND VGND VPWR
+ VPWR _06316_ sky130_fd_sc_hd__and2b_1
XFILLER_14_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07701__B net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14564_ clknet_leaf_13_clk _00950_ VGND VGND VPWR VPWR cpuregs\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11776_ mem_do_wdata _02419_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__or2_1
XANTENNA__09643__A2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13515_ net2100 net295 net421 VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__mux2_1
XFILLER_14_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10727_ cpuregs\[17\]\[10\] net626 net607 _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__o211a_1
X_14495_ clknet_leaf_94_clk _00884_ VGND VGND VPWR VPWR instr_sltu sky130_fd_sc_hd__dfxtp_1
XFILLER_158_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13446_ _04894_ _05032_ _04893_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__o21a_1
XANTENNA__08052__A2_N net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10658_ net827 _05345_ _05347_ _05349_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__a211o_1
XFILLER_167_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload14 clknet_4_15_0_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__inv_8
Xclkload25 clknet_leaf_199_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__bufinv_16
Xclkload36 clknet_leaf_189_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__clkinv_8
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload47 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload47/X sky130_fd_sc_hd__clkbuf_8
X_13377_ _02282_ _02283_ _02287_ net397 net2556 VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__o32a_1
X_10589_ cpuregs\[4\]\[7\] cpuregs\[5\]\[7\] net659 VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__mux2_1
Xclkload58 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload58/Y sky130_fd_sc_hd__inv_6
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload69 clknet_leaf_149_clk VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__inv_8
X_15116_ clknet_leaf_28_clk _01468_ VGND VGND VPWR VPWR cpuregs\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12328_ net1148 decoded_imm_j\[10\] net743 VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__and3_1
XFILLER_141_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15047_ clknet_leaf_108_clk _01399_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_12259_ net2816 net381 net369 net2876 VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__a22o_1
XANTENNA__07148__B net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08959__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12163__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13360__C1 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06820_ instr_sll net1145 instr_add instr_andi VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__or4_1
XFILLER_68_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06751_ genblk2.pcpi_div.divisor\[20\] VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_75_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_8
X_09470_ net2825 _04342_ net1235 VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08421_ reg_pc\[20\] _03821_ reg_pc\[21\] VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13105__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08352_ _03771_ _03772_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_154_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ _02845_ _02843_ _02838_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_154_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12944__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08283_ net1014 _03725_ net981 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__mux2_2
Xclkload8 clknet_4_8_0_clk VGND VGND VPWR VPWR clkload8/X sky130_fd_sc_hd__clkbuf_8
XFILLER_137_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09819__A decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07234_ net1048 net6 net1057 net1052 VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__o211a_1
XANTENNA__11729__B1 _06243_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07165_ net1071 _02709_ _02710_ _02716_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_115_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout302_A _03849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1044_A net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07948__A2 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07096_ _02655_ _02656_ net952 _02654_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout1211_A net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12154__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13351__C1 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10704__A1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout671_A net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout769_A _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11295__S net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09806_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__inv_2
Xfanout278 _03873_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout289 _03860_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_2
X_07998_ net1143 _03508_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__nor2_1
X_09737_ _04430_ _04516_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12457__A1 net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06949_ _02526_ _02527_ _02529_ _02530_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_leaf_66_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout557_X net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09668_ _04465_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__nand2_1
XFILLER_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07802__A net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08619_ genblk1.genblk1.pcpi_mul.rd\[21\] genblk1.genblk1.pcpi_mul.next_rs2\[22\]
+ net1104 VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand3_1
X_09599_ reg_pc\[5\] net877 _04426_ net847 VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__a22o_1
XANTENNA__13015__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11630_ _06213_ _06216_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__nor2_1
XFILLER_30_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09625__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _02388_ mem_rdata_q\[13\] mem_rdata_q\[12\] VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__nor3_1
XANTENNA__12854__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13300_ net556 _02197_ _02217_ _02219_ net391 VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__a311o_1
XANTENNA__10640__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10512_ net987 decoded_imm\[4\] net858 VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a21o_1
X_14280_ clknet_leaf_100_clk _00734_ VGND VGND VPWR VPWR count_cycle\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11492_ instr_lh _02455_ _06156_ net3026 VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__a22o_1
XFILLER_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10882__B net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13231_ _04947_ _04959_ _04958_ _04948_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__a211o_1
X_10443_ cpuregs\[12\]\[0\] cpuregs\[13\]\[0\] net685 VGND VGND VPWR VPWR _05143_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11196__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12393__A0 _03751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13162_ net1396 net287 net433 VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__mux2_1
XFILLER_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10374_ _04879_ _05079_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__and2_1
XFILLER_163_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10943__A1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12113_ _06553_ _06554_ _06556_ net869 VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11994__A net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13093_ net296 net2335 net441 VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__mux2_1
XFILLER_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12145__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09010__A0 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12044_ net1015 _06496_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10403__A net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_X net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout790 net791 VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output221_A net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12448__A1 net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13995_ clknet_leaf_68_clk _00449_ VGND VGND VPWR VPWR cpuregs\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_148_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15734_ net1169 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
X_12946_ net356 net2434 net451 VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__mux2_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08367__X _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11505__Y _06163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ mem_rdata_q\[14\] net6 net962 VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__mux2_1
XFILLER_61_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14616_ clknet_leaf_93_clk _01002_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dfxtp_1
X_11828_ _06297_ _06298_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__nand2_1
X_15596_ clknet_leaf_180_clk _01932_ VGND VGND VPWR VPWR cpuregs\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12049__B net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07150__C net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14547_ clknet_leaf_24_clk _00933_ VGND VGND VPWR VPWR cpuregs\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11759_ net2548 net113 net729 VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__mux2_1
XANTENNA__11423__A2 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14478_ clknet_leaf_96_clk _00867_ VGND VGND VPWR VPWR instr_lbu sky130_fd_sc_hd__dfxtp_1
Xclkload103 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload103/Y sky130_fd_sc_hd__clkinv_4
Xclkload114 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload114/Y sky130_fd_sc_hd__bufinv_16
XPHY_EDGE_ROW_157_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload125 clknet_leaf_54_clk VGND VGND VPWR VPWR clkload125/Y sky130_fd_sc_hd__inv_6
X_13429_ net998 net393 _02331_ _02333_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__a22o_1
Xclkload136 clknet_leaf_69_clk VGND VGND VPWR VPWR clkload136/Y sky130_fd_sc_hd__bufinv_16
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload147 clknet_leaf_130_clk VGND VGND VPWR VPWR clkload147/Y sky130_fd_sc_hd__inv_6
Xclkload158 clknet_leaf_118_clk VGND VGND VPWR VPWR clkload158/Y sky130_fd_sc_hd__bufinv_16
Xclkload169 clknet_leaf_87_clk VGND VGND VPWR VPWR clkload169/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08052__B2 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08970_ genblk1.genblk1.pcpi_mul.rd\[23\] genblk1.genblk1.pcpi_mul.rd\[55\] net956
+ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07921_ _03294_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14430__D alu_out\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07852_ net258 net992 VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__and2_1
XFILLER_111_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06803_ net1006 VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__inv_2
Xinput1 mem_rdata[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_166_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07783_ _03298_ _03300_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__and2_1
XANTENNA__12939__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09304__A1 net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08107__A2 net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09522_ _04377_ _04378_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__nor2_1
XANTENNA__08277__X net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11111__A1 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09313__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09453_ _04332_ _04333_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__nor2_1
X_08404_ _03811_ _03814_ net767 VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__mux2_2
X_09384_ net1803 net322 net399 VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__mux2_1
XANTENNA__09607__A2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08335_ reg_pc\[3\] reg_pc\[2\] reg_pc\[4\] VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07618__A1 net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout1161_A net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_A net519 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08266_ reg_out\[10\] reg_next_pc\[10\] net921 VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__mux2_1
XFILLER_165_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07217_ net5 net22 net1048 VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__mux2_1
XANTENNA__06841__A2 reg_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08197_ _03465_ _03685_ _03681_ VGND VGND VPWR VPWR alu_out\[29\] sky130_fd_sc_hd__o21ai_2
XFILLER_134_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1047_X net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07148_ net1080 net1066 VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__nor2_2
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10925__A1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10207__B net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07079_ net1121 _02640_ genblk2.pcpi_div.dividend\[23\] VGND VGND VPWR VPWR _02642_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12127__B1 net993 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1214_X net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ count_cycle\[32\] count_cycle\[33\] count_cycle\[34\] _04821_ VGND VGND VPWR
+ VPWR _04826_ sky130_fd_sc_hd__and4_2
Xfanout1007 net1008 VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__clkbuf_4
Xfanout1018 net1019 VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__buf_4
Xfanout1029 net1030 VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__buf_2
XFILLER_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10223__A decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12849__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_X net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11753__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_12800_ net579 net1884 net465 VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__mux2_1
X_13780_ clknet_leaf_179_clk _00234_ VGND VGND VPWR VPWR cpuregs\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_10992_ _05656_ _05657_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__a21oi_4
XFILLER_55_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09223__S net495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11325__Y _05999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12731_ net1326 net884 _02099_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_26_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ clknet_leaf_42_clk _01789_ VGND VGND VPWR VPWR cpuregs\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07251__B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12662_ net1212 genblk1.genblk1.pcpi_mul.next_rs2\[30\] net905 net3003 _02080_ VGND
+ VGND VPWR VPWR _01335_ sky130_fd_sc_hd__a221o_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14401_ clknet_leaf_131_clk alu_out\[1\] VGND VGND VPWR VPWR alu_out_q\[1\] sky130_fd_sc_hd__dfxtp_1
X_11613_ is_alu_reg_imm mem_rdata_q\[30\] _06183_ _06199_ VGND VGND VPWR VPWR _06203_
+ sky130_fd_sc_hd__and4_1
XANTENNA__12584__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15381_ clknet_leaf_9_clk _01720_ VGND VGND VPWR VPWR cpuregs\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12593_ net322 net2215 net468 VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__mux2_1
XFILLER_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14332_ clknet_leaf_178_clk _06719_ VGND VGND VPWR VPWR reg_out\[12\] sky130_fd_sc_hd__dfxtp_1
X_11544_ net29 net28 net27 VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__or3b_1
XFILLER_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14263_ clknet_leaf_122_clk _00717_ VGND VGND VPWR VPWR count_cycle\[8\] sky130_fd_sc_hd__dfxtp_1
X_11475_ net1083 _06143_ net857 VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_59_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13214_ net569 _03189_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_94_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10426_ _02437_ _02491_ _05125_ _05128_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__nand4_1
X_14194_ clknet_leaf_132_clk _00648_ VGND VGND VPWR VPWR reg_pc\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13145_ net1946 net351 net431 VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__mux2_1
X_10357_ cpuregs\[17\]\[31\] net638 net613 _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__o211a_1
XANTENNA__12613__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08302__S net925 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13076_ net403 net1639 net440 VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _04914_ _04915_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__nand2b_1
XFILLER_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12027_ _06482_ _06481_ _06479_ net861 VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11663__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13978_ clknet_leaf_198_clk _00432_ VGND VGND VPWR VPWR cpuregs\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09133__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12929_ net175 net174 _06611_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__and3b_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15648_ clknet_leaf_34_clk _01984_ VGND VGND VPWR VPWR cpuregs\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08972__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13251__D1 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15579_ clknet_leaf_15_clk _01915_ VGND VGND VPWR VPWR cpuregs\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08120_ _03332_ net935 VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__nor2_1
XANTENNA__09470__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08051_ net770 _03554_ _03555_ _03551_ VGND VGND VPWR VPWR alu_out\[13\] sky130_fd_sc_hd__a31o_1
XFILLER_135_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07002_ net1118 _02575_ net2961 VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__a21oi_1
XFILLER_116_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap732 _06182_ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__buf_1
XANTENNA__10027__B net1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09773__A1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09308__S net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07617__A net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08953_ net2601 _04253_ net943 VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__mux2_1
XANTENNA__13338__B _05675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07904_ net1051 net1180 VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__and2b_1
XANTENNA__14511__Q decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1702 reg_sh\[0\] VGND VGND VPWR VPWR net3016 sky130_fd_sc_hd__dlygate4sd3_1
X_08884_ genblk1.genblk1.pcpi_mul.rd\[62\] genblk1.genblk1.pcpi_mul.next_rs2\[63\]
+ net1107 VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__nand3_1
Xhold1713 genblk1.genblk1.pcpi_mul.next_rs2\[30\] VGND VGND VPWR VPWR net3027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1724 count_cycle\[23\] VGND VGND VPWR VPWR net3038 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1007_A net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1735 net176 VGND VGND VPWR VPWR net3049 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07835_ net1168 net1033 VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__or2_1
XFILLER_84_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1746 count_instr\[37\] VGND VGND VPWR VPWR net3060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1757 genblk1.genblk1.pcpi_mul.next_rs2\[34\] VGND VGND VPWR VPWR net3071 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout467_A net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07766_ net1047 net1178 VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__or2_1
XANTENNA__09043__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09505_ net1226 _04366_ _04367_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__and3_1
X_07697_ net829 _03212_ _03214_ _03216_ net790 VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout634_A net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08167__B net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09436_ count_instr\[10\] _04320_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_140_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09367_ net1898 net577 net400 VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout801_A net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_X net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1164_X net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07498__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08318_ _03742_ _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__or2_4
X_09298_ net1894 net586 net481 VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__mux2_1
X_08249_ latched_branch latched_store VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__nand2_1
XANTENNA__14335__D _06722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1749_A decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10218__A decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11260_ cpuregs\[3\]\[25\] net642 net602 _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__o211a_1
XFILLER_119_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout791_X net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10211_ decoded_imm\[14\] net1022 VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__nand2_1
XANTENNA__11748__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11191_ _05866_ _05867_ net815 VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__mux2_1
XFILLER_134_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09218__S net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10142_ _04858_ _04859_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput190 net190 VGND VGND VPWR VPWR pcpi_insn[27] sky130_fd_sc_hd__buf_2
X_10073_ _04814_ _04815_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__nor2_1
X_14950_ clknet_leaf_34_clk _01302_ VGND VGND VPWR VPWR cpuregs\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11323__B2 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13901_ clknet_leaf_56_clk _00355_ VGND VGND VPWR VPWR cpuregs\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09742__A decoded_imm_j\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input28_A mem_rdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14881_ clknet_leaf_33_clk _01233_ VGND VGND VPWR VPWR cpuregs\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12579__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13264__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_57_clk _00286_ VGND VGND VPWR VPWR cpuregs\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13763_ clknet_leaf_15_clk _00217_ VGND VGND VPWR VPWR cpuregs\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_10975_ cpuregs\[22\]\[17\] cpuregs\[23\]\[17\] net646 VGND VGND VPWR VPWR _05658_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15502_ clknet_leaf_171_clk _01838_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dfxtp_1
X_12714_ net1192 genblk1.genblk1.pcpi_mul.next_rs1\[6\] net914 net1037 VGND VGND VPWR
+ VPWR _02091_ sky130_fd_sc_hd__a22o_1
XFILLER_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13694_ clknet_leaf_119_clk _00148_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15433_ clknet_leaf_22_clk _01772_ VGND VGND VPWR VPWR cpuregs\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12645_ net1202 genblk1.genblk1.pcpi_mul.next_rs2\[22\] net916 net248 VGND VGND VPWR
+ VPWR _02072_ sky130_fd_sc_hd__a22o_1
XFILLER_157_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15364_ clknet_leaf_38_clk _01703_ VGND VGND VPWR VPWR cpuregs\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12576_ net576 net2283 net468 VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__mux2_1
XFILLER_129_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14315_ clknet_leaf_101_clk _00769_ VGND VGND VPWR VPWR count_cycle\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11527_ mem_rdata_q\[20\] net2349 net736 VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__mux2_1
XFILLER_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15295_ clknet_leaf_66_clk _01636_ VGND VGND VPWR VPWR cpuregs\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold309 net41 VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ clknet_leaf_75_clk _00700_ VGND VGND VPWR VPWR reg_next_pc\[23\] sky130_fd_sc_hd__dfxtp_1
X_11458_ _06126_ _06127_ net805 VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11658__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10409_ net250 net1158 _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__or3_2
X_14177_ clknet_leaf_109_clk _00631_ VGND VGND VPWR VPWR count_instr\[48\] sky130_fd_sc_hd__dfxtp_1
X_11389_ cpuregs\[22\]\[28\] cpuregs\[23\]\[28\] net688 VGND VGND VPWR VPWR _06061_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12343__A mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13128_ net286 net2399 net437 VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__mux2_1
XANTENNA__07230__A2 decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13059_ net1646 net82 net533 VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1009 cpuregs\[7\]\[5\] VGND VGND VPWR VPWR net2323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08967__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09652__A net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08191__B1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07620_ net1080 decoded_imm_j\[16\] VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__or2_1
XFILLER_38_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ count_instr\[59\] net1133 net1141 count_cycle\[59\] VGND VGND VPWR VPWR _03077_
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15162__Q mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07482_ count_instr\[54\] net1133 net1141 count_cycle\[54\] VGND VGND VPWR VPWR _03013_
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09221_ net1997 net307 net494 VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__mux2_1
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10737__S net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13113__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08246__A1 net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09152_ net1509 net318 net501 VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__mux2_1
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08103_ net1144 _03337_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__nor2_1
XANTENNA__12952__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09083_ net1395 net312 net510 VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__mux2_1
XANTENNA__10038__A _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08034_ _03535_ _03540_ VGND VGND VPWR VPWR alu_out\[11\] sky130_fd_sc_hd__nand2_1
Xhold810 cpuregs\[31\]\[29\] VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 cpuregs\[4\]\[8\] VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold832 cpuregs\[18\]\[21\] VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 cpuregs\[19\]\[11\] VGND VGND VPWR VPWR net2157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_171_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13349__A _02408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold854 cpuregs\[17\]\[29\] VGND VGND VPWR VPWR net2168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold865 cpuregs\[5\]\[25\] VGND VGND VPWR VPWR net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 cpuregs\[29\]\[19\] VGND VGND VPWR VPWR net2190 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09038__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold887 cpuregs\[23\]\[20\] VGND VGND VPWR VPWR net2201 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__B1 net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold898 cpuregs\[17\]\[2\] VGND VGND VPWR VPWR net2212 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09985_ _04451_ _04748_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__nor2_1
XFILLER_89_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout584_A _03751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08936_ genblk1.genblk1.pcpi_mul.rd\[6\] genblk1.genblk1.pcpi_mul.rd\[38\] net955
+ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__mux2_1
XFILLER_76_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_186_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1510 count_cycle\[46\] VGND VGND VPWR VPWR net2824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 _06592_ VGND VGND VPWR VPWR net2835 sky130_fd_sc_hd__dlygate4sd3_1
X_08867_ _04195_ _04198_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__nand2_1
XANTENNA__12399__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1532 _01357_ VGND VGND VPWR VPWR net2846 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout372_X net372 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A _05120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1543 count_cycle\[3\] VGND VGND VPWR VPWR net2857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 _01065_ VGND VGND VPWR VPWR net2868 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12700__B net912 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1565 genblk2.pcpi_div.quotient_msk\[31\] VGND VGND VPWR VPWR net2879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1576 genblk1.genblk1.pcpi_mul.next_rs2\[16\] VGND VGND VPWR VPWR net2890 sky130_fd_sc_hd__dlygate4sd3_1
X_07818_ net1159 net1012 VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__xor2_2
XANTENNA__13058__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08798_ net889 _04141_ _04143_ net2576 net1195 VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__a32o_1
Xhold1587 _01363_ VGND VGND VPWR VPWR net2901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 instr_sb VGND VGND VPWR VPWR net2912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11069__B1 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07749_ net255 net996 VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__or2_1
XANTENNA__10220__B net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10760_ net813 _05446_ _05448_ net828 VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__o211a_1
XFILLER_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07810__A net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09419_ _04310_ net1231 _04309_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__and3b_1
XFILLER_139_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10691_ cpuregs\[17\]\[9\] net627 net607 _05381_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout804_X net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13023__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12430_ genblk1.genblk1.pcpi_mul.mul_counter\[2\] _06666_ genblk1.genblk1.pcpi_mul.mul_counter\[3\]
+ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__o21a_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08237__A1 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10044__A1 _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12361_ net1376 net578 net361 VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__mux2_1
XFILLER_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12862__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14100_ clknet_leaf_178_clk _00554_ VGND VGND VPWR VPWR cpuregs\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07996__B1 net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11312_ cpuregs\[24\]\[26\] net703 VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__or2_1
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15080_ clknet_leaf_103_clk _01432_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12292_ decoded_imm\[27\] net733 VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_91_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14031_ clknet_leaf_45_clk _00485_ VGND VGND VPWR VPWR cpuregs\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11243_ net804 _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__or2_1
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11174_ cpuregs\[19\]\[22\] net633 net597 VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__o21a_1
XFILLER_80_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10125_ count_cycle\[47\] _04846_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__and2_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10056_ count_cycle\[20\] count_cycle\[21\] count_cycle\[22\] _04798_ VGND VGND VPWR
+ VPWR _04804_ sky130_fd_sc_hd__and4_1
X_14933_ clknet_leaf_181_clk _01285_ VGND VGND VPWR VPWR cpuregs\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13049__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10411__A net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14864_ clknet_leaf_182_clk _01216_ VGND VGND VPWR VPWR cpuregs\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13815_ clknet_leaf_182_clk _00269_ VGND VGND VPWR VPWR cpuregs\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14795_ clknet_leaf_67_clk _01147_ VGND VGND VPWR VPWR decoded_imm\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13746_ clknet_leaf_29_clk _00200_ VGND VGND VPWR VPWR cpuregs\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_10958_ cpuregs\[4\]\[17\] cpuregs\[5\]\[17\] net659 VGND VGND VPWR VPWR _05641_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13441__B _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07684__C1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13677_ clknet_leaf_147_clk _00131_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_10889_ cpuregs\[14\]\[15\] cpuregs\[15\]\[15\] net647 VGND VGND VPWR VPWR _05574_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ net2830 net886 _02063_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__a21o_1
X_15416_ clknet_leaf_11_clk _01755_ VGND VGND VPWR VPWR cpuregs\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08228__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08228__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13221__B2 net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09976__A1 net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15347_ clknet_leaf_12_clk _01687_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
X_12559_ net2553 net389 _02040_ _02041_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__a22o_1
XANTENNA__10586__A2 decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15278_ clknet_leaf_198_clk _01619_ VGND VGND VPWR VPWR cpuregs\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold106 cpuregs\[14\]\[22\] VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 cpuregs\[14\]\[3\] VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold128 cpuregs\[30\]\[23\] VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 cpuregs\[29\]\[13\] VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ clknet_leaf_174_clk _00683_ VGND VGND VPWR VPWR reg_next_pc\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_146_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 net609 VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_2
XANTENNA__15157__Q mem_rdata_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout619 net620 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ _04543_ _04549_ _04558_ net1149 VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__o31a_1
XFILLER_113_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06982_ net951 _02557_ _02558_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__or3_1
XFILLER_140_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08721_ genblk1.genblk1.pcpi_mul.next_rs2\[38\] net1099 genblk1.genblk1.pcpi_mul.rd\[37\]
+ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_124_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13108__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1190 net1191 VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ _04018_ _04019_ _04013_ _04016_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_87_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10510__A2 decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07603_ reg_pc\[30\] decoded_imm\[30\] _03115_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__a21oi_1
X_08583_ net1196 net2880 net890 _03961_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__a22o_1
XFILLER_42_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12947__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07534_ _03047_ _03049_ _03060_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__a21o_1
XANTENNA__12263__A2 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08285__X net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09321__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07465_ _02994_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__nand2_1
XFILLER_23_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09204_ net1897 net525 net492 VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13212__A1 reg_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07396_ count_instr\[48\] net1132 net1140 count_cycle\[48\] VGND VGND VPWR VPWR _02933_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08219__B2 net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09135_ net1825 net573 net501 VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__mux2_1
XANTENNA__11223__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10991__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11774__A1 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09066_ net1361 net543 net511 VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__mux2_1
XFILLER_162_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08017_ net770 _03525_ _03520_ VGND VGND VPWR VPWR alu_out\[9\] sky130_fd_sc_hd__a21o_1
XANTENNA_fanout799_A net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold640 cpuregs\[4\]\[15\] VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 net138 VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold662 cpuregs\[2\]\[13\] VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold673 cpuregs\[2\]\[22\] VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 instr_beq VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold695 cpuregs\[8\]\[16\] VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout966_A net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10215__B net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09968_ _04723_ _04725_ _04732_ _04740_ _04724_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__a311o_1
X_08919_ net1203 net2708 net895 _04236_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__a22o_1
XANTENNA__08400__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09899_ _04677_ _04678_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__xnor2_1
Xhold1340 instr_slt VGND VGND VPWR VPWR net2654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13018__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1351 genblk1.genblk1.pcpi_mul.rdx\[60\] VGND VGND VPWR VPWR net2665 sky130_fd_sc_hd__dlygate4sd3_1
X_11930_ _06259_ _06393_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__nor2_1
Xhold1362 genblk1.genblk1.pcpi_mul.rd\[44\] VGND VGND VPWR VPWR net2676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10231__A decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1373 genblk2.pcpi_div.divisor\[42\] VGND VGND VPWR VPWR net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 net154 VGND VGND VPWR VPWR net2698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1395 genblk1.genblk1.pcpi_mul.mul_counter\[2\] VGND VGND VPWR VPWR net2709 sky130_fd_sc_hd__dlygate4sd3_1
X_11861_ _06329_ _06330_ _06307_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout921_X net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12857__S net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11761__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13600_ clknet_leaf_24_clk _00055_ VGND VGND VPWR VPWR cpuregs\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10812_ cpuregs\[1\]\[13\] net549 _05498_ net799 net823 VGND VGND VPWR VPWR _05499_
+ sky130_fd_sc_hd__a221o_1
X_14580_ clknet_leaf_69_clk net1466 VGND VGND VPWR VPWR latched_rd\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12254__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11792_ genblk2.pcpi_div.divisor\[29\] genblk2.pcpi_div.dividend\[29\] VGND VGND
+ VPWR VPWR _06263_ sky130_fd_sc_hd__nand2b_1
XANTENNA__13451__B2 is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09231__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07540__A _02702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13531_ net404 net2019 net416 VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__mux2_1
XFILLER_43_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10743_ cpuregs\[22\]\[11\] cpuregs\[23\]\[11\] net664 VGND VGND VPWR VPWR _05432_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13462_ net1710 net526 net424 VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__mux2_1
X_10674_ cpuregs\[9\]\[9\] net628 net607 _05364_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__o211a_1
XANTENNA__13203__A1 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1280 VGND VGND VPWR VPWR picorv32_1280/HI trace_data[2] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15201_ clknet_leaf_15_clk _01550_ VGND VGND VPWR VPWR cpuregs\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12413_ net317 net1919 net474 VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1291 VGND VGND VPWR VPWR picorv32_1291/HI trace_data[13] sky130_fd_sc_hd__conb_1
XANTENNA__12592__S net470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13393_ net558 _02277_ _02301_ net566 reg_pc\[23\] VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__a32o_1
XFILLER_138_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15132_ clknet_leaf_1_clk _01484_ VGND VGND VPWR VPWR cpuregs\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12344_ net1151 decoded_imm_j\[3\] _06617_ mem_rdata_q\[10\] net734 VGND VGND VPWR
+ VPWR _06653_ sky130_fd_sc_hd__a221o_1
X_15063_ clknet_leaf_104_clk _01415_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12275_ net2760 _06613_ _06615_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__a21bo_1
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10406__A net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14014_ clknet_leaf_10_clk _00468_ VGND VGND VPWR VPWR cpuregs\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12714__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11226_ cpuregs\[20\]\[24\] cpuregs\[21\]\[24\] net687 VGND VGND VPWR VPWR _05902_
+ sky130_fd_sc_hd__mux2_1
XFILLER_134_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output251_A net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11936__S net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11157_ cpuregs\[10\]\[22\] net682 VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__or2_1
XANTENNA__06944__A1 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10108_ _04836_ _04837_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__nor2_1
X_11088_ cpuregs\[6\]\[20\] cpuregs\[7\]\[20\] net661 VGND VGND VPWR VPWR _05768_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12340__B _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10039_ count_cycle\[16\] _04791_ net1206 VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__a21oi_1
X_14916_ clknet_leaf_111_clk _01268_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12493__A2 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14847_ clknet_leaf_31_clk _01199_ VGND VGND VPWR VPWR cpuregs\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12245__A2 net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14778_ clknet_leaf_154_clk _00033_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09141__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11453__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13729_ clknet_leaf_116_clk _00183_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_07250_ _02790_ _02794_ net991 VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08980__S net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07181_ _02710_ _02724_ _02723_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__o21ai_1
XFILLER_118_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08082__C1 net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10964__C1 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout405 _03785_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10035__B net1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout416 _02357_ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_2
Xfanout427 net428 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_4
X_09822_ _04592_ _04597_ _04606_ _04590_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__o211a_1
Xfanout438 _02126_ VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__buf_4
XANTENNA__06800__Y _02408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout449 net450 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09316__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09753_ decoded_imm_j\[11\] _04432_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__nor2_1
X_06965_ genblk2.pcpi_div.quotient\[4\] genblk2.pcpi_div.quotient\[5\] genblk2.pcpi_div.quotient\[6\]
+ _02525_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__or4_1
X_08704_ _04062_ _04063_ _04057_ _04060_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__a211o_1
X_09684_ net2740 net878 _04479_ _04481_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__a22o_1
X_06896_ is_lb_lh_lw_lbu_lhu _02436_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__and2_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09840__A net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08635_ net1210 net2897 net899 _04005_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__a22o_1
XANTENNA__10495__A1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ genblk1.genblk1.pcpi_mul.rd\[13\] genblk1.genblk1.pcpi_mul.next_rs2\[14\]
+ net1093 VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__and3_1
XANTENNA__13433__A1 net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09051__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07517_ net1073 _03037_ _03038_ _03045_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__a31o_1
XANTENNA__11444__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08497_ _03882_ net761 _03886_ _03887_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout714_A _02083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10798__A2 net620 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07448_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10992__Y _05675_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07379_ count_instr\[15\] net1136 net977 _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__a211o_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout502_X net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12944__A0 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09118_ net1702 net305 net507 VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__mux2_1
XANTENNA__07359__X _02898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ _02362_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nor2_1
XFILLER_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09049_ net314 net2329 net514 VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__mux2_1
XANTENNA__10226__A decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12060_ net867 _06509_ _06510_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__and3_1
Xhold470 cpuregs\[28\]\[16\] VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold481 cpuregs\[16\]\[4\] VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__A1 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_X net969 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07179__B2 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold492 cpuregs\[13\]\[12\] VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net779 _05683_ _05692_ net776 VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__o211a_1
XANTENNA__11756__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10183__B1 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12441__A net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11380__C1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09226__S net495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout950 net952 VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__buf_2
XFILLER_49_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout961 _02462_ VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__clkbuf_4
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13256__B _05316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout972 net975 VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout983 _02416_ VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout994 net995 VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__clkbuf_4
XFILLER_18_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12962_ net293 net2227 net453 VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__mux2_1
Xhold1170 cpuregs\[17\]\[28\] VGND VGND VPWR VPWR net2484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A mem_rdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11913_ _06265_ _06383_ _06264_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__o21ba_1
X_14701_ clknet_leaf_163_clk _01086_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10486__A1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1181 cpuregs\[3\]\[28\] VGND VGND VPWR VPWR net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 cpuregs\[18\]\[31\] VGND VGND VPWR VPWR net2506 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ mem_rdata_q\[30\] net24 net965 VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__mux2_1
XFILLER_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12587__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07351__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13272__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14632_ clknet_leaf_170_clk _01017_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_11844_ genblk2.pcpi_div.divisor\[3\] genblk2.pcpi_div.dividend\[3\] VGND VGND VPWR
+ VPWR _06315_ sky130_fd_sc_hd__nand2b_1
XFILLER_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12227__A2 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13424__A1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14563_ clknet_leaf_14_clk _00949_ VGND VGND VPWR VPWR cpuregs\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11775_ _06245_ _06249_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__and2_1
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08313__A1_N net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13514_ net1726 net299 net421 VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__mux2_1
X_10726_ cpuregs\[16\]\[10\] net668 VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__or2_1
X_14494_ clknet_leaf_94_clk _00883_ VGND VGND VPWR VPWR instr_slt sky130_fd_sc_hd__dfxtp_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13445_ _02343_ _02344_ _02347_ net397 net994 VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__o32a_1
X_10657_ cpuregs\[18\]\[8\] net553 _05348_ net780 VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__o22a_1
XANTENNA__11738__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload15/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__07269__X _02814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload26 clknet_leaf_178_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__bufinv_16
Xclkload37 clknet_leaf_190_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__bufinv_16
X_13376_ net558 _02262_ _02284_ _02286_ net393 VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__a311o_1
XANTENNA__08305__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10588_ cpuregs\[6\]\[7\] cpuregs\[7\]\[7\] net673 VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__mux2_1
Xclkload48 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__clkinv_4
XFILLER_170_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload59 clknet_leaf_176_clk VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__clkinv_4
XFILLER_115_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12327_ net744 _06618_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__and2_1
X_15115_ clknet_leaf_46_clk _01467_ VGND VGND VPWR VPWR cpuregs\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15046_ clknet_leaf_112_clk _01398_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_12258_ net2731 net377 net364 net2816 VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__a22o_1
XFILLER_123_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13447__A net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11209_ cpuregs\[10\]\[23\] net662 VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_79_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12189_ genblk2.pcpi_div.quotient_msk\[8\] net274 net2933 VGND VGND VPWR VPWR _06587_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_69_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09136__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10477__B2 net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08420_ reg_out\[21\] alu_out_q\[21\] net1155 VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__mux2_1
XFILLER_52_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11414__B net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08351_ reg_pc\[7\] reg_pc\[6\] _03764_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__and3_1
XANTENNA__15170__Q mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14428__D alu_out\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07302_ net1063 net1029 _02844_ net1077 _02840_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ reg_out\[18\] reg_next_pc\[18\] net922 VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07645__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload9 clknet_4_9_0_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_12
X_07233_ _02774_ _02776_ _02778_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__a21o_1
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10745__S net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13121__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07164_ net1062 _02708_ _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_132_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14514__Q decoded_imm_j\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07095_ net1122 genblk2.pcpi_div.quotient\[25\] _02651_ net952 VGND VGND VPWR VPWR
+ _02656_ sky130_fd_sc_hd__a31o_1
XANTENNA__07339__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12960__S net454 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout497_A net499 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1204_A net1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09046__S net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A mem_rdata[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09805_ _04590_ _04591_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__nand2_1
XANTENNA__08189__A2_N net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout279 _03873_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_1
X_07997_ _03280_ _03501_ _03282_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout664_A net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ _04516_ _04430_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__nand2b_1
X_06948_ genblk2.pcpi_div.dividend\[4\] net1125 _02528_ net949 VGND VGND VPWR VPWR
+ _02530_ sky130_fd_sc_hd__a31o_1
XANTENNA__10468__A1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09667_ decoded_imm_j\[1\] _04422_ _04457_ _04456_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout452_X net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06879_ net1066 _02474_ _02476_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__and3_1
XFILLER_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08618_ genblk1.genblk1.pcpi_mul.rd\[21\] genblk1.genblk1.pcpi_mul.next_rs2\[22\]
+ net1104 VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__and3_1
XANTENNA__07802__B net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08186__A net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09598_ _03762_ reg_next_pc\[5\] net923 VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__mux2_1
XFILLER_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08549_ _03925_ _03928_ _03930_ _03931_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__o211a_1
XFILLER_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11560_ net3018 net561 _06178_ _06180_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__a22o_1
XANTENNA__12090__B1 net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10511_ net1176 net860 _05207_ _03228_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__o22a_1
XFILLER_155_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ _02370_ net1061 _02454_ mem_do_rdata net1232 VGND VGND VPWR VPWR _06156_
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13031__S net446 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13230_ _03263_ net568 VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__nor2_1
XFILLER_155_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10442_ net831 _05137_ _05139_ _05141_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__a211o_1
XFILLER_152_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13161_ net2389 net290 net434 VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__mux2_1
XFILLER_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10373_ instr_lui is_lui_auipc_jal VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__and2b_1
XFILLER_123_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12112_ net999 _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__xnor2_1
XFILLER_163_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13092_ net299 net1985 net441 VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__mux2_1
XFILLER_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12043_ net1016 _06492_ net721 VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_57_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07572__A1 net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout780 net781 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07572__B2 net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout791 net795 VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12448__A2 net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13994_ clknet_leaf_45_clk _00448_ VGND VGND VPWR VPWR cpuregs\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input13_X net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15733_ net125 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_1
XFILLER_45_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12945_ net403 net2142 net451 VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__mux2_1
XFILLER_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output214_A net1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11120__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ mem_rdata_q\[13\] net5 net963 VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__mux2_1
XFILLER_61_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14615_ clknet_leaf_115_clk _01001_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dfxtp_1
X_11827_ genblk2.pcpi_div.dividend\[12\] genblk2.pcpi_div.divisor\[12\] VGND VGND
+ VPWR VPWR _06298_ sky130_fd_sc_hd__nand2b_1
X_15595_ clknet_leaf_21_clk _01931_ VGND VGND VPWR VPWR cpuregs\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12049__C net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12081__B1 net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14546_ clknet_leaf_21_clk _00932_ VGND VGND VPWR VPWR cpuregs\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11758_ net1520 net112 net728 VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10709_ cpuregs\[8\]\[10\] net666 VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__or2_1
XANTENNA__10631__B2 net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14477_ clknet_leaf_95_clk _00866_ VGND VGND VPWR VPWR instr_lw sky130_fd_sc_hd__dfxtp_1
X_11689_ net1854 net542 net374 VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__mux2_1
XANTENNA__12346__A mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload104 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload104/Y sky130_fd_sc_hd__inv_6
X_13428_ _04879_ _02332_ net393 VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__a21oi_1
Xclkload115 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload115/X sky130_fd_sc_hd__clkbuf_4
Xclkload126 clknet_leaf_55_clk VGND VGND VPWR VPWR clkload126/Y sky130_fd_sc_hd__clkinv_8
Xclkload137 clknet_leaf_70_clk VGND VGND VPWR VPWR clkload137/Y sky130_fd_sc_hd__inv_12
XANTENNA__11187__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload148 clknet_leaf_131_clk VGND VGND VPWR VPWR clkload148/X sky130_fd_sc_hd__clkbuf_8
Xclkload159 clknet_leaf_119_clk VGND VGND VPWR VPWR clkload159/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13359_ net557 _02247_ _02271_ net565 reg_pc\[19\] VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__a32o_1
XFILLER_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13333__B1 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07920_ _03335_ _03348_ _03437_ _03408_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__o31a_1
X_15029_ clknet_leaf_137_clk _01381_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11344__C1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07851_ _03368_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__inv_2
XANTENNA__10698__A1 net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15165__Q mem_rdata_q\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06802_ net1009 VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__inv_2
XFILLER_96_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 mem_rdata[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
X_07782_ net1164 net1026 VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__or2_1
XFILLER_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11647__A0 decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09521_ net2796 _04376_ net1226 VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13116__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09452_ net3042 _04330_ net1228 VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08403_ _03812_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__nor2_1
XANTENNA__14509__Q decoded_imm_j\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09068__A1 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09383_ net2226 net325 net401 VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__mux2_1
XANTENNA__12955__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08334_ reg_pc\[4\] reg_pc\[3\] reg_pc\[2\] VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__and3_1
XANTENNA__07618__A2 decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08293__X net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08265_ net1031 _03716_ net980 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__mux2_1
XANTENNA_fanout412_A _02358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1154_A net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07216_ _02761_ _02762_ _02760_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__a21o_1
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08196_ _03314_ _03684_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07147_ count_instr\[0\] net1135 net977 _02699_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__a211o_1
XFILLER_145_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07078_ genblk2.pcpi_div.dividend\[23\] net1121 _02640_ VGND VGND VPWR VPWR _02641_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout781_A net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A net880 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13324__B1 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10138__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1008 net217 VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__buf_4
Xfanout1019 net210 VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1207_X net1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input5_X net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07554__A1 genblk2.pcpi_div.pcpi_rd\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10223__B net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07813__A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09719_ _04511_ _04512_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__and2b_1
X_10991_ net772 _05665_ _05673_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__and3_1
XANTENNA__13026__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12730_ net1190 genblk1.genblk1.pcpi_mul.next_rs1\[14\] net914 net1021 VGND VGND
+ VPWR VPWR _02099_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _02398_ net913 VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__nor2_1
X_11612_ net3005 net563 _06185_ _06201_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__a22o_1
X_14400_ clknet_leaf_127_clk alu_out\[0\] VGND VGND VPWR VPWR alu_out_q\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_169_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15380_ clknet_leaf_10_clk _01719_ VGND VGND VPWR VPWR cpuregs\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12592_ net327 net2425 net470 VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__mux2_1
XANTENNA__10613__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11543_ net2557 _06168_ net547 VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__mux2_1
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14331_ clknet_leaf_177_clk _06718_ VGND VGND VPWR VPWR reg_out\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14262_ clknet_leaf_122_clk _00716_ VGND VGND VPWR VPWR count_cycle\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11474_ net1083 decoded_imm\[30\] VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__or2_1
XFILLER_125_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12366__A1 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13213_ _02136_ _02142_ _02143_ net397 net1047 VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__o32a_1
X_10425_ net1087 is_sb_sh_sw mem_do_prefetch VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14193_ clknet_leaf_132_clk _00647_ VGND VGND VPWR VPWR reg_pc\[1\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_94_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10916__A2 _05599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13144_ net1409 net357 net431 VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__mux2_1
XFILLER_152_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10356_ cpuregs\[16\]\[31\] net692 VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__or2_1
XFILLER_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12613__B net1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13075_ net407 net1631 net439 VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__mux2_1
X_10287_ decoded_imm\[17\] net1017 net1018 decoded_imm\[16\] VGND VGND VPWR VPWR _04993_
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ net1021 net721 _06480_ net861 VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__a31o_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08378__X _03794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13977_ clknet_leaf_191_clk _00431_ VGND VGND VPWR VPWR cpuregs\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12928_ net174 _06611_ net175 VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__and3b_1
XFILLER_62_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15647_ clknet_leaf_71_clk _01983_ VGND VGND VPWR VPWR cpuregs\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12859_ net289 net2383 net461 VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__mux2_1
XANTENNA__12054__B1 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15578_ clknet_leaf_12_clk _01914_ VGND VGND VPWR VPWR cpuregs\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14529_ clknet_leaf_80_clk _00918_ VGND VGND VPWR VPWR decoded_imm_j\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08050_ _03288_ _03553_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07001_ genblk2.pcpi_div.quotient\[11\] _02565_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__or2_1
XFILLER_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06802__A net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11580__A2 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08952_ genblk1.genblk1.pcpi_mul.rd\[14\] genblk1.genblk1.pcpi_mul.rd\[46\] net954
+ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__mux2_1
XFILLER_88_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07617__B decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07903_ net1178 net1049 VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__nand2b_1
X_08883_ genblk1.genblk1.pcpi_mul.next_rs2\[63\] net1107 genblk1.genblk1.pcpi_mul.rd\[62\]
+ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__a21o_1
Xhold1703 reg_next_pc\[25\] VGND VGND VPWR VPWR net3017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07536__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1714 count_instr\[2\] VGND VGND VPWR VPWR net3028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1725 count_cycle\[4\] VGND VGND VPWR VPWR net3039 sky130_fd_sc_hd__dlygate4sd3_1
X_07834_ net1168 net1033 VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__nand2_1
Xhold1736 genblk2.pcpi_div.dividend\[23\] VGND VGND VPWR VPWR net3050 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1747 reg_pc\[16\] VGND VGND VPWR VPWR net3061 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1758 genblk2.pcpi_div.quotient_msk\[27\] VGND VGND VPWR VPWR net3072 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10978__B net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09324__S net482 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07765_ _03281_ _03282_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout362_A net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08159__A1_N net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09504_ count_instr\[33\] count_instr\[32\] _04363_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__nand3_1
X_07696_ cpuregs\[27\]\[3\] net629 net595 _03215_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__o211a_1
XFILLER_112_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10843__A1 net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09435_ _04320_ _04321_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__nor2_1
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout627_A net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09366_ net1737 net581 net402 VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__mux2_1
XANTENNA__13242__C1 _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11399__A2 _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08317_ latched_rd\[0\] _03743_ latched_rd\[1\] VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__or3b_4
X_09297_ latched_rd\[1\] latched_rd\[0\] _04289_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__nor3_2
XANTENNA_fanout415_X net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_X net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08248_ net1157 net940 _03707_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__a21o_1
XANTENNA_fanout996_A net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10218__B net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08179_ _03443_ _03669_ net990 VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__mux2_1
XFILLER_107_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10210_ decoded_imm\[15\] net1020 VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__nor2_1
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07808__A net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11190_ cpuregs\[20\]\[23\] cpuregs\[21\]\[23\] net697 VGND VGND VPWR VPWR _05867_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout784_X net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10141_ net3001 _04856_ net1235 VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__o21ai_1
XFILLER_134_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10234__A decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput180 net180 VGND VGND VPWR VPWR pcpi_insn[18] sky130_fd_sc_hd__buf_2
XANTENNA__11308__C1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput191 net191 VGND VGND VPWR VPWR pcpi_insn[28] sky130_fd_sc_hd__buf_2
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10072_ net2987 _04813_ net1236 VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__o21ai_1
XFILLER_88_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07527__A1 genblk2.pcpi_div.pcpi_rd\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11764__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11323__A2 net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13900_ clknet_leaf_54_clk _00354_ VGND VGND VPWR VPWR cpuregs\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_14880_ clknet_leaf_72_clk _01232_ VGND VGND VPWR VPWR cpuregs\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09234__S net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13264__B _05351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13831_ clknet_leaf_71_clk _00285_ VGND VGND VPWR VPWR cpuregs\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07262__B decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10974_ _05644_ _05647_ _03171_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__o21a_1
X_13762_ clknet_leaf_14_clk _00216_ VGND VGND VPWR VPWR cpuregs\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15501_ clknet_leaf_174_clk _01837_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dfxtp_2
X_12713_ net1364 net883 _02090_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__a21o_1
XFILLER_71_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12595__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13693_ clknet_leaf_105_clk _00147_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13280__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15432_ clknet_leaf_29_clk _01771_ VGND VGND VPWR VPWR cpuregs\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12644_ net2763 net895 _02071_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__a21o_1
XFILLER_129_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15363_ clknet_leaf_102_clk genblk1.genblk1.pcpi_mul.instr_any_mul VGND VGND VPWR
+ VPWR genblk1.genblk1.pcpi_mul.pcpi_wait sky130_fd_sc_hd__dfxtp_1
X_12575_ net580 net2319 net469 VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__mux2_1
XANTENNA__10409__A net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14314_ clknet_leaf_101_clk _00768_ VGND VGND VPWR VPWR count_cycle\[59\] sky130_fd_sc_hd__dfxtp_1
X_11526_ mem_rdata_q\[19\] net2101 net742 VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__mux2_1
X_15294_ clknet_leaf_51_clk _01635_ VGND VGND VPWR VPWR cpuregs\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12339__A1 decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12339__B2 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11457_ cpuregs\[22\]\[30\] cpuregs\[23\]\[30\] net689 VGND VGND VPWR VPWR _06127_
+ sky130_fd_sc_hd__mux2_1
X_14245_ clknet_leaf_76_clk _00699_ VGND VGND VPWR VPWR reg_next_pc\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10180__D_N net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11011__A1 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10408_ net248 _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__or2_1
X_14176_ clknet_leaf_111_clk _00630_ VGND VGND VPWR VPWR count_instr\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11388_ net832 _06055_ _06057_ _06059_ net793 VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__a2111o_1
XANTENNA_output89_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10415__Y _05120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12343__B _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10339_ cpuregs\[1\]\[31\] net639 net613 _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__o211a_1
X_13127_ net290 net2509 net437 VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__mux2_1
XFILLER_98_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13058_ net1373 net81 net536 VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__mux2_1
XANTENNA__09933__A _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12009_ genblk2.pcpi_div.dividend\[12\] _06467_ net271 VGND VGND VPWR VPWR _01021_
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09144__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07550_ net20 net938 net937 VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11078__A1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07481_ net15 net938 net936 VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_122_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09220_ net1993 net310 net494 VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__mux2_1
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07900__B net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09151_ net1875 net323 net501 VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__mux2_1
XANTENNA__11422__B net707 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08102_ _03338_ _03593_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__or2_1
XFILLER_159_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07454__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09082_ net1704 net316 net510 VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__mux2_1
XFILLER_163_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13527__A0 net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08033_ _03364_ _03538_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a21o_1
XANTENNA__10753__S net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold800 cpuregs\[3\]\[3\] VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 cpuregs\[2\]\[29\] VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 cpuregs\[25\]\[26\] VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09319__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold833 cpuregs\[19\]\[18\] VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 cpuregs\[13\]\[27\] VGND VGND VPWR VPWR net2158 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13349__B net759 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold855 cpuregs\[5\]\[29\] VGND VGND VPWR VPWR net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 cpuregs\[17\]\[13\] VGND VGND VPWR VPWR net2180 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__A1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold877 cpuregs\[23\]\[0\] VGND VGND VPWR VPWR net2191 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__B2 net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold888 cpuregs\[3\]\[8\] VGND VGND VPWR VPWR net2202 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09984_ net1152 _04755_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__nand2_1
Xhold899 cpuregs\[11\]\[16\] VGND VGND VPWR VPWR net2213 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1117_A net1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08935_ net2539 _04244_ net944 VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout577_A _03756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1500 genblk1.genblk1.pcpi_mul.next_rs2\[15\] VGND VGND VPWR VPWR net2814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 count_instr\[21\] VGND VGND VPWR VPWR net2825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13365__A net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1522 count_instr\[42\] VGND VGND VPWR VPWR net2836 sky130_fd_sc_hd__dlygate4sd3_1
X_08866_ _04199_ _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nand2_1
Xhold1533 genblk2.pcpi_div.quotient_msk\[30\] VGND VGND VPWR VPWR net2847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08182__A1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1544 genblk2.pcpi_div.quotient_msk\[3\] VGND VGND VPWR VPWR net2858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09054__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1555 genblk1.genblk1.pcpi_mul.rd\[37\] VGND VGND VPWR VPWR net2869 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1566 genblk1.genblk1.pcpi_mul.rd\[15\] VGND VGND VPWR VPWR net2880 sky130_fd_sc_hd__dlygate4sd3_1
X_07817_ _03323_ _03327_ _03330_ _03333_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__or4_1
Xhold1577 genblk2.pcpi_div.divisor\[30\] VGND VGND VPWR VPWR net2891 sky130_fd_sc_hd__dlygate4sd3_1
X_08797_ _04142_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__inv_2
Xhold1588 genblk1.genblk1.pcpi_mul.next_rs2\[6\] VGND VGND VPWR VPWR net2902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_A net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1599 genblk1.genblk1.pcpi_mul.rd\[47\] VGND VGND VPWR VPWR net2913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11069__A1 cpu_state\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07748_ net255 net996 VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__nand2_1
XANTENNA__07650__X _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout911_A net913 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07679_ net801 _03197_ net549 cpuregs\[1\]\[3\] net829 VGND VGND VPWR VPWR _03199_
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12018__B1 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07810__B net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09418_ count_instr\[4\] _04307_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__and2_1
X_10690_ cpuregs\[16\]\[9\] net671 VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_33_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09349_ net1655 net330 net475 VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__mux2_1
XANTENNA__10229__A decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12360_ net1387 net582 net362 VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__mux2_1
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11759__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11311_ _05983_ _05984_ net807 VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout999_X net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07996__A1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12291_ mem_rdata_q\[28\] _06622_ _06624_ _06620_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__a211o_1
XANTENNA__11986__C net1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14030_ clknet_leaf_39_clk _00484_ VGND VGND VPWR VPWR cpuregs\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11242_ cpuregs\[12\]\[24\] cpuregs\[13\]\[24\] net686 VGND VGND VPWR VPWR _05918_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11173_ cpuregs\[17\]\[22\] net633 net610 _05850_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__o211a_1
XFILLER_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_42_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09753__A decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10124_ _04846_ _04847_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__nor2_1
XFILLER_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10055_ _04802_ _04803_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__nor2_1
X_14932_ clknet_leaf_182_clk _01284_ VGND VGND VPWR VPWR cpuregs\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14863_ clknet_leaf_180_clk _01215_ VGND VGND VPWR VPWR cpuregs\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13814_ clknet_leaf_188_clk _00268_ VGND VGND VPWR VPWR cpuregs\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12257__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14794_ clknet_leaf_67_clk _01146_ VGND VGND VPWR VPWR decoded_imm\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13745_ clknet_leaf_17_clk _00199_ VGND VGND VPWR VPWR cpuregs\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10957_ cpuregs\[6\]\[17\] cpuregs\[7\]\[17\] net659 VGND VGND VPWR VPWR _05640_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09673__B2 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08308__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13676_ clknet_leaf_150_clk _00130_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_10888_ cpuregs\[12\]\[15\] cpuregs\[13\]\[15\] net647 VGND VGND VPWR VPWR _05573_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12338__B decoded_imm_j\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15415_ clknet_leaf_41_clk _01754_ VGND VGND VPWR VPWR cpuregs\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ net1194 genblk1.genblk1.pcpi_mul.next_rs2\[13\] net915 net238 VGND VGND VPWR
+ VPWR _02063_ sky130_fd_sc_hd__a22o_1
XANTENNA__08228__A2 net1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07436__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11232__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15346_ clknet_leaf_12_clk _01686_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12558_ net874 _02038_ _02039_ net389 VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__a31oi_1
XFILLER_157_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11509_ net193 net3048 net746 VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__mux2_1
X_15277_ clknet_leaf_191_clk _01618_ VGND VGND VPWR VPWR cpuregs\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold107 cpuregs\[22\]\[26\] VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ net2536 net871 VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__or2_1
Xhold118 cpuregs\[26\]\[23\] VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09139__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold129 cpuregs\[16\]\[8\] VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ clknet_leaf_175_clk _00682_ VGND VGND VPWR VPWR reg_next_pc\[5\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_60_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14159_ clknet_leaf_94_clk _00613_ VGND VGND VPWR VPWR count_instr\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_146_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout609 _03148_ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkbuf_4
X_06981_ net1119 _02556_ genblk2.pcpi_div.quotient\[9\] VGND VGND VPWR VPWR _02558_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08720_ net893 _04075_ _04077_ net2650 net1201 VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_124_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1180 net97 VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__buf_4
X_08651_ genblk1.genblk1.pcpi_mul.rd\[26\] genblk1.genblk1.pcpi_mul.next_rs2\[27\]
+ net1105 VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__nand3_1
Xfanout1191 net1205 VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__buf_2
XFILLER_94_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15173__Q mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10321__B net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07602_ _03117_ _03119_ _03124_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__or3_1
XANTENNA__12248__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08582_ _03959_ _03960_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09602__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07533_ _03058_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__nand2_1
XANTENNA__13124__S net438 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11433__A net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11471__A1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07675__B1 net811 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07464_ _02976_ _02983_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_157_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09203_ net1587 net539 net492 VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07395_ net8 net939 net936 VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12963__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08219__A2 net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13212__A2 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09134_ net1620 net578 net501 VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1067_A net1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09065_ net1386 net573 net511 VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1234_A net1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08016_ _03351_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09049__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold630 cpuregs\[3\]\[15\] VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold641 cpuregs\[28\]\[17\] VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold652 cpuregs\[4\]\[28\] VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12723__B2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold663 cpuregs\[4\]\[17\] VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 cpuregs\[27\]\[17\] VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 cpuregs\[4\]\[30\] VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1022_X net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold696 cpuregs\[4\]\[31\] VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09967_ _04448_ _04449_ net1129 VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout861_A net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08918_ _04156_ _04158_ _04155_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__a21bo_1
XFILLER_40_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09898_ _04664_ _04668_ _04662_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__a21oi_1
Xhold1330 reg_next_pc\[26\] VGND VGND VPWR VPWR net2644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 _00002_ VGND VGND VPWR VPWR net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 genblk2.pcpi_div.divisor\[46\] VGND VGND VPWR VPWR net2666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 genblk2.pcpi_div.divisor\[13\] VGND VGND VPWR VPWR net2677 sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ _04186_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__inv_2
XANTENNA__10231__B net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_X net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1374 is_sll_srl_sra VGND VGND VPWR VPWR net2688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 mem_rdata_q\[0\] VGND VGND VPWR VPWR net2699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 is_alu_reg_reg VGND VGND VPWR VPWR net2710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12239__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11860_ _06307_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08476__X _03873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ cpuregs\[2\]\[13\] cpuregs\[3\]\[13\] net660 VGND VGND VPWR VPWR _05498_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _06261_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout914_X net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12439__A net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13034__S net446 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11343__A net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13530_ net407 net1870 net416 VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__mux2_1
XANTENNA__07666__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10742_ net828 _05426_ _05428_ _05430_ net789 VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11462__B2 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10673_ cpuregs\[8\]\[9\] net667 VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__or2_1
X_13461_ net1583 net537 net424 VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__mux2_1
XFILLER_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_1270 VGND VGND VPWR VPWR picorv32_1270/HI eoi[28] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15200_ clknet_leaf_38_clk _01549_ VGND VGND VPWR VPWR cpuregs\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xpicorv32_1281 VGND VGND VPWR VPWR picorv32_1281/HI trace_data[3] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12412_ net323 net1738 net472 VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1292 VGND VGND VPWR VPWR picorv32_1292/HI trace_data[14] sky130_fd_sc_hd__conb_1
X_13392_ net1007 net756 VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__or2_1
X_15131_ clknet_leaf_0_clk _01483_ VGND VGND VPWR VPWR cpuregs\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ mem_rdata_q\[23\] _06223_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__and2_1
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12174__A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12274_ _06250_ _06614_ _06612_ _06239_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__a211o_1
X_15062_ clknet_leaf_105_clk net2108 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14013_ clknet_leaf_199_clk _00467_ VGND VGND VPWR VPWR cpuregs\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12714__B2 net1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11225_ cpuregs\[22\]\[24\] cpuregs\[23\]\[24\] net687 VGND VGND VPWR VPWR _05901_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11156_ cpuregs\[9\]\[22\] net633 net610 _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__o211a_1
XANTENNA_output244_A net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10107_ net2841 _04835_ net1225 VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10422__A net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11087_ net772 _05758_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__and3_1
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10038_ _04791_ _04792_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__nor2_1
X_14915_ clknet_leaf_125_clk _01267_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14846_ clknet_leaf_38_clk _01198_ VGND VGND VPWR VPWR cpuregs\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11494__D_N net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14777_ clknet_leaf_154_clk _00032_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_170_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11989_ _06335_ _06338_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12349__A mem_rdata_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13728_ clknet_leaf_122_clk _00182_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07657__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13659_ clknet_leaf_108_clk _00113_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_185_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07180_ net1065 net1045 _02728_ _02730_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__a211o_1
X_15329_ clknet_leaf_52_clk _01669_ VGND VGND VPWR VPWR cpuregs\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15168__Q mem_rdata_q\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10316__B net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout406 _03785_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12181__A2 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout417 _02357_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_4
X_09821_ _04592_ _04597_ _04590_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__o21ai_1
Xfanout428 net430 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_4
Xfanout439 net440 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__buf_4
XANTENNA_clkload12_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12531__B net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13119__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09752_ decoded_imm_j\[11\] _04432_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06964_ genblk2.pcpi_div.dividend\[7\] net1119 _02541_ net948 VGND VGND VPWR VPWR
+ _02543_ sky130_fd_sc_hd__a31o_1
XANTENNA__08137__A1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08703_ genblk1.genblk1.pcpi_mul.rd\[34\] genblk1.genblk1.pcpi_mul.next_rs2\[35\]
+ net1101 VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__nand3_1
X_06895_ is_jalr_addi_slti_sltiu_xori_ori_andi is_lui_auipc_jal net1088 VGND VGND
+ VPWR VPWR _02491_ sky130_fd_sc_hd__or3b_1
XANTENNA__12958__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09683_ net1187 _04425_ _04480_ _02489_ net848 VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__o221a_1
XFILLER_94_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11692__A1 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08634_ _04003_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09332__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11434__Y _06105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08565_ genblk1.genblk1.pcpi_mul.next_rs2\[14\] net1093 genblk1.genblk1.pcpi_mul.rd\[13\]
+ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__a21o_1
XANTENNA__13433__A2 net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09637__B2 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07516_ net358 _03039_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__o21bai_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12641__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08496_ _03886_ _03887_ _03882_ net761 VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__a211o_1
XFILLER_168_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07447_ reg_pc\[19\] decoded_imm\[19\] _02954_ _02978_ _02979_ VGND VGND VPWR VPWR
+ _02980_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_170_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_170_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_137_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout707_A _03139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07378_ count_instr\[47\] net1132 net1140 count_cycle\[47\] VGND VGND VPWR VPWR _02916_
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12706__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09117_ net2094 net310 net506 VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1237_X net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10955__B1 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09048_ net317 net2346 net513 VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__mux2_1
XFILLER_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold460 cpuregs\[2\]\[2\] VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12722__A _02404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold471 cpuregs\[30\]\[1\] VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold482 cpuregs\[27\]\[7\] VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net787 _05687_ _05689_ _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__or4_1
Xhold493 net153 VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12172__A2 net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10183__A1 net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout940 _02693_ VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13029__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout951 net952 VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout962 net965 VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10242__A decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout973 net974 VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout984 _02381_ VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__clkbuf_4
Xfanout995 net224 VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__buf_4
XFILLER_46_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12961_ net297 net2035 net454 VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_18_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1160 cpuregs\[18\]\[3\] VGND VGND VPWR VPWR net2474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11772__S net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14700_ clknet_leaf_152_clk _01085_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1171 cpuregs\[1\]\[3\] VGND VGND VPWR VPWR net2485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 cpuregs\[11\]\[25\] VGND VGND VPWR VPWR net2496 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _06369_ _06376_ _06379_ _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__o31a_1
XFILLER_85_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12880__A0 mem_rdata_q\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12892_ mem_rdata_q\[29\] net22 net964 VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__mux2_1
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1193 cpuregs\[11\]\[1\] VGND VGND VPWR VPWR net2507 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_47_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09242__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13272__B _05386_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ clknet_leaf_137_clk _01016_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10891__C1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11843_ genblk2.pcpi_div.divisor\[3\] genblk2.pcpi_div.dividend\[3\] VGND VGND VPWR
+ VPWR _06314_ sky130_fd_sc_hd__and2b_1
XFILLER_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14562_ clknet_leaf_41_clk _00948_ VGND VGND VPWR VPWR cpuregs\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11774_ net170 net133 net536 VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__mux2_1
X_13513_ net2013 net303 net421 VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__mux2_1
X_10725_ _05413_ _05414_ net814 VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__mux2_1
X_14493_ clknet_leaf_95_clk _00882_ VGND VGND VPWR VPWR instr_sll sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_161_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_161_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06862__A1 net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13444_ reg_pc\[29\] net566 _02345_ _02346_ net393 VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__a2111o_1
X_10656_ cpuregs\[19\]\[8\] net626 net594 VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__o21a_1
XANTENNA_output194_A net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__12108__S net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload27 clknet_leaf_180_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__inv_6
X_10587_ net1171 net855 _05279_ _05280_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__a22o_1
X_13375_ net710 _02263_ _02285_ net566 reg_pc\[21\] VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__a32o_1
XANTENNA__10417__A net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload38 clknet_leaf_192_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__clkinv_2
Xclkload49 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload49/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09800__B2 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15114_ clknet_leaf_39_clk _01466_ VGND VGND VPWR VPWR cpuregs\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12326_ decoded_imm\[11\] net745 _06641_ _06642_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__o22a_1
XFILLER_142_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15045_ clknet_leaf_112_clk net1579 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12257_ genblk2.pcpi_div.divisor\[20\] net377 net364 net2731 VGND VGND VPWR VPWR
+ _01126_ sky130_fd_sc_hd__a22o_1
XANTENNA_output71_A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13360__A1 net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07285__X _02829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11208_ cpuregs\[9\]\[23\] net623 net606 _05884_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_112_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12188_ net749 _06586_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nor2_1
X_11139_ net824 _05813_ _05815_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__a211o_1
XFILLER_110_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11123__B1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12871__A0 mem_rdata_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10477__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09152__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14829_ clknet_leaf_179_clk _01181_ VGND VGND VPWR VPWR cpuregs\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09619__B2 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08350_ reg_pc\[6\] _03764_ reg_pc\[7\] VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__a21oi_1
X_07301_ genblk1.genblk1.pcpi_mul.pcpi_rd\[10\] genblk2.pcpi_div.pcpi_rd\[10\] net1110
+ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__mux2_1
X_08281_ net1017 _03724_ net981 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_154_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_152_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_152_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_119_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13179__A1 _03799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07232_ _02774_ _02776_ _02778_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__nand3_1
XFILLER_20_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11729__A2 _06242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07163_ net1049 net1067 _02711_ net1082 _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07094_ net1122 _02651_ genblk2.pcpi_div.quotient\[25\] VGND VGND VPWR VPWR _02655_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_160_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13351__A1 net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09327__S net482 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13357__B net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A _04888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14530__Q decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09804_ decoded_imm_j\[15\] _04436_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__or2_1
XFILLER_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout269 net272 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_4
X_07996_ net968 _03317_ net934 _03315_ _03506_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_2_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ _04522_ _04525_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__or2_1
X_06947_ net1125 _02528_ net3058 VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11114__B1 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout657_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13373__A net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09666_ _04463_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__and2_1
X_06878_ _02474_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__nand2_1
XANTENNA__09062__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08617_ genblk1.genblk1.pcpi_mul.next_rs2\[22\] net1102 genblk1.genblk1.pcpi_mul.rd\[21\]
+ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__a21o_1
XFILLER_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout445_X net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09597_ reg_pc\[4\] net878 _04425_ net848 VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout824_A net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_X net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08548_ _03930_ _03931_ _03925_ _03928_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a211o_1
XFILLER_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout612_X net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ genblk1.genblk1.pcpi_mul.mul_waiting net1223 VGND VGND VPWR VPWR _03875_
+ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_143_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_143_clk sky130_fd_sc_hd__clkbuf_8
X_10510_ net987 decoded_imm\[3\] net856 VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__a21o_1
X_11490_ latched_branch _06150_ _06155_ _03740_ net1232 VGND VGND VPWR VPWR _00813_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_21_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08406__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10441_ cpuregs\[0\]\[0\] net555 _05140_ net785 VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__o22a_1
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13160_ net1375 net295 net433 VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__mux2_1
X_10372_ net999 net992 _02474_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__mux2_1
XFILLER_124_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout981_X net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12111_ net1001 _06549_ net724 VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__o21ai_1
X_13091_ net304 net1902 net442 VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__mux2_1
XFILLER_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12042_ genblk2.pcpi_div.dividend\[17\] _06495_ net269 VGND VGND VPWR VPWR _01026_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09237__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12145__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold290 cpuregs\[13\]\[23\] VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11068__A net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07572__A2 net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout770 net771 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout781 net782 VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout792 net795 VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12598__S net470 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13993_ clknet_leaf_49_clk _00447_ VGND VGND VPWR VPWR cpuregs\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12448__A3 net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15732_ net1173 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11656__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12944_ net408 net2185 net451 VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__mux2_1
X_12875_ mem_rdata_q\[12\] net4 net963 VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output207_A net1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14614_ clknet_leaf_114_clk _01000_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dfxtp_1
X_11826_ genblk2.pcpi_div.divisor\[12\] genblk2.pcpi_div.dividend\[12\] VGND VGND
+ VPWR VPWR _06297_ sky130_fd_sc_hd__nand2b_1
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12605__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15594_ clknet_leaf_29_clk _01930_ VGND VGND VPWR VPWR cpuregs\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08285__A0 net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14545_ clknet_leaf_73_clk _00931_ VGND VGND VPWR VPWR cpuregs\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11757_ net1644 net111 net730 VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_134_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_134_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_99_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ net813 _05395_ _05397_ net828 VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__o211a_1
XANTENNA__10631__A2 net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14476_ clknet_leaf_95_clk _00865_ VGND VGND VPWR VPWR instr_lh sky130_fd_sc_hd__dfxtp_1
X_11688_ net2193 net573 net374 VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__mux2_1
XANTENNA__12346__B _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13427_ reg_pc\[27\] _05079_ _06034_ is_lui_auipc_jal VGND VGND VPWR VPWR _02332_
+ sky130_fd_sc_hd__o2bb2a_1
Xclkload105 clknet_leaf_40_clk VGND VGND VPWR VPWR clkload105/Y sky130_fd_sc_hd__clkinv_8
X_10639_ cpuregs\[10\]\[8\] net666 VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__or2_1
Xclkload116 clknet_leaf_33_clk VGND VGND VPWR VPWR clkload116/Y sky130_fd_sc_hd__bufinv_16
Xclkload127 clknet_leaf_56_clk VGND VGND VPWR VPWR clkload127/X sky130_fd_sc_hd__clkbuf_8
XFILLER_155_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload138 clknet_leaf_71_clk VGND VGND VPWR VPWR clkload138/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload149 clknet_leaf_132_clk VGND VGND VPWR VPWR clkload149/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13358_ net1014 net755 VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_77_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12309_ net3056 net743 _06632_ _06633_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__o22a_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13289_ net1029 net752 VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__or2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09147__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13333__A1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09537__B1 net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15028_ clknet_leaf_137_clk net1336 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_110_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07850_ _03366_ _03367_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__and2_2
XANTENNA__08986__S net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06801_ net1012 VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__inv_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07781_ net1164 net1026 VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__nor2_1
Xinput3 mem_rdata[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_49_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09520_ count_instr\[39\] count_instr\[38\] count_instr\[37\] _04372_ VGND VGND VPWR
+ VPWR _04377_ sky130_fd_sc_hd__and4_1
XANTENNA__07903__B net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11647__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09451_ count_instr\[15\] _04330_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__and2_1
XFILLER_80_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08402_ reg_pc\[17\] reg_pc\[16\] _03805_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__and3_1
XFILLER_52_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09382_ net1811 net330 net399 VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09610__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08333_ reg_out\[4\] alu_out_q\[4\] net1154 VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_125_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10083__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08264_ reg_out\[9\] reg_next_pc\[9\] net921 VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__mux2_1
XFILLER_165_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08028__B1 net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07215_ _02760_ _02761_ _02762_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__nand3_1
XANTENNA__14525__Q decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08195_ net1145 _03682_ _03683_ _03447_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__o22a_1
XANTENNA__12971__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07146_ count_instr\[32\] net1130 net1140 count_cycle\[32\] VGND VGND VPWR VPWR _02699_
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07077_ genblk2.pcpi_div.dividend\[22\] genblk2.pcpi_div.dividend\[21\] _02631_ VGND
+ VGND VPWR VPWR _02640_ sky130_fd_sc_hd__or3_1
XFILLER_161_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09057__S net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout774_A _03170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1009 net216 VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout395_X net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout941_A _02693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07979_ _03308_ net934 VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_145_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11616__A mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09718_ decoded_imm_j\[8\] _04429_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__or2_1
XANTENNA__07813__B net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10990_ net822 _05668_ _05670_ _05672_ net787 VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__a2111o_1
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_98_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09649_ reg_pc\[30\] net880 _04451_ net850 VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout827_X net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ net2730 net902 _02079_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__a21o_1
XFILLER_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11611_ net2727 net562 _06184_ _06201_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__a22o_1
XFILLER_24_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12591_ net331 net1913 net467 VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_116_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_169_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13042__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14330_ clknet_leaf_173_clk _06717_ VGND VGND VPWR VPWR reg_out\[10\] sky130_fd_sc_hd__dfxtp_1
X_11542_ net29 net27 net28 _06167_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__and4b_1
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14435__Q net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13012__A0 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14261_ clknet_leaf_123_clk _00715_ VGND VGND VPWR VPWR count_cycle\[6\] sky130_fd_sc_hd__dfxtp_1
X_11473_ _06124_ _06125_ _06142_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__a21oi_4
XFILLER_109_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13212_ reg_pc\[1\] net565 _02139_ _02140_ net392 VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__a221o_1
X_10424_ _02439_ _02493_ _05126_ _05121_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_59_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14192_ clknet_leaf_94_clk _00646_ VGND VGND VPWR VPWR count_instr\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13143_ net1367 net404 net432 VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__mux2_1
XANTENNA__07242__A1 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10355_ _05059_ _05060_ net806 VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__mux2_1
XANTENNA__12182__A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12613__C net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13074_ net521 net1895 net439 VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__mux2_1
X_10286_ decoded_imm\[16\] net1018 _04991_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12025_ net721 _06480_ net1021 VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13217__S net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13976_ clknet_leaf_190_clk _00430_ VGND VGND VPWR VPWR cpuregs\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12927_ net279 net2404 net458 VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__mux2_1
XFILLER_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15646_ clknet_leaf_35_clk _01982_ VGND VGND VPWR VPWR cpuregs\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08394__X _03807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12858_ net293 net2492 net461 VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__mux2_1
XFILLER_61_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11809_ genblk2.pcpi_div.divisor\[18\] genblk2.pcpi_div.dividend\[18\] VGND VGND
+ VPWR VPWR _06280_ sky130_fd_sc_hd__nand2b_1
Xclkbuf_leaf_107_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_8
X_15577_ clknet_leaf_42_clk _01913_ VGND VGND VPWR VPWR cpuregs\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12789_ net1221 genblk1.genblk1.pcpi_mul.next_rs1\[57\] net2367 net906 net762 VGND
+ VGND VPWR VPWR _01428_ sky130_fd_sc_hd__a221o_1
X_14528_ clknet_leaf_28_clk _00917_ VGND VGND VPWR VPWR decoded_imm_j\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13003__A0 _03749_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07481__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14459_ clknet_leaf_64_clk _00848_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07000_ genblk2.pcpi_div.dividend\[12\] net1118 _02572_ net947 VGND VGND VPWR VPWR
+ _02574_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10368__A1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08951_ net2430 _04252_ net943 VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__mux2_1
XANTENNA__15176__Q mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07902_ net1177 net1046 VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__and2b_1
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08882_ net904 _04212_ _04214_ net2721 net1217 VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__a32o_1
Xhold1704 instr_bne VGND VGND VPWR VPWR net3018 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07473__X _03005_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1715 instr_rdinstr VGND VGND VPWR VPWR net3029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1726 count_instr\[19\] VGND VGND VPWR VPWR net3040 sky130_fd_sc_hd__dlygate4sd3_1
X_07833_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__and2_1
Xhold1737 count_instr\[50\] VGND VGND VPWR VPWR net3051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1748 count_cycle\[32\] VGND VGND VPWR VPWR net3062 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_162_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13127__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07633__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07764_ net1171 net1039 VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nor2_1
XFILLER_65_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09503_ count_instr\[32\] _04363_ count_instr\[33\] VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__a21o_1
XANTENNA__12293__A1 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12966__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07695_ cpuregs\[26\]\[3\] net677 VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__or2_1
XANTENNA__09694__C1 net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1097_A net1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09434_ count_instr\[9\] _04318_ net1225 VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10843__A2 net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09340__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09365_ net2262 net584 net401 VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout522_A net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09997__B1 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08316_ latched_rd\[2\] latched_rd\[4\] latched_rd\[3\] VGND VGND VPWR VPWR _03744_
+ sky130_fd_sc_hd__or3_1
XFILLER_166_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09296_ _04289_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__inv_2
XFILLER_20_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08247_ net258 net941 _03706_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__a21o_1
XANTENNA__07472__A1 genblk2.pcpi_div.pcpi_rd\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_X net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11005__C1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12348__A2 net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08480__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08178_ _03296_ _03663_ _03295_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10359__B2 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A net898 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07224__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_A net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09295__B _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07129_ genblk2.pcpi_div.dividend\[30\] _02678_ net1123 VGND VGND VPWR VPWR _02684_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07224__B2 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07808__B net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ count_cycle\[51\] count_cycle\[52\] _04854_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput170 net170 VGND VGND VPWR VPWR mem_wstrb[3] sky130_fd_sc_hd__buf_2
XANTENNA__10234__B net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput181 net181 VGND VGND VPWR VPWR pcpi_insn[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout777_X net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput192 net192 VGND VGND VPWR VPWR pcpi_insn[29] sky130_fd_sc_hd__buf_2
X_10071_ count_cycle\[26\] count_cycle\[27\] _04811_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__and3_1
XFILLER_121_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07824__A net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13037__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13830_ clknet_leaf_36_clk _00284_ VGND VGND VPWR VPWR cpuregs\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13761_ clknet_leaf_41_clk _00215_ VGND VGND VPWR VPWR cpuregs\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_10973_ net791 _05651_ _05653_ _05655_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__or4_1
X_15500_ clknet_leaf_133_clk _01836_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dfxtp_1
XFILLER_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12712_ net1192 genblk1.genblk1.pcpi_mul.next_rs1\[5\] net914 net231 VGND VGND VPWR
+ VPWR _02090_ sky130_fd_sc_hd__a22o_1
X_13692_ clknet_leaf_106_clk _00146_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09250__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13280__B _05421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15431_ clknet_leaf_18_clk _01770_ VGND VGND VPWR VPWR cpuregs\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_71_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12643_ net1202 genblk1.genblk1.pcpi_mul.next_rs2\[21\] net916 net247 VGND VGND VPWR
+ VPWR _02071_ sky130_fd_sc_hd__a22o_1
X_15362_ clknet_leaf_64_clk _01702_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09988__B1 net1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12574_ net585 net2350 net469 VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__mux2_1
XANTENNA__10409__B net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14313_ clknet_leaf_101_clk _00767_ VGND VGND VPWR VPWR count_cycle\[58\] sky130_fd_sc_hd__dfxtp_1
X_11525_ mem_rdata_q\[18\] net2611 net742 VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__mux2_1
XFILLER_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15293_ clknet_leaf_56_clk _01634_ VGND VGND VPWR VPWR cpuregs\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13500__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12339__A2 net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14244_ clknet_leaf_76_clk _00698_ VGND VGND VPWR VPWR reg_next_pc\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11456_ cpuregs\[20\]\[30\] cpuregs\[21\]\[30\] net688 VGND VGND VPWR VPWR _06126_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10407_ net1159 net247 _05111_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__or3_1
X_14175_ clknet_leaf_111_clk _00629_ VGND VGND VPWR VPWR count_instr\[46\] sky130_fd_sc_hd__dfxtp_1
X_11387_ cpuregs\[27\]\[28\] net637 net598 _06058_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__o211a_1
XFILLER_125_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11020__S net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13126_ net296 net2294 net437 VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__mux2_1
XFILLER_125_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10338_ cpuregs\[0\]\[31\] net694 VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__or2_1
XFILLER_124_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10770__A1 net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11955__S net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13057_ net2467 net80 net536 VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__mux2_1
X_10269_ _04935_ _04936_ _04973_ _04934_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__a31o_1
XFILLER_78_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12008_ net862 _06346_ _06463_ _06465_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__a32o_1
XANTENNA__09652__C decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08191__A2 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13959_ clknet_leaf_60_clk _00413_ VGND VGND VPWR VPWR cpuregs\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11690__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07480_ _02993_ _02997_ _03008_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_122_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12027__B2 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15629_ clknet_leaf_192_clk _01965_ VGND VGND VPWR VPWR cpuregs\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09150_ net2073 net327 net502 VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__mux2_1
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08101_ _03339_ _03589_ _03400_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__o21ai_1
X_09081_ net1598 net320 net508 VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__mux2_1
XFILLER_135_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08032_ _03364_ _03538_ net770 VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__o21ai_1
XFILLER_163_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11538__A0 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold801 cpuregs\[25\]\[9\] VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold812 cpuregs\[11\]\[14\] VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 cpuregs\[1\]\[20\] VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 cpuregs\[6\]\[10\] VGND VGND VPWR VPWR net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 cpuregs\[5\]\[13\] VGND VGND VPWR VPWR net2159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold856 reg_sh\[1\] VGND VGND VPWR VPWR net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold867 cpuregs\[5\]\[11\] VGND VGND VPWR VPWR net2181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 cpuregs\[17\]\[10\] VGND VGND VPWR VPWR net2192 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _04751_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold889 cpuregs\[19\]\[2\] VGND VGND VPWR VPWR net2203 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_164_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08934_ genblk1.genblk1.pcpi_mul.rd\[5\] genblk1.genblk1.pcpi_mul.rd\[37\] net955
+ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__mux2_1
XANTENNA__10622__X _05315_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08299__X net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1012_A net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1501 genblk1.genblk1.pcpi_mul.rd\[60\] VGND VGND VPWR VPWR net2815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09335__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1512 genblk1.genblk1.pcpi_mul.next_rs2\[44\] VGND VGND VPWR VPWR net2826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13365__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08865_ genblk1.genblk1.pcpi_mul.next_rs2\[60\] net1105 genblk1.genblk1.pcpi_mul.rd\[59\]
+ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a21o_1
Xhold1523 genblk1.genblk1.pcpi_mul.pcpi_rd\[6\] VGND VGND VPWR VPWR net2837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout472_A _06664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10513__A1 net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1534 count_cycle\[6\] VGND VGND VPWR VPWR net2848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 genblk2.pcpi_div.quotient_msk\[13\] VGND VGND VPWR VPWR net2859 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1556 genblk1.genblk1.pcpi_mul.rd\[49\] VGND VGND VPWR VPWR net2870 sky130_fd_sc_hd__dlygate4sd3_1
X_07816_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__inv_2
Xhold1567 genblk2.pcpi_div.quotient\[21\] VGND VGND VPWR VPWR net2881 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08796_ genblk1.genblk1.pcpi_mul.next_rs2\[49\] net1094 _04138_ _04140_ VGND VGND
+ VPWR VPWR _04142_ sky130_fd_sc_hd__and4_1
Xhold1578 count_instr\[28\] VGND VGND VPWR VPWR net2892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 genblk2.pcpi_div.divisor\[28\] VGND VGND VPWR VPWR net2903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11069__A2 _05748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07747_ _02478_ _03264_ _03265_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__or3_1
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout737_A net738 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout358_X net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07678_ net618 net796 VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__nor2_1
XANTENNA__09070__S net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12018__A1 net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09417_ count_instr\[4\] _04307_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__or2_1
XANTENNA__11613__B mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10029__B1 net1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ net1955 net333 net475 VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__mux2_1
XFILLER_166_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10229__B net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09279_ net1525 net336 net484 VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__mux2_1
XFILLER_166_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11310_ cpuregs\[30\]\[26\] cpuregs\[31\]\[26\] net703 VGND VGND VPWR VPWR _05984_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07819__A net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11529__A0 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12290_ decoded_imm\[28\] net739 VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__and2_1
XANTENNA__08414__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11241_ cpuregs\[14\]\[24\] cpuregs\[15\]\[24\] net686 VGND VGND VPWR VPWR _05917_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10245__A net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12741__A2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11172_ cpuregs\[16\]\[22\] net682 VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__or2_1
XFILLER_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10123_ net2824 _04845_ net1228 VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__o21ai_1
XFILLER_103_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09245__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input33_A mem_ready VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10054_ net2972 _04800_ net1235 VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__o21ai_1
X_14931_ clknet_leaf_180_clk _01283_ VGND VGND VPWR VPWR cpuregs\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10504__A1 net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09370__A1 net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14862_ clknet_leaf_19_clk _01214_ VGND VGND VPWR VPWR cpuregs\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_13813_ clknet_leaf_190_clk _00267_ VGND VGND VPWR VPWR cpuregs\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14793_ clknet_leaf_67_clk _01145_ VGND VGND VPWR VPWR decoded_imm\[29\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13744_ clknet_leaf_31_clk _00198_ VGND VGND VPWR VPWR cpuregs\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10956_ net1161 net855 _05638_ _05639_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07684__A1 net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13675_ clknet_leaf_150_clk _00129_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10887_ _05569_ _05571_ net782 VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__a21o_1
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15414_ clknet_leaf_9_clk _01753_ VGND VGND VPWR VPWR cpuregs\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ net2629 net887 _02062_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__a21o_1
XFILLER_157_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15345_ clknet_leaf_189_clk _01685_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
X_12557_ genblk2.pcpi_div.divisor\[59\] net874 VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__or2_1
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07288__X _02832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11508_ net2648 net2645 net747 VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__mux2_1
XANTENNA__10440__B1 net611 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15276_ clknet_leaf_185_clk _01617_ VGND VGND VPWR VPWR cpuregs\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08324__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12488_ _05104_ net718 net1164 VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__a21bo_1
Xhold108 cpuregs\[31\]\[13\] VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold119 cpuregs\[16\]\[14\] VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ clknet_leaf_132_clk _00681_ VGND VGND VPWR VPWR reg_next_pc\[4\] sky130_fd_sc_hd__dfxtp_1
X_11439_ cpuregs\[4\]\[30\] cpuregs\[5\]\[30\] net688 VGND VGND VPWR VPWR _06109_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09944__A net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14158_ clknet_leaf_94_clk _00612_ VGND VGND VPWR VPWR count_instr\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11940__B1 net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11685__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13109_ net403 net2121 net436 VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__mux2_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14089_ clknet_leaf_56_clk _00543_ VGND VGND VPWR VPWR cpuregs\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_06980_ net1119 genblk2.pcpi_div.quotient\[9\] _02556_ VGND VGND VPWR VPWR _02557_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09155__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09361__A1 _03870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1170 net126 VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__clkbuf_4
X_08650_ genblk1.genblk1.pcpi_mul.next_rs2\[27\] net1108 genblk1.genblk1.pcpi_mul.rd\[26\]
+ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_124_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07183__B decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1181 net97 VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__buf_4
Xfanout1192 net1198 VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__buf_2
XANTENNA__08994__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07601_ net1069 net992 _03123_ net1085 _03122_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__a221o_1
X_08581_ _03953_ _03956_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__nand2_1
XANTENNA__13445__B1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07532_ reg_pc\[26\] decoded_imm\[26\] VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__or2_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07463_ _02992_ _02993_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__nand2_1
X_09202_ net1536 net542 net493 VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07394_ _02924_ _02929_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__nand2_1
XANTENNA__07427__A1 genblk2.pcpi_div.pcpi_rd\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09133_ net1474 net581 net502 VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__mux2_1
XANTENNA__11223__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13140__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_A net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09064_ net1434 net577 net508 VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__mux2_1
XANTENNA__08234__S net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10982__A1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08015_ net988 _03521_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14533__Q decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold620 cpuregs\[31\]\[30\] VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 cpuregs\[2\]\[26\] VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1227_A net1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold642 cpuregs\[7\]\[25\] VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 cpuregs\[7\]\[4\] VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold664 cpuregs\[27\]\[13\] VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold675 cpuregs\[25\]\[28\] VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10734__A1 net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold686 cpuregs\[4\]\[14\] VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 cpuregs\[27\]\[26\] VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A net696 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09966_ _04738_ _04739_ net2639 net879 VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12280__A is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1015_X net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09065__S net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08917_ net1196 net2640 net888 _04235_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__a22o_1
X_09897_ net1127 _04443_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__xor2_1
XFILLER_112_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_96_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_8
Xhold1320 genblk2.pcpi_div.divisor\[60\] VGND VGND VPWR VPWR net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout475_X net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_A net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1331 mem_rdata_q\[1\] VGND VGND VPWR VPWR net2645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09352__A1 net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1342 genblk1.genblk1.pcpi_mul.pcpi_rd\[20\] VGND VGND VPWR VPWR net2656 sky130_fd_sc_hd__dlygate4sd3_1
X_08848_ genblk1.genblk1.pcpi_mul.next_rs2\[57\] net1103 _04182_ _04184_ VGND VGND
+ VPWR VPWR _04186_ sky130_fd_sc_hd__and4_1
Xhold1353 reg_next_pc\[17\] VGND VGND VPWR VPWR net2667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 _01118_ VGND VGND VPWR VPWR net2678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 reg_next_pc\[10\] VGND VGND VPWR VPWR net2689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1386 genblk1.genblk1.pcpi_mul.next_rs2\[2\] VGND VGND VPWR VPWR net2700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08779_ net885 _04125_ _04127_ net2871 net1194 VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__a32o_1
Xhold1397 genblk1.genblk1.pcpi_mul.rdx\[40\] VGND VGND VPWR VPWR net2711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout642_X net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ net797 _05494_ _05496_ net838 VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__a211o_1
XFILLER_14_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08409__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ genblk2.pcpi_div.dividend\[29\] genblk2.pcpi_div.divisor\[29\] VGND VGND
+ VPWR VPWR _06261_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_0_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12439__B _02507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10741_ cpuregs\[27\]\[11\] net625 net593 _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__o211a_1
XANTENNA__11462__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13460_ net1929 net544 net423 VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__mux2_1
X_10672_ net813 _05360_ _05362_ net828 VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__o211a_1
Xpicorv32_1260 VGND VGND VPWR VPWR picorv32_1260/HI eoi[18] sky130_fd_sc_hd__conb_1
Xpicorv32_1271 VGND VGND VPWR VPWR picorv32_1271/HI eoi[29] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12411_ net326 net1891 net474 VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__mux2_1
XFILLER_138_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_1282 VGND VGND VPWR VPWR picorv32_1282/HI trace_data[4] sky130_fd_sc_hd__conb_1
X_13391_ net1012 net756 _02299_ net710 VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__o211a_1
Xpicorv32_1293 VGND VGND VPWR VPWR picorv32_1293/HI trace_data[15] sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_20_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13050__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15130_ clknet_leaf_9_clk _01482_ VGND VGND VPWR VPWR cpuregs\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08091__A1 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12342_ decoded_imm\[4\] net745 _06650_ _06651_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__o22a_1
X_15061_ clknet_leaf_105_clk net2505 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_12273_ mem_do_rdata mem_do_rinst mem_state\[1\] mem_state\[0\] VGND VGND VPWR VPWR
+ _06614_ sky130_fd_sc_hd__or4b_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14012_ clknet_leaf_197_clk _00466_ VGND VGND VPWR VPWR cpuregs\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09764__A net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11224_ net835 _05895_ _05897_ _05899_ net794 VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__a2111o_1
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09591__A1 reg_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12190__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11155_ cpuregs\[8\]\[22\] net682 VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__or2_1
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10106_ count_cycle\[38\] count_cycle\[39\] count_cycle\[40\] _04831_ VGND VGND VPWR
+ VPWR _04836_ sky130_fd_sc_hd__and4_1
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11086_ net824 _05761_ _05763_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__a211o_1
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output237_A net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10037_ net2720 _04790_ net1224 VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__o21ai_1
X_14914_ clknet_leaf_124_clk _01266_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11150__A1 net840 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13427__B1 _06034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14845_ clknet_leaf_43_clk _01197_ VGND VGND VPWR VPWR cpuregs\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11557__A_N mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13225__S net757 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14776_ clknet_leaf_154_clk _00031_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11988_ net1032 net723 _06448_ net862 VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__a31o_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07223__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13727_ clknet_leaf_142_clk _00181_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10939_ cpuregs\[16\]\[16\] net655 VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__or2_1
XANTENNA__09498__X _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13658_ clknet_leaf_107_clk _00112_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ _02392_ net912 VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__nor2_1
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13589_ net1320 VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_11_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
X_15328_ clknet_leaf_50_clk _01668_ VGND VGND VPWR VPWR cpuregs\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08082__A1 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10964__A1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07290__C1 _02829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15259_ clknet_leaf_20_clk _01600_ VGND VGND VPWR VPWR cpuregs\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12705__A2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout407 net408 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_2
X_09820_ _04604_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__and2_1
Xfanout418 _02357_ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_4
Xfanout429 net430 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkbuf_8
X_09751_ net2689 net875 _04539_ _04542_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__a22o_1
XANTENNA__11428__B net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06963_ net1119 _02541_ genblk2.pcpi_div.dividend\[7\] VGND VGND VPWR VPWR _02542_
+ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_78_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_8
X_08702_ genblk1.genblk1.pcpi_mul.next_rs2\[35\] net1101 genblk1.genblk1.pcpi_mul.rd\[34\]
+ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__a21o_1
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09682_ _04425_ _04471_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__xnor2_1
X_06894_ _02445_ _02490_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__and2_1
XFILLER_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07345__B1 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08633_ _03997_ _04000_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__nand2_1
XFILLER_94_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13135__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ net885 _03943_ _03945_ net2574 net1192 VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__a32o_1
XANTENNA__09637__A2 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07133__S net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07648__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07515_ net1067 net1005 _03043_ net1082 _03042_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__a221o_1
XANTENNA__12974__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08495_ genblk1.genblk1.pcpi_mul.rd\[2\] genblk1.genblk1.pcpi_mul.next_rs2\[3\] net1098
+ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout435_A net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12641__B2 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07446_ reg_pc\[19\] decoded_imm\[19\] decoded_imm\[18\] reg_pc\[18\] VGND VGND VPWR
+ VPWR _02979_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_137_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07377_ net936 _02912_ net358 VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout602_A _03153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09116_ net1882 net312 net506 VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__mux2_1
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10955__A1 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09047_ net322 net2137 net513 VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__mux2_1
XFILLER_135_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12157__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09022__A0 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold450 cpuregs\[31\]\[16\] VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold461 cpuregs\[15\]\[2\] VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 cpuregs\[28\]\[30\] VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12722__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold483 cpuregs\[28\]\[19\] VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 cpuregs\[2\]\[16\] VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10523__A net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10183__A2 _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11380__A1 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout930 _03462_ VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 _02693_ VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09949_ _04446_ _04447_ net1129 VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__o21a_1
Xfanout952 net953 VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 net965 VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_69_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10242__B net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout974 net975 VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 _02381_ VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net997 VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__buf_4
X_12960_ net301 net2172 net454 VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__mux2_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1150 cpuregs\[11\]\[18\] VGND VGND VPWR VPWR net2464 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07336__B1 _02876_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11911_ _06376_ _06377_ _06380_ _06381_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__o31a_1
XANTENNA__07832__A net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1161 cpuregs\[18\]\[20\] VGND VGND VPWR VPWR net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 cpuregs\[11\]\[30\] VGND VGND VPWR VPWR net2486 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ mem_rdata_q\[28\] net21 net964 VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__mux2_1
XANTENNA__12880__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1183 cpuregs\[11\]\[0\] VGND VGND VPWR VPWR net2497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13409__B1 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1194 genblk1.genblk1.pcpi_mul.next_rs1\[60\] VGND VGND VPWR VPWR net2508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13045__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ clknet_leaf_137_clk _01015_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11842_ genblk2.pcpi_div.dividend\[4\] genblk2.pcpi_div.divisor\[4\] VGND VGND VPWR
+ VPWR _06313_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_64_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ clknet_leaf_1_clk _00947_ VGND VGND VPWR VPWR cpuregs\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11773_ _06245_ _06248_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__and2_1
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13512_ net1947 net305 net422 VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__mux2_1
X_10724_ cpuregs\[20\]\[10\] cpuregs\[21\]\[10\] net668 VGND VGND VPWR VPWR _05414_
+ sky130_fd_sc_hd__mux2_1
X_14492_ clknet_leaf_93_clk _00881_ VGND VGND VPWR VPWR instr_sub sky130_fd_sc_hd__dfxtp_1
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13443_ net996 net757 net558 _02321_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_24_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06862__A2 net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10655_ cpuregs\[17\]\[8\] net626 net607 _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__o211a_1
XFILLER_127_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload17 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload17/X sky130_fd_sc_hd__clkbuf_4
X_13374_ net1002 net760 VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__or2_1
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload28 clknet_leaf_181_clk VGND VGND VPWR VPWR clkload28/X sky130_fd_sc_hd__clkbuf_4
X_10586_ net1077 decoded_imm\[6\] net860 VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__o21a_1
X_15113_ clknet_leaf_49_clk _01465_ VGND VGND VPWR VPWR cpuregs\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xclkload39 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__inv_6
X_12325_ is_beq_bne_blt_bge_bltu_bgeu mem_rdata_q\[7\] decoded_imm_j\[11\] net1151
+ net734 VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__a221o_1
XANTENNA__12148__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15044_ clknet_leaf_112_clk _01396_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_12256_ net2818 net377 net364 genblk2.pcpi_div.divisor\[20\] VGND VGND VPWR VPWR
+ _01125_ sky130_fd_sc_hd__a22o_1
XFILLER_170_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11207_ cpuregs\[8\]\[23\] net662 VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_112_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12124__S net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12187_ net2909 net274 net2937 VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11138_ cpuregs\[18\]\[21\] net554 _05816_ net784 VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_118_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11069_ cpu_state\[3\] _05748_ net856 VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11123__A1 net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12320__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12871__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11264__A net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14828_ clknet_leaf_24_clk _01180_ VGND VGND VPWR VPWR cpuregs\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09619__A2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14759_ clknet_leaf_139_clk _00044_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_07300_ count_cycle\[10\] net972 net841 _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_127_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08280_ reg_out\[17\] reg_next_pc\[17\] net922 VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07231_ _02761_ _02777_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__and2_1
X_07162_ count_cycle\[1\] net972 net842 _02713_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__o211a_1
XANTENNA__15179__Q mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07093_ genblk2.pcpi_div.dividend\[25\] _02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_132_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12139__B1 net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09608__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07917__A net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14811__Q decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07636__B net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09803_ decoded_imm_j\[15\] _04436_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__nand2_1
XFILLER_115_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07995_ _03318_ net928 VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nand2_1
XANTENNA__12969__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09734_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06946_ genblk2.pcpi_div.dividend\[3\] genblk2.pcpi_div.dividend\[2\] genblk2.pcpi_div.dividend\[1\]
+ genblk2.pcpi_div.dividend\[0\] VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_2_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09343__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09665_ decoded_imm_j\[3\] _04424_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__or2_1
XANTENNA__13373__B net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A _03156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06877_ reg_sh\[1\] reg_sh\[0\] VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__nor2_1
X_08616_ net895 _03987_ _03989_ net2559 net1203 VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__a32o_1
XANTENNA__10873__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09596_ _03757_ reg_next_pc\[4\] net923 VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__mux2_2
X_08547_ genblk1.genblk1.pcpi_mul.rd\[10\] genblk1.genblk1.pcpi_mul.next_rs2\[11\]
+ net1092 VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout1082_X net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10625__B1 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08478_ genblk1.genblk1.pcpi_mul.mul_waiting net1237 VGND VGND VPWR VPWR _03874_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07429_ net358 _02958_ _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout605_X net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08046__A1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10440_ cpuregs\[1\]\[0\] net635 net611 VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__o21a_1
XANTENNA__08046__B2 net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10371_ net569 _05076_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__nor2_1
XFILLER_164_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12110_ _06372_ _06373_ _06548_ net869 VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__a31o_1
XFILLER_152_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07827__A net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13090_ net305 net2318 net441 VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__mux2_1
XFILLER_123_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12041_ _06494_ _06493_ _06491_ net861 VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__a2bb2o_1
Xhold280 cpuregs\[12\]\[31\] VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 cpuregs\[24\]\[30\] VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10253__A decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10561__C1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout760 _04884_ VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__buf_2
XANTENNA__07891__A_N net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout771 _03464_ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__clkbuf_4
Xfanout782 _03152_ VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__buf_2
X_13992_ clknet_leaf_71_clk _00446_ VGND VGND VPWR VPWR cpuregs\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_184_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout793 net795 VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__buf_2
XANTENNA__09253__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15731_ net1175 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_1
X_12943_ net521 net2202 net451 VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__mux2_1
XFILLER_19_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10864__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12874_ mem_rdata_q\[11\] net3 net963 VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14613_ clknet_leaf_104_clk _00999_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dfxtp_1
X_11825_ genblk2.pcpi_div.divisor\[13\] genblk2.pcpi_div.dividend\[13\] VGND VGND
+ VPWR VPWR _06296_ sky130_fd_sc_hd__nand2b_1
XANTENNA_output102_A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15593_ clknet_leaf_22_clk _01929_ VGND VGND VPWR VPWR cpuregs\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_199_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12605__B2 net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13503__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14544_ clknet_leaf_46_clk _00930_ VGND VGND VPWR VPWR cpuregs\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11756_ net1437 net110 net727 VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10707_ net800 _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__or2_1
X_14475_ clknet_leaf_96_clk _00864_ VGND VGND VPWR VPWR instr_lb sky130_fd_sc_hd__dfxtp_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11687_ net1853 net578 net374 VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13426_ _02463_ _02325_ _02326_ _02330_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__a31o_1
X_10638_ cpuregs\[9\]\[8\] net628 net608 _05329_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__o211a_1
XFILLER_128_944 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload106 clknet_leaf_41_clk VGND VGND VPWR VPWR clkload106/X sky130_fd_sc_hd__clkbuf_8
XFILLER_139_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload117 clknet_leaf_72_clk VGND VGND VPWR VPWR clkload117/X sky130_fd_sc_hd__clkbuf_4
Xclkload128 clknet_leaf_58_clk VGND VGND VPWR VPWR clkload128/Y sky130_fd_sc_hd__inv_12
XFILLER_143_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload139 clknet_leaf_78_clk VGND VGND VPWR VPWR clkload139/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_114_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10862__S net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13357_ _02411_ net755 VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nand2_1
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10569_ _05261_ _05262_ net800 VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12308_ net1146 decoded_imm_j\[19\] net970 mem_rdata_q\[19\] VGND VGND VPWR VPWR
+ _06633_ sky130_fd_sc_hd__a22o_1
X_13288_ net567 _05456_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__nor2_1
XANTENNA__08332__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10434__Y _05134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15027_ clknet_leaf_138_clk net1543 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12239_ genblk2.pcpi_div.divisor\[2\] net385 net371 net2898 VGND VGND VPWR VPWR _01108_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11344__A1 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11693__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06800_ net1016 VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__inv_2
X_07780_ net1164 net1026 VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nand2_1
Xinput4 mem_rdata[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
XANTENNA__15462__Q mem_wordsize\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09450_ _04330_ _04331_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__nor2_1
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08401_ reg_pc\[16\] _03805_ reg_pc\[17\] VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_135_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09381_ net2004 net333 net399 VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__mux2_1
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11722__A net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08332_ net577 net2474 net528 VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__mux2_1
XANTENNA__06816__A net1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08263_ net1033 _03715_ net980 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07214_ reg_pc\[5\] decoded_imm\[5\] VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__nand2_1
XANTENNA__08028__A1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08194_ _02399_ net997 net990 VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__a21o_1
X_07145_ net1051 net1066 _02697_ net1086 VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout300_A _03852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10772__S net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_144_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09338__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07647__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07076_ _02636_ _02637_ _02639_ net949 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_160_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10791__C1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12493__B1_N net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07539__B1 _03065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10801__A net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07978_ _03490_ _03491_ _03486_ VGND VGND VPWR VPWR alu_out\[4\] sky130_fd_sc_hd__a21o_1
XANTENNA__08478__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09073__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09717_ decoded_imm_j\[8\] _04429_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__and2_1
XANTENNA__11616__B mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06929_ _02509_ _02512_ _02513_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout934_A _03459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09648_ _03866_ reg_next_pc\[30\] net924 VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__mux2_1
XANTENNA__10846__B1 net811 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09801__S net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ count_instr\[60\] _04413_ net1209 VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_26_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ net2608 net563 _06183_ _06202_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__a22o_1
X_12590_ net335 net2031 net467 VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__mux2_1
XFILLER_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11541_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__inv_2
XANTENNA__11271__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08019__A1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14260_ clknet_leaf_129_clk _00714_ VGND VGND VPWR VPWR count_cycle\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11472_ net774 _06133_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__and3_1
XANTENNA__08019__B2 net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13211_ net958 _04953_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_162_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10423_ net1089 _05125_ _02503_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__o21ai_1
X_14191_ clknet_leaf_94_clk _00645_ VGND VGND VPWR VPWR count_instr\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09248__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13142_ net1588 net407 net431 VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__mux2_1
X_10354_ cpuregs\[22\]\[31\] cpuregs\[23\]\[31\] net693 VGND VGND VPWR VPWR _05060_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07242__A2 _02783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13073_ net526 net1716 net439 VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__mux2_1
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10285_ _04987_ _04989_ _04990_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__a21oi_1
X_12024_ net1025 net1023 _06470_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__or3_1
XFILLER_78_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12402__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout590 net592 VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__buf_2
XFILLER_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13975_ clknet_leaf_183_clk _00429_ VGND VGND VPWR VPWR cpuregs\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkload9_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12926_ net284 net2253 net458 VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__mux2_1
XFILLER_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07702__B1 _03148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ clknet_leaf_16_clk _01981_ VGND VGND VPWR VPWR cpuregs\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12857_ net298 net2252 net462 VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__mux2_1
X_11808_ genblk2.pcpi_div.dividend\[19\] genblk2.pcpi_div.divisor\[19\] VGND VGND
+ VPWR VPWR _06279_ sky130_fd_sc_hd__and2b_1
X_12788_ net1221 net2286 net2491 net906 net762 VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__a221o_1
X_15576_ clknet_leaf_9_clk _01912_ VGND VGND VPWR VPWR cpuregs\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08327__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11739_ net1735 net1175 net729 VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__mux2_1
X_14527_ clknet_leaf_28_clk _00916_ VGND VGND VPWR VPWR decoded_imm_j\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07466__C1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14458_ clknet_leaf_64_clk _00847_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dfxtp_1
XANTENNA__06923__X _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11688__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13409_ net710 _02289_ _02315_ net566 reg_pc\[25\] VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__a32o_1
X_14389_ clknet_leaf_84_clk _00810_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dfxtp_1
XFILLER_116_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09158__S net503 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14361__Q net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08950_ genblk1.genblk1.pcpi_mul.rd\[13\] genblk1.genblk1.pcpi_mul.rd\[45\] net954
+ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__mux2_1
XANTENNA__07186__B net1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08997__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07901_ net1176 _02402_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__nand2_1
XFILLER_97_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ _04213_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08194__B1 net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1705 decoded_imm\[2\] VGND VGND VPWR VPWR net3019 sky130_fd_sc_hd__dlygate4sd3_1
X_07832_ net1167 net1031 VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__nand2_1
Xhold1716 count_cycle\[35\] VGND VGND VPWR VPWR net3030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1727 count_cycle\[13\] VGND VGND VPWR VPWR net3041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1738 is_compare VGND VGND VPWR VPWR net3052 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1749 decoded_imm\[15\] VGND VGND VPWR VPWR net3063 sky130_fd_sc_hd__dlygate4sd3_1
X_07763_ _03280_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__inv_2
XFILLER_38_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09502_ count_instr\[32\] _04363_ _04365_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__o21a_1
XFILLER_65_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07694_ cpuregs\[25\]\[3\] net629 net609 _03213_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__o211a_1
XFILLER_92_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09433_ count_instr\[9\] _04318_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__and2_1
XANTENNA__12548__A net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout348_A _03799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13143__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09364_ net2150 net586 net401 VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__mux2_1
XANTENNA__13242__A1 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08237__S net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08315_ latched_branch latched_store net850 VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09997__A1 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07457__C1 _02988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ latched_rd\[2\] _03743_ _04280_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__or3_1
XANTENNA__12982__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08246_ net256 net941 _03705_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__a21o_1
XFILLER_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13379__A _02410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08177_ net966 _03290_ _03291_ net929 _03667_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__a221o_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12283__A net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08480__B net1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10359__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_X net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09068__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07128_ _02681_ _02682_ _02683_ net948 VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07224__A2 net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A net898 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10515__B net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07059_ genblk2.pcpi_div.quotient\[18\] genblk2.pcpi_div.quotient\[19\] _02610_ VGND
+ VGND VPWR VPWR _02625_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_37_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11308__A1 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput160 net160 VGND VGND VPWR VPWR mem_wdata[3] sky130_fd_sc_hd__buf_2
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06983__A1 net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput171 net171 VGND VGND VPWR VPWR pcpi_insn[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput182 net182 VGND VGND VPWR VPWR pcpi_insn[1] sky130_fd_sc_hd__buf_2
XFILLER_0_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput193 net193 VGND VGND VPWR VPWR pcpi_insn[2] sky130_fd_sc_hd__buf_2
X_10070_ _04813_ net1236 _04812_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout672_X net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07824__B net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10819__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13760_ clknet_leaf_8_clk _00214_ VGND VGND VPWR VPWR cpuregs\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10972_ cpuregs\[11\]\[17\] net621 net590 _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__o211a_1
XFILLER_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07840__A net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12711_ net1688 net884 _02089_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__a21o_1
X_13691_ clknet_leaf_106_clk _00145_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13053__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11362__A net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12642_ net2752 net895 _02070_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__a21o_1
X_15430_ clknet_leaf_29_clk _01769_ VGND VGND VPWR VPWR cpuregs\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15361_ clknet_leaf_62_clk _01701_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
X_12573_ net588 net1910 net470 VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__mux2_1
XFILLER_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11524_ mem_rdata_q\[17\] net2109 net742 VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__mux2_1
X_14312_ clknet_leaf_101_clk _00766_ VGND VGND VPWR VPWR count_cycle\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09767__A decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15292_ clknet_4_10_0_clk _01633_ VGND VGND VPWR VPWR cpuregs\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14243_ clknet_leaf_76_clk _00697_ VGND VGND VPWR VPWR reg_next_pc\[20\] sky130_fd_sc_hd__dfxtp_1
X_11455_ _06112_ _06115_ _03171_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__o21a_1
XFILLER_125_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12744__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10406_ net244 _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_74_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14174_ clknet_leaf_111_clk _00628_ VGND VGND VPWR VPWR count_instr\[45\] sky130_fd_sc_hd__dfxtp_1
X_11386_ cpuregs\[26\]\[28\] net690 VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__or2_1
XANTENNA__10755__C1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output267_A net267 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13125_ net299 net2500 net437 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__mux2_1
X_10337_ _05041_ _05042_ net818 VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__mux2_1
XFILLER_140_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13056_ net1596 net79 net533 VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__mux2_1
X_10268_ _04936_ _04973_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__nand2_1
X_12007_ net1027 net723 _06464_ net862 VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__a31oi_1
XFILLER_94_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10199_ decoded_imm\[24\] net1004 VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13472__A1 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13958_ clknet_leaf_30_clk _00412_ VGND VGND VPWR VPWR cpuregs\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12909_ net349 net1960 net455 VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__mux2_1
XANTENNA__12680__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13889_ clknet_leaf_41_clk _00343_ VGND VGND VPWR VPWR cpuregs\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ clknet_leaf_178_clk _01964_ VGND VGND VPWR VPWR cpuregs\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08057__S net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07439__C1 _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15559_ clknet_leaf_45_clk _01895_ VGND VGND VPWR VPWR cpuregs\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11786__A1 genblk2.pcpi_div.outsign VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08100_ net1159 net1013 net932 _03598_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__a31o_1
XANTENNA__09677__A decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09080_ net2103 net324 net510 VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__mux2_1
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07454__A2 net1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08031_ net1143 _03536_ _03537_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__a21o_1
XANTENNA__09396__B net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06813__B net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold802 cpuregs\[13\]\[7\] VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold813 cpuregs\[30\]\[16\] VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold824 cpuregs\[11\]\[13\] VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 cpuregs\[27\]\[19\] VGND VGND VPWR VPWR net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 cpuregs\[10\]\[4\] VGND VGND VPWR VPWR net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 cpuregs\[17\]\[15\] VGND VGND VPWR VPWR net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _04752_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__nand2_1
Xhold868 cpuregs\[18\]\[9\] VGND VGND VPWR VPWR net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 cpuregs\[27\]\[4\] VGND VGND VPWR VPWR net2193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09616__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08933_ net2635 _04243_ net944 VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__mux2_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_A _03852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13138__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08864_ genblk1.genblk1.pcpi_mul.rd\[59\] genblk1.genblk1.pcpi_mul.next_rs2\[60\]
+ net1108 VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__nand3_1
XANTENNA__12042__S net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1502 genblk2.pcpi_div.divisor\[22\] VGND VGND VPWR VPWR net2816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07644__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10351__A net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1513 _01350_ VGND VGND VPWR VPWR net2827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1524 genblk1.genblk1.pcpi_mul.rd\[17\] VGND VGND VPWR VPWR net2838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10513__A2 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1535 instr_lhu VGND VGND VPWR VPWR net2849 sky130_fd_sc_hd__dlygate4sd3_1
X_07815_ _03331_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__and2_1
Xhold1546 count_cycle\[43\] VGND VGND VPWR VPWR net2860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12977__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1557 genblk1.genblk1.pcpi_mul.rd\[45\] VGND VGND VPWR VPWR net2871 sky130_fd_sc_hd__dlygate4sd3_1
X_08795_ genblk1.genblk1.pcpi_mul.next_rs2\[49\] net1094 _04138_ _04140_ VGND VGND
+ VPWR VPWR _04141_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_142_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1568 genblk2.pcpi_div.quotient_msk\[26\] VGND VGND VPWR VPWR net2882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1579 genblk2.pcpi_div.quotient_msk\[18\] VGND VGND VPWR VPWR net2893 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_A _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11734__X _06244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07746_ net1066 reg_sh\[4\] _02473_ _02701_ decoded_imm_j\[4\] VGND VGND VPWR VPWR
+ _03265_ sky130_fd_sc_hd__a32o_1
XANTENNA__12266__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09351__S net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07677_ cpuregs\[2\]\[3\] cpuregs\[3\]\[3\] net675 VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__mux2_1
XANTENNA__12671__C1 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout632_A net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07142__A1 net1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09416_ _04307_ _04308_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__nor2_1
XFILLER_41_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13214__A_N net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09347_ net1784 net338 net476 VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__mux2_1
XFILLER_12_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout420_X net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1162_X net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_X net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09278_ net1454 net339 net484 VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__mux2_1
X_08229_ net1056 net1171 net240 net1055 VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__a22o_1
XFILLER_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07819__B net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11240_ _05913_ _05915_ net785 VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__a21o_1
XFILLER_153_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11171_ _05847_ _05848_ net804 VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__mux2_1
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07835__A net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10122_ count_cycle\[44\] count_cycle\[45\] count_cycle\[46\] _04841_ VGND VGND VPWR
+ VPWR _04846_ sky130_fd_sc_hd__and4_1
XFILLER_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08430__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13048__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10053_ count_cycle\[20\] count_cycle\[21\] _04798_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__and3_1
X_14930_ clknet_leaf_19_clk _01282_ VGND VGND VPWR VPWR cpuregs\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input26_A mem_rdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14861_ clknet_leaf_179_clk _01213_ VGND VGND VPWR VPWR cpuregs\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13812_ clknet_leaf_178_clk _00266_ VGND VGND VPWR VPWR cpuregs\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_14792_ clknet_leaf_86_clk _01144_ VGND VGND VPWR VPWR decoded_imm\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12257__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09261__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10955_ net1078 _05637_ net855 VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__a21oi_1
X_13743_ clknet_leaf_44_clk _00197_ VGND VGND VPWR VPWR cpuregs\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12188__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13674_ clknet_leaf_150_clk _00128_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_10886_ cpuregs\[1\]\[15\] net549 _05570_ net798 net822 VGND VGND VPWR VPWR _05571_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_14_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15413_ clknet_leaf_9_clk _01752_ VGND VGND VPWR VPWR cpuregs\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12625_ net1194 genblk1.genblk1.pcpi_mul.next_rs2\[12\] net915 net1165 VGND VGND
+ VPWR VPWR _02062_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11768__A1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13511__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07436__A2 net1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12556_ _05116_ net719 _02397_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__a21o_1
X_15344_ clknet_leaf_189_clk _01684_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11507_ net2554 mem_rdata_q\[0\] net746 VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__mux2_1
XFILLER_156_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15275_ clknet_leaf_185_clk _01616_ VGND VGND VPWR VPWR cpuregs\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12487_ net1164 net715 _05104_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__or3b_1
XFILLER_144_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold109 cpuregs\[26\]\[24\] VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ cpuregs\[6\]\[30\] cpuregs\[7\]\[30\] net692 VGND VGND VPWR VPWR _06108_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output94_A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14226_ clknet_leaf_132_clk _00680_ VGND VGND VPWR VPWR reg_next_pc\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11966__S net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14157_ clknet_leaf_100_clk _00611_ VGND VGND VPWR VPWR count_instr\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10870__S net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11369_ cpuregs\[1\]\[28\] net551 _06040_ net805 net832 VGND VGND VPWR VPWR _06041_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__06920__Y _02508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06947__A1 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12651__A _02396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11940__A1 net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13108_ net407 net2207 net435 VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__mux2_1
X_14088_ clknet_leaf_59_clk _00542_ VGND VGND VPWR VPWR cpuregs\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13039_ net1348 net92 net535 VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__mux2_1
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1160 net243 VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__clkbuf_4
Xfanout1171 net125 VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1182 net1187 VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__clkbuf_4
Xfanout1193 net1197 VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__buf_2
X_07600_ genblk1.genblk1.pcpi_mul.pcpi_rd\[30\] genblk2.pcpi_div.pcpi_rd\[30\] net1112
+ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__mux2_1
XFILLER_54_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08580_ _03957_ _03958_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nand2_1
XANTENNA__12248__A2 net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13445__B2 net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09171__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07531_ reg_pc\[26\] decoded_imm\[26\] VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__nand2_1
X_07462_ _02992_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__and2_1
XANTENNA__07675__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09201_ net1916 net573 net494 VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__mux2_1
XANTENNA__11208__B1 net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06883__B1 _02478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07393_ _02924_ _02929_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__or2_1
XFILLER_33_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09132_ net2225 net585 net502 VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__mux2_1
XFILLER_31_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14814__Q decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09063_ net1404 net581 net511 VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__mux2_1
XFILLER_108_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08014_ net1168 net1033 _03522_ net1143 VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__a211o_1
XANTENNA__12708__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold610 net201 VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_135_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold621 cpuregs\[31\]\[25\] VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 cpuregs\[12\]\[12\] VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 cpuregs\[8\]\[7\] VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 cpuregs\[27\]\[27\] VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold665 cpuregs\[6\]\[27\] VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__06938__A1 genblk2.pcpi_div.outsign VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold676 cpuregs\[4\]\[0\] VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09346__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold687 net47 VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold698 cpuregs\[23\]\[8\] VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net1185 _04449_ net849 VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout582_A _03753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12280__B is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08916_ _04134_ _04136_ _04133_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__a21bo_1
XFILLER_100_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09896_ net851 _04675_ _04676_ net881 net2565 VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__a32o_1
XFILLER_112_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1310 genblk1.genblk1.pcpi_mul.rd\[2\] VGND VGND VPWR VPWR net2624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1008_X net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1321 genblk1.genblk1.pcpi_mul.pcpi_rd\[4\] VGND VGND VPWR VPWR net2635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 genblk1.genblk1.pcpi_mul.rdx\[8\] VGND VGND VPWR VPWR net2646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 genblk2.pcpi_div.divisor\[15\] VGND VGND VPWR VPWR net2657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08847_ genblk1.genblk1.pcpi_mul.next_rs2\[57\] net1103 _04182_ _04184_ VGND VGND
+ VPWR VPWR _04185_ sky130_fd_sc_hd__a22o_1
Xhold1354 genblk1.genblk1.pcpi_mul.next_rs2\[8\] VGND VGND VPWR VPWR net2668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout847_A net852 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1365 genblk1.genblk1.pcpi_mul.rdx\[44\] VGND VGND VPWR VPWR net2679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13392__A net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1376 genblk2.pcpi_div.divisor\[52\] VGND VGND VPWR VPWR net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1387 count_cycle\[48\] VGND VGND VPWR VPWR net2701 sky130_fd_sc_hd__dlygate4sd3_1
X_08778_ _04126_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__inv_2
XANTENNA__12239__A2 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1398 genblk1.genblk1.pcpi_mul.rdx\[16\] VGND VGND VPWR VPWR net2712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09081__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07729_ cpuregs\[28\]\[4\] cpuregs\[29\]\[4\] net701 VGND VGND VPWR VPWR _03248_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__A1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_X net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ cpuregs\[26\]\[11\] net665 VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__or2_1
XFILLER_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07666__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10671_ net800 _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout802_X net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpicorv32_1250 VGND VGND VPWR VPWR picorv32_1250/HI eoi[8] sky130_fd_sc_hd__conb_1
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12410_ net330 net2218 net471 VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__mux2_1
XFILLER_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpicorv32_1261 VGND VGND VPWR VPWR picorv32_1261/HI eoi[19] sky130_fd_sc_hd__conb_1
Xpicorv32_1272 VGND VGND VPWR VPWR picorv32_1272/HI eoi[30] sky130_fd_sc_hd__conb_1
XFILLER_167_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13390_ net998 _04884_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__or2_1
Xpicorv32_1283 VGND VGND VPWR VPWR picorv32_1283/HI trace_data[5] sky130_fd_sc_hd__conb_1
XANTENNA__08425__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1294 VGND VGND VPWR VPWR picorv32_1294/HI trace_data[16] sky130_fd_sc_hd__conb_1
X_12341_ net1151 decoded_imm_j\[4\] _06617_ mem_rdata_q\[11\] net734 VGND VGND VPWR
+ VPWR _06651_ sky130_fd_sc_hd__a221o_1
XFILLER_127_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08091__A2 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15060_ clknet_leaf_104_clk _01412_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_12272_ net1234 net268 _06612_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__a21o_1
X_14011_ clknet_leaf_196_clk _00465_ VGND VGND VPWR VPWR cpuregs\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11223_ cpuregs\[27\]\[24\] net640 net601 _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__o211a_1
XFILLER_122_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09256__S net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11154_ net804 _05829_ _05831_ net831 VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__o211a_1
XFILLER_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11087__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10105_ _04835_ net1225 _04834_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__and3b_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11085_ cpuregs\[18\]\[20\] net552 _05764_ net782 VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__o22a_1
XANTENNA__12478__A2 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10422__C net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10036_ count_cycle\[13\] count_cycle\[14\] count_cycle\[15\] _04786_ VGND VGND VPWR
+ VPWR _04791_ sky130_fd_sc_hd__and4_2
X_14913_ clknet_leaf_124_clk _01265_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input29_X net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output132_A net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13506__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12410__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14844_ clknet_leaf_13_clk _01196_ VGND VGND VPWR VPWR cpuregs\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13427__B2 is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06909__A net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08303__A0 net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14775_ clknet_leaf_153_clk _00030_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11987_ net723 _06448_ net1031 VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13726_ clknet_leaf_141_clk _00180_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10938_ _05620_ _05621_ net798 VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07657__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13657_ clknet_leaf_107_clk _00111_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10869_ cpuregs\[20\]\[14\] cpuregs\[21\]\[14\] net664 VGND VGND VPWR VPWR _05555_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12608_ net2700 net894 _02053_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__a21o_1
XFILLER_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13588_ net1323 VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_1
X_15327_ clknet_leaf_57_clk _01667_ VGND VGND VPWR VPWR cpuregs\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12539_ net1158 _05113_ net719 VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__o21ai_1
XFILLER_144_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15258_ clknet_leaf_32_clk _01599_ VGND VGND VPWR VPWR cpuregs\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11696__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14209_ clknet_leaf_26_clk _00663_ VGND VGND VPWR VPWR reg_pc\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15189_ clknet_leaf_179_clk _01538_ VGND VGND VPWR VPWR cpuregs\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11374__C1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09166__S net499 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout408 net409 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_2
Xfanout419 net422 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13627__D net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06962_ genblk2.pcpi_div.dividend\[6\] _02538_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__or2_1
X_09750_ net1183 _04431_ _04541_ _02489_ net846 VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__o221a_1
XFILLER_67_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08701_ net894 _04059_ _04061_ net2918 net1202 VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__a32o_1
X_09681_ _04477_ _04478_ _02480_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__o21ai_1
X_06893_ instr_jal _02479_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__nor2_1
XFILLER_95_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08632_ _04001_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__nand2_1
XANTENNA__07922__B net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13418__A1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11429__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08563_ _03944_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__inv_2
XANTENNA__14809__Q decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07514_ genblk1.genblk1.pcpi_mul.pcpi_rd\[24\] genblk2.pcpi_div.pcpi_rd\[24\] net1112
+ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__mux2_1
X_08494_ genblk1.genblk1.pcpi_mul.next_rs2\[3\] net1098 genblk1.genblk1.pcpi_mul.rd\[2\]
+ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__a21o_1
XANTENNA__07648__A2 decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10101__B1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07445_ _02953_ _02965_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout330_A _03818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13151__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net430 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07376_ net936 _02913_ _02387_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__a21o_1
XFILLER_149_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09115_ net1653 net316 net506 VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__mux2_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12990__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09270__A1 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10955__A2 _05637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ net326 net2411 net515 VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__mux2_1
XFILLER_164_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout797_A net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold440 cpuregs\[24\]\[15\] VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10804__A net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1125_X net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold451 cpuregs\[2\]\[25\] VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09076__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold462 cpuregs\[15\]\[15\] VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 cpuregs\[15\]\[28\] VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold484 cpuregs\[28\]\[9\] VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 cpuregs\[26\]\[19\] VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout964_A net965 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout920 net921 VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__clkbuf_4
Xfanout931 _03462_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__buf_2
XANTENNA__10183__A3 _04883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09948_ net1129 _04448_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__xor2_1
Xfanout942 _02690_ VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__buf_4
Xfanout953 _02508_ VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__clkbuf_4
Xfanout964 net965 VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__clkbuf_4
Xfanout975 _02421_ VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 _02379_ VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__clkbuf_4
Xfanout997 net223 VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__buf_4
X_09879_ net1184 _04441_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__or2_1
Xhold1140 cpuregs\[19\]\[23\] VGND VGND VPWR VPWR net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 cpuregs\[9\]\[23\] VGND VGND VPWR VPWR net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 genblk1.genblk1.pcpi_mul.next_rs1\[59\] VGND VGND VPWR VPWR net2476 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _06371_ _06373_ _06370_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__a21o_1
XANTENNA__07832__B net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1173 reg_next_pc\[23\] VGND VGND VPWR VPWR net2487 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13409__A1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12890_ mem_rdata_q\[27\] net20 net964 VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__mux2_1
XFILLER_73_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1184 net54 VGND VGND VPWR VPWR net2498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1195 cpuregs\[11\]\[28\] VGND VGND VPWR VPWR net2509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10891__A1 net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11841_ genblk2.pcpi_div.divisor\[4\] genblk2.pcpi_div.dividend\[4\] VGND VGND VPWR
+ VPWR _06312_ sky130_fd_sc_hd__nand2b_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ clknet_leaf_0_clk _00946_ VGND VGND VPWR VPWR cpuregs\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11772_ net169 net132 net536 VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__mux2_1
X_10723_ cpuregs\[22\]\[10\] cpuregs\[23\]\[10\] net668 VGND VGND VPWR VPWR _05413_
+ sky130_fd_sc_hd__mux2_1
X_13511_ net1678 net308 net420 VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__mux2_1
X_14491_ clknet_leaf_93_clk _00880_ VGND VGND VPWR VPWR instr_add sky130_fd_sc_hd__dfxtp_1
XANTENNA__13061__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13442_ net710 _02322_ _02336_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__and3_1
X_10654_ cpuregs\[16\]\[8\] net668 VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__or2_1
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08155__S net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07279__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13373_ net1010 net756 VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__or2_1
XFILLER_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08064__A2 net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10585_ net1077 _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__nand2_1
Xclkload18 clknet_leaf_4_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload29 clknet_leaf_182_clk VGND VGND VPWR VPWR clkload29/X sky130_fd_sc_hd__clkbuf_4
X_15112_ clknet_leaf_49_clk _01464_ VGND VGND VPWR VPWR cpuregs\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_39_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12324_ is_sb_sh_sw _06223_ mem_rdata_q\[31\] VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__o21a_1
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09549__C1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13297__A _02404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12255_ net2769 net377 net364 net2818 VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__a22o_1
X_15043_ clknet_leaf_125_clk _01395_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12405__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07295__A net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11206_ net798 _05880_ _05882_ net825 VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__o211a_1
XFILLER_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12186_ net751 net2686 VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ cpuregs\[19\]\[21\] net622 net591 VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__o21a_1
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11068_ net1075 decoded_imm\[19\] VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__or2_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12320__B2 mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10019_ _04780_ net1223 _04779_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__and3b_1
XFILLER_110_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10867__D1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14827_ clknet_leaf_23_clk _01179_ VGND VGND VPWR VPWR cpuregs\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14758_ clknet_leaf_141_clk _00043_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13709_ clknet_leaf_124_clk _00163_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14689_ clknet_leaf_143_clk _01074_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07230_ reg_pc\[5\] decoded_imm\[5\] _02747_ _02748_ _02746_ VGND VGND VPWR VPWR
+ _02777_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14364__Q net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07161_ count_instr\[33\] net1130 net977 _02712_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__a211o_1
XFILLER_157_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09685__A decoded_imm_j\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07092_ genblk2.pcpi_div.dividend\[24\] _02647_ net1121 VGND VGND VPWR VPWR _02653_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_146_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13336__B1 net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09802_ net2642 net875 _04589_ net845 VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__a22o_1
XFILLER_140_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07994_ _03500_ _03505_ VGND VGND VPWR VPWR alu_out\[6\] sky130_fd_sc_hd__nand2_1
XANTENNA__09624__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06945_ net1125 genblk2.pcpi_div.quotient\[4\] _02525_ net953 VGND VGND VPWR VPWR
+ _02527_ sky130_fd_sc_hd__a31o_1
X_09733_ _04522_ _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout280_A _03873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13146__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09664_ decoded_imm_j\[3\] _04424_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__nand2_1
X_06876_ reg_sh\[4\] _02473_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__or2_2
XFILLER_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07144__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08615_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__inv_2
XANTENNA__12985__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09595_ reg_pc\[3\] net878 _04424_ net848 VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout545_A net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12075__B1 net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08546_ genblk1.genblk1.pcpi_mul.next_rs2\[11\] net1091 genblk1.genblk1.pcpi_mul.rd\[10\]
+ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__a21o_1
XANTENNA__15619__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08477_ net278 net2506 net530 VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__mux2_1
XFILLER_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout712_A _02083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1075_X net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07428_ net1065 net1014 _02962_ net1079 _02961_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout500_X net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07359_ _02811_ _02897_ net1060 VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__o21a_1
XFILLER_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10370_ _05057_ _05058_ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__a21oi_4
XFILLER_136_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11629__D_N mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13327__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09029_ net580 net2524 net514 VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__mux2_1
XFILLER_151_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11547__A_N net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07827__B net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11338__C1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ net1016 net721 _06492_ net861 VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__a31o_1
Xhold270 cpuregs\[28\]\[27\] VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07557__A1 net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold281 cpuregs\[14\]\[17\] VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__B net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout967_X net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold292 cpuregs\[29\]\[20\] VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout750 net751 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__buf_2
XANTENNA__07843__A net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout772 _03170_ VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__buf_4
X_13991_ clknet_leaf_71_clk _00445_ VGND VGND VPWR VPWR cpuregs\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xfanout783 net784 VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__clkbuf_4
Xfanout794 net795 VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13056__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15730_ net122 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
X_12942_ net526 net2261 net451 VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__mux2_1
XFILLER_74_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12873_ mem_rdata_q\[10\] net2 net964 VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__mux2_1
XFILLER_46_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ clknet_leaf_104_clk _00998_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ genblk2.pcpi_div.dividend\[13\] genblk2.pcpi_div.divisor\[13\] VGND VGND
+ VPWR VPWR _06295_ sky130_fd_sc_hd__and2b_1
XFILLER_33_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15592_ clknet_leaf_31_clk _01928_ VGND VGND VPWR VPWR cpuregs\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14543_ clknet_leaf_39_clk _00929_ VGND VGND VPWR VPWR cpuregs\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12196__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11755_ net1546 net109 net727 VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__mux2_1
X_10706_ cpuregs\[12\]\[10\] cpuregs\[13\]\[10\] net664 VGND VGND VPWR VPWR _05396_
+ sky130_fd_sc_hd__mux2_1
X_14474_ clknet_leaf_88_clk _00863_ VGND VGND VPWR VPWR instr_jalr sky130_fd_sc_hd__dfxtp_2
XFILLER_140_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11686_ net1696 net582 net375 VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__mux2_1
XFILLER_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13425_ net710 _02308_ _02328_ _02329_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__a31o_1
X_10637_ cpuregs\[8\]\[8\] net667 VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__or2_1
Xclkload107 clknet_leaf_42_clk VGND VGND VPWR VPWR clkload107/Y sky130_fd_sc_hd__bufinv_16
XFILLER_128_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload118 clknet_leaf_73_clk VGND VGND VPWR VPWR clkload118/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload129 clknet_leaf_59_clk VGND VGND VPWR VPWR clkload129/Y sky130_fd_sc_hd__inv_6
X_10568_ cpuregs\[30\]\[6\] cpuregs\[31\]\[6\] net670 VGND VGND VPWR VPWR _05262_
+ sky130_fd_sc_hd__mux2_1
X_13356_ net569 _05748_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_114_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13318__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12307_ mem_rdata_q\[31\] _06618_ net733 VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__a21o_2
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13287_ net960 _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__nor2_1
X_10499_ cpuregs\[16\]\[1\] net688 VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__or2_1
X_15026_ clknet_leaf_139_clk _01378_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_12238_ genblk2.pcpi_div.divisor\[1\] net385 net371 net2964 VGND VGND VPWR VPWR _01107_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11259__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11974__S net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12169_ genblk2.pcpi_div.quotient_msk\[28\] net380 net368 net2732 VGND VGND VPWR
+ VPWR _01070_ sky130_fd_sc_hd__a22o_1
Xinput5 mem_rdata[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08400_ reg_out\[17\] alu_out_q\[17\] net1154 VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__mux2_1
X_09380_ net1886 net337 net399 VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__mux2_1
XFILLER_101_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08331_ _03754_ _03755_ net767 VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__mux2_2
XANTENNA__06816__B instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08262_ reg_out\[8\] reg_next_pc\[8\] net921 VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__mux2_1
XFILLER_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07213_ reg_pc\[5\] decoded_imm\[5\] VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__or2_1
X_08193_ _03266_ _03675_ _03267_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07144_ genblk1.genblk1.pcpi_mul.pcpi_rd\[0\] genblk2.pcpi_div.pcpi_rd\[0\] net1112
+ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__mux2_1
XANTENNA__07236__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06832__A _02379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07075_ genblk2.pcpi_div.quotient\[22\] _02638_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1035_A net1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07539__A1 net1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout495_A _04286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07539__B2 net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10543__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09354__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout662_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07977_ _03306_ _03489_ net770 VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__o21a_1
XANTENNA__08478__B net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09716_ net2560 net876 _04510_ net852 VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__a22o_1
X_06928_ genblk2.pcpi_div.dividend\[0\] net1126 genblk2.pcpi_div.dividend\[1\] VGND
+ VGND VPWR VPWR _02513_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout450_X net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09647_ reg_pc\[29\] net880 _04450_ net850 VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__a22o_1
XFILLER_28_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06859_ net1060 cpu_state\[6\] VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout548_X net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07711__A1 decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09578_ _04413_ _04414_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__nor2_1
XFILLER_24_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08529_ _03909_ _03912_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__nand2_1
XANTENNA__13260__A2 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11540_ _06165_ net26 net23 VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__or3b_1
XFILLER_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ net832 _06136_ _06138_ _06140_ net793 VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__a2111o_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10422_ net1081 net1088 net1068 VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__or3_2
X_13210_ net1051 decoded_imm\[0\] _04951_ _04952_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__a22o_1
X_14190_ clknet_leaf_94_clk _00644_ VGND VGND VPWR VPWR count_instr\[61\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10353_ cpuregs\[20\]\[31\] cpuregs\[21\]\[31\] net693 VGND VGND VPWR VPWR _05059_
+ sky130_fd_sc_hd__mux2_1
X_13141_ net1472 net520 net431 VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__mux2_1
XFILLER_151_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13072_ net537 net1770 net439 VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__mux2_1
X_10284_ decoded_imm\[16\] net1018 VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12023_ _06349_ _06350_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10534__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09264__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10711__B net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout580 _03753_ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__buf_1
XANTENNA__07292__B decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout591 net592 VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkbuf_4
X_13974_ clknet_leaf_190_clk _00428_ VGND VGND VPWR VPWR cpuregs\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input11_X net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12925_ net285 net2314 net457 VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__mux2_1
XANTENNA__10837__B2 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output212_A net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13514__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12039__B1 net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15644_ clknet_leaf_45_clk _01980_ VGND VGND VPWR VPWR cpuregs\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12856_ net302 net2287 net462 VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__mux2_1
XANTENNA__11542__B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11807_ genblk2.pcpi_div.divisor\[20\] genblk2.pcpi_div.dividend\[20\] VGND VGND
+ VPWR VPWR _06278_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15575_ clknet_leaf_9_clk _01911_ VGND VGND VPWR VPWR cpuregs\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12787_ net1219 net2236 net2286 net907 net763 VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__a221o_1
XFILLER_15_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13251__A2 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11034__S net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14526_ clknet_leaf_28_clk _00915_ VGND VGND VPWR VPWR decoded_imm_j\[16\] sky130_fd_sc_hd__dfxtp_1
X_11738_ net1876 net122 net727 VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__mux2_1
X_14457_ clknet_leaf_90_clk _00846_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dfxtp_1
X_11669_ net26 net23 _06165_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__or3_2
XANTENNA__07748__A net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ net994 net760 VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__or2_1
XANTENNA__08343__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14388_ clknet_leaf_85_clk _00809_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dfxtp_4
X_13339_ net1018 net752 net556 _02233_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__o211a_1
XFILLER_115_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10174__A net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09963__A net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07900_ net1172 net1041 VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__and2b_1
X_15009_ clknet_leaf_115_clk _01361_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_166_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ _04205_ _04208_ _04210_ _04211_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__o211a_1
XFILLER_96_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09174__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1706 genblk2.pcpi_div.dividend\[13\] VGND VGND VPWR VPWR net3020 sky130_fd_sc_hd__dlygate4sd3_1
X_07831_ net1167 net1031 VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__or2_1
XFILLER_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1717 genblk2.pcpi_div.pcpi_wait VGND VGND VPWR VPWR net3031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1728 count_instr\[15\] VGND VGND VPWR VPWR net3042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1739 count_instr\[6\] VGND VGND VPWR VPWR net3053 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07762_ net1171 net1039 VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__nand2_1
X_09501_ count_instr\[32\] _04363_ net1207 VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__a21oi_1
X_07693_ cpuregs\[24\]\[3\] net677 VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__or2_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07154__C1 net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09432_ _04318_ _04319_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_140_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14817__Q decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09363_ latched_rd\[1\] latched_rd\[0\] _04290_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__and3b_4
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08314_ latched_rd\[2\] latched_rd\[3\] latched_rd\[4\] VGND VGND VPWR VPWR _03742_
+ sky130_fd_sc_hd__or3b_1
XANTENNA__11253__A1 _02396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09294_ net2077 net278 net486 VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__mux2_1
XFILLER_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08245_ net255 net941 _03704_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__a21o_1
XFILLER_166_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1152_A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout508_A _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09349__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11005__A1 net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08176_ _03289_ net935 VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_183_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08253__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13379__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08480__C net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07127_ genblk2.pcpi_div.dividend\[30\] _02679_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10764__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1038_X net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07058_ genblk2.pcpi_div.dividend\[20\] net1117 _02622_ net947 VGND VGND VPWR VPWR
+ _02624_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_37_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput150 net150 VGND VGND VPWR VPWR mem_wdata[23] sky130_fd_sc_hd__buf_2
XFILLER_161_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput161 net161 VGND VGND VPWR VPWR mem_wdata[4] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A net882 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput172 net172 VGND VGND VPWR VPWR pcpi_insn[10] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_198_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput183 net183 VGND VGND VPWR VPWR pcpi_insn[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput194 net194 VGND VGND VPWR VPWR pcpi_insn[30] sky130_fd_sc_hd__buf_2
XFILLER_0_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10516__B1 net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1205_X net1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input3_X net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09084__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10971_ cpuregs\[10\]\[17\] net655 VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__or2_1
XANTENNA__10958__S net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_X net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12710_ net1198 net1339 net914 net1041 VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__a22o_1
XANTENNA__07696__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13690_ clknet_leaf_106_clk _00144_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07160__A2 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12641_ net1202 genblk1.genblk1.pcpi_mul.next_rs2\[20\] net916 net245 VGND VGND VPWR
+ VPWR _02070_ sky130_fd_sc_hd__a22o_1
XFILLER_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11244__A1 net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15360_ clknet_leaf_64_clk _01700_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12572_ _04275_ _06663_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__or2_2
XANTENNA__07999__A1 net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09400__X _04298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14311_ clknet_leaf_101_clk _00765_ VGND VGND VPWR VPWR count_cycle\[56\] sky130_fd_sc_hd__dfxtp_1
X_11523_ mem_rdata_q\[16\] net1973 net742 VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__mux2_1
XFILLER_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15291_ clknet_leaf_60_clk _01632_ VGND VGND VPWR VPWR cpuregs\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09259__S net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14242_ clknet_leaf_27_clk _00696_ VGND VGND VPWR VPWR reg_next_pc\[19\] sky130_fd_sc_hd__dfxtp_1
X_11454_ net793 _06119_ _06121_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__or4_2
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12744__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10405_ net1160 net1161 _05108_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__or3_1
XANTENNA__12744__B2 net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11385_ cpuregs\[25\]\[28\] net637 net612 _06056_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_74_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14173_ clknet_leaf_111_clk _00627_ VGND VGND VPWR VPWR count_instr\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13124_ net304 net2496 net438 VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_113_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10336_ cpuregs\[4\]\[31\] cpuregs\[5\]\[31\] net695 VGND VGND VPWR VPWR _05042_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13509__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_13055_ net2001 net78 net533 VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__mux2_1
XANTENNA__10281__X _04987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10267_ _04938_ _04964_ _04967_ _04970_ _04972_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__a41o_1
XANTENNA__12413__S net474 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_940 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12006_ net723 _06464_ net1026 VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__a21o_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10198_ decoded_imm\[25\] net1002 VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07923__A1 _02396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10868__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13957_ clknet_leaf_30_clk _00411_ VGND VGND VPWR VPWR cpuregs\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12649__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11553__A net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12908_ net352 net2006 net455 VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__mux2_1
XANTENNA__10286__A2 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13888_ clknet_leaf_2_clk _00342_ VGND VGND VPWR VPWR cpuregs\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08338__S net531 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15627_ clknet_leaf_21_clk _01963_ VGND VGND VPWR VPWR cpuregs\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12839_ net520 net2110 net460 VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09958__A net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15558_ clknet_leaf_39_clk _01894_ VGND VGND VPWR VPWR cpuregs\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08100__A1 net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11786__A2 _05120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11699__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14509_ clknet_leaf_80_clk _00898_ VGND VGND VPWR VPWR decoded_imm_j\[5\] sky130_fd_sc_hd__dfxtp_1
X_15489_ clknet_leaf_56_clk _01825_ VGND VGND VPWR VPWR cpuregs\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10994__B1 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08030_ _03358_ _03529_ net988 _03357_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__o211a_1
XANTENNA__09169__S net499 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput30 mem_rdata[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14372__Q net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12735__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold803 cpuregs\[7\]\[9\] VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 cpuregs\[6\]\[30\] VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 cpuregs\[7\]\[15\] VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold836 cpuregs\[25\]\[0\] VGND VGND VPWR VPWR net2150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09693__A net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold847 cpuregs\[10\]\[0\] VGND VGND VPWR VPWR net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 cpuregs\[3\]\[25\] VGND VGND VPWR VPWR net2172 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ net1129 _04451_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__or2_1
Xhold869 cpuregs\[11\]\[4\] VGND VGND VPWR VPWR net2183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08932_ genblk1.genblk1.pcpi_mul.rd\[4\] genblk1.genblk1.pcpi_mul.rd\[36\] net955
+ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_103_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1503 net134 VGND VGND VPWR VPWR net2817 sky130_fd_sc_hd__dlygate4sd3_1
X_08863_ net902 _04196_ _04198_ net2707 net1213 VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__a32o_1
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1514 genblk2.pcpi_div.quotient_msk\[22\] VGND VGND VPWR VPWR net2828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 genblk2.pcpi_div.quotient_msk\[19\] VGND VGND VPWR VPWR net2839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1536 pcpi_timeout_counter\[0\] VGND VGND VPWR VPWR net2850 sky130_fd_sc_hd__dlygate4sd3_1
X_07814_ net248 net1009 VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__nand2_1
Xhold1547 pcpi_timeout_counter\[1\] VGND VGND VPWR VPWR net2861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13448__C1 _02501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08794_ genblk1.genblk1.pcpi_mul.rd\[48\] genblk1.genblk1.pcpi_mul.rdx\[48\] VGND
+ VGND VPWR VPWR _04140_ sky130_fd_sc_hd__or2_1
Xhold1558 genblk1.genblk1.pcpi_mul.rd\[3\] VGND VGND VPWR VPWR net2872 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1569 genblk1.genblk1.pcpi_mul.rd\[7\] VGND VGND VPWR VPWR net2883 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09632__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07745_ net987 _03263_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout360_A net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09667__A1 decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13154__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07676_ net801 _03193_ _03195_ net838 VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__a211o_1
XFILLER_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07142__A2 _02384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09415_ net2982 _04305_ net1231 VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12993__S net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout625_A net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09346_ net1580 net340 net475 VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__mux2_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout413_X net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09277_ net1577 net343 net485 VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1155_X net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09079__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08228_ net1056 net1173 net239 net942 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__a22o_1
XFILLER_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout994_A net995 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08159_ net966 _03269_ _03270_ net935 VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__o2bb2a_1
X_11170_ cpuregs\[22\]\[22\] cpuregs\[23\]\[22\] net682 VGND VGND VPWR VPWR _05848_
+ sky130_fd_sc_hd__mux2_1
XFILLER_161_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout782_X net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10121_ _04845_ net1228 _04844_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__and3b_1
XANTENNA__07835__B net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10052_ _04800_ _04801_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14860_ clknet_leaf_23_clk _01212_ VGND VGND VPWR VPWR cpuregs\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07851__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13811_ clknet_leaf_24_clk _00265_ VGND VGND VPWR VPWR cpuregs\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_input19_A mem_rdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14791_ clknet_leaf_67_clk _01143_ VGND VGND VPWR VPWR decoded_imm\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09658__A1 decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12469__A net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13064__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11373__A net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13742_ clknet_leaf_36_clk _00196_ VGND VGND VPWR VPWR cpuregs\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_10954_ net1075 decoded_imm\[16\] VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13673_ clknet_leaf_149_clk _00127_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[43\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_191_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_191_clk sky130_fd_sc_hd__clkbuf_8
X_10885_ cpuregs\[2\]\[15\] cpuregs\[3\]\[15\] net656 VGND VGND VPWR VPWR _05570_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15412_ clknet_leaf_10_clk _01751_ VGND VGND VPWR VPWR cpuregs\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12624_ net1194 net2629 net887 net3004 _02061_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_100_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15343_ clknet_leaf_189_clk _01683_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
X_12555_ net254 net716 _05116_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__or3b_1
XANTENNA__12408__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11506_ _02380_ decoder_pseudo_trigger VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__or2_1
X_15274_ clknet_leaf_185_clk _01615_ VGND VGND VPWR VPWR cpuregs\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10440__A2 net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12486_ _06709_ _06710_ net2687 net386 VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_156_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12717__B2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14225_ clknet_leaf_132_clk _00679_ VGND VGND VPWR VPWR reg_next_pc\[2\] sky130_fd_sc_hd__dfxtp_1
X_11437_ net256 net857 _06106_ _06107_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__a22o_1
XANTENNA__10728__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07585__X _03109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output87_A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14156_ clknet_leaf_100_clk _00610_ VGND VGND VPWR VPWR count_instr\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11368_ cpuregs\[2\]\[28\] cpuregs\[3\]\[28\] net691 VGND VGND VPWR VPWR _06040_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12651__B net913 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11548__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13107_ net521 net2408 net435 VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__mux2_1
XANTENNA__11940__A2 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07745__B _03263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10319_ _04904_ _05024_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__nor2_1
X_14087_ clknet_leaf_60_clk _00541_ VGND VGND VPWR VPWR cpuregs\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11299_ cpuregs\[12\]\[26\] cpuregs\[13\]\[26\] net703 VGND VGND VPWR VPWR _05973_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_163_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ net1464 net91 net535 VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__mux2_1
XFILLER_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1150 net1152 VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__buf_2
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1161 net242 VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__clkbuf_4
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1172 net1173 VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1183 net1187 VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1197 VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__buf_2
XFILLER_94_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07761__A net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14989_ clknet_leaf_119_clk _01341_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09649__B2 net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07530_ net1073 _03049_ _03050_ _03057_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__a31o_1
XANTENNA__12653__B1 net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14367__Q net266 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07461_ reg_pc\[21\] decoded_imm\[21\] VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_182_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_182_clk sky130_fd_sc_hd__clkbuf_8
X_09200_ net1609 net577 net493 VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__mux2_1
XANTENNA__06883__A1 net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12405__A0 _03799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07392_ _02906_ _02925_ _02927_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_33_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07700__S net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09131_ net2071 net586 net502 VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__mux2_1
XANTENNA__08085__B1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09062_ net1950 net583 net510 VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__mux2_1
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12708__A1 net1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08013_ _03315_ _03508_ _03355_ _03317_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_135_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold600 cpuregs\[6\]\[11\] VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__B1 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold611 cpuregs\[27\]\[24\] VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 cpuregs\[13\]\[29\] VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13381__A1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold633 cpuregs\[15\]\[24\] VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold644 cpuregs\[22\]\[7\] VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 cpuregs\[8\]\[23\] VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 cpuregs\[15\]\[18\] VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 cpuregs\[27\]\[16\] VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13149__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold688 cpuregs\[22\]\[30\] VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 cpuregs\[15\]\[25\] VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ net985 _04734_ _04737_ net1185 VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__o211a_1
XANTENNA__07655__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08915_ net1194 net2679 net886 _04234_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__a22o_1
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10081__B net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12988__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09895_ net1184 _04442_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__or2_1
Xhold1300 genblk1.genblk1.pcpi_mul.rd\[1\] VGND VGND VPWR VPWR net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 genblk1.genblk1.pcpi_mul.rdx\[28\] VGND VGND VPWR VPWR net2625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 net197 VGND VGND VPWR VPWR net2636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12892__A0 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08846_ genblk1.genblk1.pcpi_mul.rd\[56\] genblk1.genblk1.pcpi_mul.rdx\[56\] VGND
+ VGND VPWR VPWR _04184_ sky130_fd_sc_hd__or2_1
Xhold1333 net143 VGND VGND VPWR VPWR net2647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06839__X _02443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1344 is_jalr_addi_slti_sltiu_xori_ori_andi VGND VGND VPWR VPWR net2658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09362__S net478 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1355 genblk2.pcpi_div.divisor\[43\] VGND VGND VPWR VPWR net2669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 net188 VGND VGND VPWR VPWR net2680 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13392__B net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1377 genblk1.genblk1.pcpi_mul.rd\[38\] VGND VGND VPWR VPWR net2691 sky130_fd_sc_hd__dlygate4sd3_1
X_08777_ _04117_ _04120_ _04122_ _04124_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__o211a_1
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout363_X net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13436__A2 _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1388 genblk2.pcpi_div.divisor\[17\] VGND VGND VPWR VPWR net2702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1399 genblk2.pcpi_div.quotient\[11\] VGND VGND VPWR VPWR net2713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07728_ cpuregs\[30\]\[4\] cpuregs\[31\]\[4\] net678 VGND VGND VPWR VPWR _03247_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout530_X net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_173_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_173_clk sky130_fd_sc_hd__clkbuf_8
X_07659_ net837 _03175_ _03177_ _03179_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__a211o_1
XFILLER_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout628_X net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10670_ cpuregs\[12\]\[9\] cpuregs\[13\]\[9\] net667 VGND VGND VPWR VPWR _05361_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07610__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1251 VGND VGND VPWR VPWR picorv32_1251/HI eoi[9] sky130_fd_sc_hd__conb_1
Xpicorv32_1262 VGND VGND VPWR VPWR picorv32_1262/HI eoi[20] sky130_fd_sc_hd__conb_1
X_09329_ net1659 net280 net481 VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1273 VGND VGND VPWR VPWR picorv32_1273/HI eoi[31] sky130_fd_sc_hd__conb_1
Xpicorv32_1284 VGND VGND VPWR VPWR picorv32_1284/HI trace_data[6] sky130_fd_sc_hd__conb_1
XFILLER_167_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpicorv32_1295 VGND VGND VPWR VPWR picorv32_1295/HI trace_data[17] sky130_fd_sc_hd__conb_1
X_12340_ mem_rdata_q\[24\] _06223_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__and2_1
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout997_X net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12271_ _02369_ _02448_ _06238_ _06252_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__a31o_1
XFILLER_153_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14010_ clknet_leaf_198_clk _00464_ VGND VGND VPWR VPWR cpuregs\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12175__A2 net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11222_ cpuregs\[26\]\[24\] net699 VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__or2_1
XANTENNA__08441__S net531 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13059__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11153_ net816 _05830_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__or2_1
XFILLER_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10104_ count_cycle\[38\] count_cycle\[39\] _04831_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__and3_1
X_11084_ cpuregs\[19\]\[20\] net622 net591 VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__o21a_1
XFILLER_103_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12898__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14912_ clknet_leaf_121_clk _01264_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_10035_ _04790_ net1224 _04789_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__and3b_1
XANTENNA__12883__A0 mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09272__S net485 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08551__B2 net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ clknet_leaf_11_clk _01195_ VGND VGND VPWR VPWR cpuregs\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output125_A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14774_ clknet_leaf_153_clk _00029_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12635__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ net1039 net1036 net1034 _06434_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__or4_2
X_13725_ clknet_leaf_146_clk _00179_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10937_ cpuregs\[22\]\[16\] cpuregs\[23\]\[16\] net655 VGND VGND VPWR VPWR _05621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_164_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_164_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_32_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13522__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13656_ clknet_leaf_113_clk _00110_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10661__A2 _05351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10868_ cpuregs\[22\]\[14\] cpuregs\[23\]\[14\] net664 VGND VGND VPWR VPWR _05554_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ net1199 genblk1.genblk1.pcpi_mul.next_rs2\[3\] net916 net119 VGND VGND VPWR
+ VPWR _02053_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12138__S net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13587_ net1319 VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10799_ cpuregs\[10\]\[12\] net652 VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__or2_1
XFILLER_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15326_ clknet_leaf_58_clk _01666_ VGND VGND VPWR VPWR cpuregs\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12538_ _02025_ net2534 net389 VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10881__S net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15257_ clknet_leaf_37_clk _01598_ VGND VGND VPWR VPWR cpuregs\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12469_ net1168 _06696_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12166__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14208_ clknet_leaf_25_clk _00662_ VGND VGND VPWR VPWR reg_pc\[16\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__07756__A net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08204__X alu_out\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15188_ clknet_leaf_19_clk _01537_ VGND VGND VPWR VPWR cpuregs\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14139_ clknet_leaf_126_clk _00593_ VGND VGND VPWR VPWR count_instr\[10\] sky130_fd_sc_hd__dfxtp_1
Xfanout409 _03782_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06961_ _02540_ _02539_ _02537_ _02536_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__a2bb2o_1
X_08700_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__inv_2
XANTENNA__12874__A0 mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09680_ _04474_ _04476_ _04473_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12601__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06892_ net1184 net985 VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__nand2_8
XANTENNA__09182__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08631_ genblk1.genblk1.pcpi_mul.next_rs2\[24\] net1103 genblk1.genblk1.pcpi_mul.rd\[23\]
+ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__a21o_1
XANTENNA__11725__B net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08562_ genblk1.genblk1.pcpi_mul.next_rs2\[13\] net1090 _03940_ _03942_ VGND VGND
+ VPWR VPWR _03944_ sky130_fd_sc_hd__and4_1
XFILLER_70_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07513_ count_cycle\[24\] net973 net843 _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__o211a_1
XFILLER_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_155_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_155_clk sky130_fd_sc_hd__clkbuf_8
X_08493_ net896 _03884_ _03885_ net2614 net1199 VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__a32o_1
XFILLER_62_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07444_ _02975_ _02976_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__and2_1
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__S net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07375_ latched_is_lh _02912_ _02811_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout323_A _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A net1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09114_ net1502 net320 net504 VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__mux2_1
XFILLER_136_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_946 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09045_ net330 net2426 net512 VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1232_A net1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09357__S net478 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold430 cpuregs\[21\]\[12\] VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08261__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold441 cpuregs\[13\]\[10\] VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold452 cpuregs\[29\]\[9\] VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10804__B decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold463 cpuregs\[13\]\[16\] VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 cpuregs\[24\]\[27\] VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__B1 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold485 cpuregs\[23\]\[29\] VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold496 cpuregs\[22\]\[18\] VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout910 _03879_ VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout921 net927 VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__clkbuf_4
X_09947_ net2644 net879 _04722_ net849 VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__a22o_1
Xfanout932 net933 VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__buf_2
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout480_X net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout943 _00015_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__buf_4
Xfanout954 net955 VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__clkbuf_4
Xfanout965 _02449_ VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12865__A0 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout976 net979 VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__buf_2
XANTENNA__11668__A1 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09878_ net1146 _04655_ _04656_ _04659_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__a31o_1
Xfanout987 _02379_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__clkbuf_2
Xfanout998 net999 VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__buf_2
XFILLER_85_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1130 cpuregs\[7\]\[1\] VGND VGND VPWR VPWR net2444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09092__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1141 genblk2.pcpi_div.divisor\[62\] VGND VGND VPWR VPWR net2455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1152 cpuregs\[19\]\[31\] VGND VGND VPWR VPWR net2466 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _04161_ _04164_ _04166_ _04168_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__o211a_1
Xhold1163 genblk1.genblk1.pcpi_mul.next_rs1\[31\] VGND VGND VPWR VPWR net2477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1174 cpuregs\[9\]\[16\] VGND VGND VPWR VPWR net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 cpuregs\[23\]\[30\] VGND VGND VPWR VPWR net2499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 cpuregs\[9\]\[26\] VGND VGND VPWR VPWR net2510 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ genblk2.pcpi_div.dividend\[5\] genblk2.pcpi_div.divisor\[5\] VGND VGND VPWR
+ VPWR _06311_ sky130_fd_sc_hd__and2b_1
XANTENNA__12617__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08297__A0 net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _06245_ _06247_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_146_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout912_X net912 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13510_ net1855 net312 net421 VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__mux2_1
X_10722_ net827 _05407_ _05409_ _05411_ net789 VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__a2111o_1
X_14490_ clknet_leaf_92_clk _00879_ VGND VGND VPWR VPWR instr_srli sky130_fd_sc_hd__dfxtp_1
XANTENNA__08436__S net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13441_ net570 _06105_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__nor2_1
X_10653_ _05343_ _05344_ net814 VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__mux2_1
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09797__B1 net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13372_ net569 _05820_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__nor2_1
XANTENNA__12276__B1_N net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10584_ _05251_ _05260_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__a21oi_2
Xclkload19 clknet_leaf_193_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinv_4
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15111_ clknet_leaf_72_clk _01463_ VGND VGND VPWR VPWR cpuregs\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12323_ decoded_imm\[12\] net743 _06632_ _06640_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__o22a_1
XFILLER_154_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12482__A net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12148__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09267__S net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15042_ clknet_leaf_124_clk _01394_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_12254_ net2702 net377 net364 genblk2.pcpi_div.divisor\[18\] VGND VGND VPWR VPWR
+ _01123_ sky130_fd_sc_hd__a22o_1
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11205_ net810 _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__or2_1
XANTENNA__08221__B1 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12185_ genblk2.pcpi_div.quotient_msk\[6\] net276 net2685 VGND VGND VPWR VPWR _06585_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_112_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ cpuregs\[17\]\[21\] net622 net610 _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__o211a_1
XANTENNA_output242_A net242 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13517__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11659__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12421__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11067_ _05729_ _05730_ _05747_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12320__A2 decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10018_ count_cycle\[7\] count_cycle\[8\] _04776_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__and3_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14826_ clknet_leaf_21_clk _01178_ VGND VGND VPWR VPWR cpuregs\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14757_ clknet_leaf_141_clk _00042_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12657__A _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_137_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_137_clk sky130_fd_sc_hd__clkbuf_8
X_11969_ net1043 net1041 _06423_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__or3_2
XANTENNA__06838__A1 net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13708_ clknet_leaf_107_clk _00162_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_14688_ clknet_leaf_155_clk _01073_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13639_ clknet_leaf_147_clk _00093_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07160_ count_instr\[1\] net1136 count_cycle\[33\] net1140 VGND VGND VPWR VPWR _02712_
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15309_ clknet_leaf_182_clk _01649_ VGND VGND VPWR VPWR cpuregs\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_07091_ _02648_ _02649_ _02651_ _02652_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_146_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12139__A2 net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09177__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10624__B _05316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14380__Q net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08212__B1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09801_ _04435_ _04588_ net1183 VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload10_A clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07993_ _03283_ _03503_ _03504_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__a21o_1
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09732_ _04523_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__and2_1
X_06944_ net1125 _02525_ genblk2.pcpi_div.quotient\[4\] VGND VGND VPWR VPWR _02526_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09663_ net848 _04461_ _04462_ net878 net2630 VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__a32o_1
XFILLER_54_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06875_ reg_sh\[4\] _02473_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout273_A net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08614_ genblk1.genblk1.pcpi_mul.next_rs2\[21\] net1102 _03984_ _03986_ VGND VGND
+ VPWR VPWR _03988_ sky130_fd_sc_hd__and4_1
X_09594_ _03754_ reg_next_pc\[3\] net923 VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__mux2_2
XANTENNA__09640__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08279__A0 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08545_ net887 _03927_ _03929_ net2749 net1193 VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout440_A net442 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_128_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_70_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1182_A net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13162__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10625__A2 decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08476_ _03871_ _03872_ net769 VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_42_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07427_ genblk1.genblk1.pcpi_mul.pcpi_rd\[18\] genblk2.pcpi_div.pcpi_rd\[18\] net1111
+ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout705_A net707 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1068_X net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07358_ net24 _02689_ _02694_ net6 _02812_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__o221a_1
XFILLER_136_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13398__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07289_ genblk1.genblk1.pcpi_mul.pcpi_rd\[9\] genblk2.pcpi_div.pcpi_rd\[9\] net1110
+ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1235_X net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09087__S net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13327__B2 net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09028_ net585 net2327 net514 VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__mux2_1
XFILLER_151_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 cpuregs\[13\]\[15\] VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold271 net43 VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 net48 VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 cpuregs\[20\]\[8\] VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout862_X net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10561__A1 net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout740 net742 VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkbuf_4
Xfanout751 _05120_ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__buf_2
XFILLER_120_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout762 _03877_ VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__buf_2
XANTENNA__12838__A0 _03774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07843__B net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout773 _03170_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__buf_4
X_13990_ clknet_leaf_35_clk _00444_ VGND VGND VPWR VPWR cpuregs\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout784 _03152_ VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__clkbuf_4
Xfanout795 _03151_ VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10849__C1 net826 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12941_ net537 net1848 net451 VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__mux2_1
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12872_ mem_rdata_q\[9\] net32 net963 VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__mux2_1
X_14611_ clknet_leaf_106_clk _00997_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ genblk2.pcpi_div.divisor\[14\] genblk2.pcpi_div.dividend\[14\] VGND VGND
+ VPWR VPWR _06294_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_29_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_8
X_15591_ clknet_leaf_45_clk _01927_ VGND VGND VPWR VPWR cpuregs\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12477__A net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13072__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10077__B1 net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14542_ clknet_leaf_88_clk _00928_ VGND VGND VPWR VPWR is_beq_bne_blt_bge_bltu_bgeu
+ sky130_fd_sc_hd__dfxtp_2
X_11754_ net1398 net107 net727 VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__mux2_1
XANTENNA__10709__B net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10705_ cpuregs\[14\]\[10\] cpuregs\[15\]\[10\] net664 VGND VGND VPWR VPWR _05395_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14473_ clknet_leaf_94_clk _00862_ VGND VGND VPWR VPWR instr_bgeu sky130_fd_sc_hd__dfxtp_1
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11685_ net2079 net584 net375 VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__mux2_1
X_13424_ net558 _02307_ _02327_ _04879_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__a31o_1
X_10636_ net800 _05325_ _05327_ net827 VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__o211a_1
XFILLER_139_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload108 clknet_leaf_43_clk VGND VGND VPWR VPWR clkload108/Y sky130_fd_sc_hd__inv_6
Xclkload119 clknet_leaf_75_clk VGND VGND VPWR VPWR clkload119/X sky130_fd_sc_hd__clkbuf_8
X_13355_ net959 _02266_ _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__and3_1
XFILLER_155_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10567_ cpuregs\[28\]\[6\] cpuregs\[29\]\[6\] net670 VGND VGND VPWR VPWR _05261_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12416__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13318__B2 net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12306_ decoded_imm\[20\] net733 net559 mem_rdata_q\[20\] net532 VGND VGND VPWR VPWR
+ _01154_ sky130_fd_sc_hd__a221o_1
X_13286_ _04977_ _04979_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__xor2_1
X_10498_ _05195_ _05196_ net805 VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__mux2_1
X_15025_ clknet_leaf_140_clk net1355 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12237_ net2579 net385 net371 genblk2.pcpi_div.divisor\[1\] VGND VGND VPWR VPWR _01106_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10537__D1 net790 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12168_ genblk2.pcpi_div.quotient_msk\[27\] net380 net368 net2843 VGND VGND VPWR
+ VPWR _01069_ sky130_fd_sc_hd__a22o_1
XFILLER_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10731__Y _05421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11119_ cpuregs\[8\]\[21\] net661 VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__or2_1
XFILLER_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12099_ net867 _06541_ _06543_ _06544_ net275 VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__o221a_1
XFILLER_49_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 mem_rdata[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_4
XFILLER_64_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14809_ clknet_leaf_77_clk _01161_ VGND VGND VPWR VPWR decoded_imm\[13\] sky130_fd_sc_hd__dfxtp_2
X_08330_ reg_pc\[3\] reg_pc\[2\] VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__xor2_1
XANTENNA__11265__C1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10178__Y _04884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06816__C instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14375__Q net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08261_ net1035 _03714_ net980 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__mux2_2
X_07212_ _02745_ _02750_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__nand2_1
XFILLER_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08192_ _03313_ _03680_ net935 _03312_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07236__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07143_ net1 net130 _02695_ net8 _02692_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__a221o_1
XANTENNA__07236__B2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10635__A net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07074_ genblk2.pcpi_div.quotient\[21\] _02628_ net1117 VGND VGND VPWR VPWR _02638_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__13309__B2 net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10791__B2 net797 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07539__A2 net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_A net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout488_A _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13157__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07976_ _03306_ _03489_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__nand2_1
XFILLER_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09715_ _04428_ _04509_ net1183 VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__mux2_1
XFILLER_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06927_ genblk2.pcpi_div.dividend\[1\] genblk2.pcpi_div.dividend\[0\] net1126 VGND
+ VGND VPWR VPWR _02512_ sky130_fd_sc_hd__and3_1
XANTENNA__12996__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout655_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_X net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09646_ _03861_ reg_next_pc\[29\] net924 VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__mux2_2
X_06858_ instr_sw instr_sh instr_sb _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__or4b_1
XANTENNA__10846__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09370__S net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09577_ net2855 _04412_ net1238 VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06789_ net254 VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout822_A net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_X net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_X net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08528_ _03913_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__nand2_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08459_ reg_pc\[28\] _03855_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout610_X net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11470_ cpuregs\[27\]\[30\] net637 net598 _06139_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__o211a_1
XFILLER_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10421_ _02379_ net880 _05123_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__and3_1
XFILLER_137_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13140_ net1463 net526 net431 VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__mux2_1
X_10352_ _05045_ _05048_ _03171_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__o21a_1
XFILLER_118_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13071_ net544 net2205 net440 VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__mux2_1
XFILLER_140_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10283_ _04988_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_76_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12022_ net3043 _06478_ net269 VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__mux2_1
XANTENNA__12523__A2 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11731__B1 _06243_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13067__S net442 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout570 _05040_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__buf_2
Xfanout581 _03753_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__clkbuf_2
Xfanout592 net596 VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__clkbuf_2
X_13973_ clknet_leaf_190_clk _00427_ VGND VGND VPWR VPWR cpuregs\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12287__B2 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12924_ net291 net2463 net458 VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__mux2_1
XANTENNA__10837__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09280__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07702__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12039__A1 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15643_ clknet_leaf_13_clk _01979_ VGND VGND VPWR VPWR cpuregs\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_85_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12855_ net306 net2395 net462 VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__mux2_1
XANTENNA_output205_A net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11806_ _06275_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__or2_1
X_15574_ clknet_leaf_12_clk _01910_ VGND VGND VPWR VPWR cpuregs\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12786_ net1219 genblk1.genblk1.pcpi_mul.next_rs1\[54\] net2236 net907 net764 VGND
+ VGND VPWR VPWR _01425_ sky130_fd_sc_hd__a221o_1
XANTENNA__11542__C net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14525_ clknet_leaf_76_clk _00914_ VGND VGND VPWR VPWR decoded_imm_j\[15\] sky130_fd_sc_hd__dfxtp_1
X_11737_ net1736 net119 net727 VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__mux2_1
XANTENNA__13530__S net416 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10470__B1 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14456_ clknet_leaf_90_clk _00845_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dfxtp_1
X_11668_ decoded_imm\[0\] net734 _06224_ _06225_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__a211o_1
X_13407_ net1004 net756 net558 _02290_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__o211a_1
X_10619_ cpuregs\[26\]\[7\] net668 VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_12_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14387_ clknet_leaf_84_clk _00808_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dfxtp_2
XANTENNA__07748__B net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11599_ net741 _06198_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__nor2_1
X_13338_ net568 _05675_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_94_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10174__B net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11985__S net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13269_ _02187_ _02188_ _02192_ net395 net1033 VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_149_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15008_ clknet_leaf_115_clk _01360_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07764__A net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08194__A2 net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07830_ _03340_ _03343_ _03347_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__or3_1
Xhold1707 genblk2.pcpi_div.dividend\[18\] VGND VGND VPWR VPWR net3021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1718 instr_xor VGND VGND VPWR VPWR net3032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1729 genblk2.pcpi_div.dividend\[14\] VGND VGND VPWR VPWR net3043 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_127_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07761_ net1181 net1053 VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__xor2_1
XFILLER_110_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09500_ _04363_ _04364_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__nor2_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07692_ _03210_ _03211_ net802 VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__mux2_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07154__B1 net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09190__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09431_ net2831 _04316_ net1225 VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13227__B1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09362_ net1903 net280 net478 VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__mux2_1
XFILLER_21_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08313_ net961 _03740_ net548 _00814_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07457__A1 net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09293_ net2499 net283 net486 VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__mux2_1
XANTENNA__07457__B2 net1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11253__A2 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ net254 net941 _03703_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__a21o_1
XFILLER_21_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08175_ _03660_ _03666_ VGND VGND VPWR VPWR alu_out\[26\] sky130_fd_sc_hd__or2_1
XANTENNA_fanout403_A net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07126_ genblk2.pcpi_div.quotient\[30\] _02680_ net952 VGND VGND VPWR VPWR _02682_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_119_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07057_ net1117 _02622_ genblk2.pcpi_div.dividend\[20\] VGND VGND VPWR VPWR _02623_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_37_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput140 net140 VGND VGND VPWR VPWR mem_wdata[14] sky130_fd_sc_hd__buf_2
Xoutput151 net151 VGND VGND VPWR VPWR mem_wdata[24] sky130_fd_sc_hd__buf_2
XANTENNA__09365__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput162 net162 VGND VGND VPWR VPWR mem_wdata[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput173 net173 VGND VGND VPWR VPWR pcpi_insn[11] sky130_fd_sc_hd__buf_2
Xoutput184 net184 VGND VGND VPWR VPWR pcpi_insn[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput195 net195 VGND VGND VPWR VPWR pcpi_insn[31] sky130_fd_sc_hd__buf_2
XANTENNA_fanout393_X net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A _03170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1100_X net1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07959_ _03284_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nand2_1
XFILLER_29_966 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10819__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10970_ cpuregs\[9\]\[17\] net621 net605 _05652_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__o211a_1
XFILLER_83_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09629_ reg_pc\[20\] net877 _04441_ net847 VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__a22o_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout825_X net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12640_ net2970 net893 _02069_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__a21o_1
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12571_ _02050_ net2589 net389 VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_50_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_51_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14310_ clknet_leaf_101_clk _00764_ VGND VGND VPWR VPWR count_cycle\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07849__A net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11522_ mem_rdata_q\[15\] net2238 net742 VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__mux2_1
X_15290_ clknet_leaf_30_clk _01631_ VGND VGND VPWR VPWR cpuregs\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12474__B net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14241_ clknet_leaf_27_clk _00695_ VGND VGND VPWR VPWR reg_next_pc\[18\] sky130_fd_sc_hd__dfxtp_1
X_11453_ cpuregs\[11\]\[30\] net637 net598 _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__o211a_1
X_10404_ net1161 _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__nor2_1
X_14172_ clknet_leaf_111_clk _00626_ VGND VGND VPWR VPWR count_instr\[43\] sky130_fd_sc_hd__dfxtp_1
X_11384_ cpuregs\[24\]\[28\] net689 VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_74_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10755__B2 net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11952__B1 _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13123_ net305 net2302 net437 VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__mux2_1
X_10335_ cpuregs\[6\]\[31\] cpuregs\[7\]\[31\] net692 VGND VGND VPWR VPWR _05041_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09275__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13054_ net1461 net77 net533 VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_3_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10266_ _04936_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__nand2_1
XFILLER_79_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10507__A1 net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12005_ net205 _06459_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__or2_1
XFILLER_87_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10197_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__inv_2
XANTENNA__11180__A1 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07871__X _03389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07923__A2 net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__S net418 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13956_ clknet_leaf_40_clk _00410_ VGND VGND VPWR VPWR cpuregs\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12649__B net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12907_ net357 net1926 net455 VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__mux2_1
XANTENNA__13209__B1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13887_ clknet_leaf_2_clk _00341_ VGND VGND VPWR VPWR cpuregs\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10691__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12838_ _03774_ net2345 net460 VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__mux2_1
X_15626_ clknet_leaf_29_clk _01962_ VGND VGND VPWR VPWR cpuregs\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07439__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12769_ net1219 net2432 net2594 net906 net763 VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__a221o_1
X_15557_ clknet_leaf_56_clk _01893_ VGND VGND VPWR VPWR cpuregs\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07439__B2 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12665__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08100__A2 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07759__A net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14508_ clknet_leaf_80_clk _00897_ VGND VGND VPWR VPWR decoded_imm_j\[4\] sky130_fd_sc_hd__dfxtp_2
X_15488_ clknet_leaf_59_clk _01824_ VGND VGND VPWR VPWR cpuregs\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08354__S net529 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10994__A1 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput20 mem_rdata[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
Xinput31 mem_rdata[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
X_14439_ clknet_leaf_64_clk net2738 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dfxtp_1
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold804 cpuregs\[27\]\[31\] VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 cpuregs\[20\]\[6\] VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 cpuregs\[2\]\[11\] VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 cpuregs\[2\]\[17\] VGND VGND VPWR VPWR net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07611__A1 net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold848 cpuregs\[9\]\[14\] VGND VGND VPWR VPWR net2162 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ net1129 _04451_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__nand2_1
XANTENNA__12604__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07611__B2 net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10913__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold859 genblk2.pcpi_div.divisor\[31\] VGND VGND VPWR VPWR net2173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09185__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08931_ net1633 _04242_ net944 VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__mux2_1
XFILLER_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11728__B net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08862_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__inv_2
Xhold1504 genblk2.pcpi_div.divisor\[19\] VGND VGND VPWR VPWR net2818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1515 genblk2.pcpi_div.quotient\[15\] VGND VGND VPWR VPWR net2829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _01060_ VGND VGND VPWR VPWR net2840 sky130_fd_sc_hd__dlygate4sd3_1
X_07813_ net248 net1009 VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__or2_1
Xhold1537 count_cycle\[22\] VGND VGND VPWR VPWR net2851 sky130_fd_sc_hd__dlygate4sd3_1
X_08793_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__inv_2
XFILLER_85_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1548 count_cycle\[53\] VGND VGND VPWR VPWR net2862 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1559 genblk2.pcpi_div.divisor\[29\] VGND VGND VPWR VPWR net2873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07744_ net775 _03254_ _03262_ _03246_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a31oi_4
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07675_ cpuregs\[5\]\[3\] net623 net811 _03194_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__o211a_1
XFILLER_65_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout353_A _03794_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1095_A net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07142__A3 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09414_ count_instr\[3\] count_instr\[2\] _04303_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__and3_1
XFILLER_34_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09345_ net1486 net343 net475 VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__mux2_1
XANTENNA__10794__S net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_A net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout618_A net620 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13170__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10434__B1 net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07669__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09276_ net1611 net347 net484 VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__mux2_1
XANTENNA__08264__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08227_ net1056 net1173 net239 net1054 VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__a22o_1
XANTENNA__07388__B decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_X net1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ _03292_ net933 _03641_ _03651_ VGND VGND VPWR VPWR alu_out\[24\] sky130_fd_sc_hd__a211o_1
XANTENNA_fanout987_A _02379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07109_ genblk2.pcpi_div.dividend\[27\] genblk2.pcpi_div.dividend\[26\] _02657_ net1123
+ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__o31a_1
XFILLER_134_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08089_ _03347_ _03582_ _03398_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__o21a_1
XANTENNA__09095__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10120_ count_cycle\[44\] count_cycle\[45\] _04841_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout775_X net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08158__A2 net933 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10051_ count_cycle\[20\] _04798_ net1235 VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__o21ai_1
XFILLER_103_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13439__B1 net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13810_ clknet_leaf_28_clk _00264_ VGND VGND VPWR VPWR cpuregs\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14790_ clknet_leaf_109_clk _00049_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_wait_q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13741_ clknet_leaf_105_clk net2516 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_waiting
+ sky130_fd_sc_hd__dfxtp_4
X_10953_ _05618_ _05619_ _05636_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_104_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13672_ clknet_leaf_148_clk _00126_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10884_ net799 _05566_ _05568_ net838 VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_14_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15411_ clknet_leaf_9_clk _01750_ VGND VGND VPWR VPWR cpuregs\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12623_ genblk1.genblk1.pcpi_mul.mul_waiting net1223 net1166 VGND VGND VPWR VPWR
+ _02061_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08682__B genblk1.genblk1.pcpi_mul.next_rs2\[32\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13080__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
X_15342_ clknet_leaf_189_clk _01682_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12554_ _02037_ net2535 net389 VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__mux2_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11505_ _02380_ decoder_pseudo_trigger VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__nor2_1
XFILLER_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15273_ clknet_leaf_188_clk _01614_ VGND VGND VPWR VPWR cpuregs\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12485_ net870 _06707_ _06708_ net386 VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__a31o_1
X_14224_ clknet_leaf_78_clk _00678_ VGND VGND VPWR VPWR reg_next_pc\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11436_ net1083 _06105_ net857 VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__a21oi_1
X_14155_ clknet_leaf_100_clk _00609_ VGND VGND VPWR VPWR count_instr\[26\] sky130_fd_sc_hd__dfxtp_1
X_11367_ _06037_ _06038_ net817 VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__mux2_1
X_13106_ net526 net2248 net435 VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__mux2_1
XFILLER_98_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10318_ _05021_ _05023_ _04905_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__o21ai_2
XANTENNA__11548__B net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14086_ clknet_leaf_30_clk _00540_ VGND VGND VPWR VPWR cpuregs\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11298_ net840 _05969_ _05971_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_163_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ net1366 net90 net535 VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__mux2_1
X_10249_ decoded_imm\[2\] net1045 VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__or2_1
Xfanout1140 instr_rdcycleh VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__buf_2
XANTENNA__12350__B1 _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1151 net1152 VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__buf_1
Xfanout1162 net241 VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__buf_4
XFILLER_120_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1173 net124 VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1184 net1186 VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__buf_4
Xfanout1195 net1196 VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__buf_2
XANTENNA__07761__B net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08349__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09649__A2 net880 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_182_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14988_ clknet_leaf_119_clk _01340_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11283__B net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13939_ clknet_leaf_176_clk _00393_ VGND VGND VPWR VPWR cpuregs\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12653__B2 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09969__A net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07460_ reg_pc\[21\] decoded_imm\[21\] VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__or2_1
XFILLER_50_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11208__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15609_ clknet_leaf_42_clk _01945_ VGND VGND VPWR VPWR cpuregs\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__06883__A2 _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_197_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07391_ _02892_ _02894_ _02907_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_33_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10416__B1 net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09130_ _04281_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14383__Q net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09061_ net1572 net587 net510 VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08012_ _03354_ _03431_ _03413_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__o21a_1
XANTENNA__13366__C1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold601 cpuregs\[13\]\[1\] VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10914__Y _05599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold612 cpuregs\[7\]\[11\] VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 cpuregs\[27\]\[0\] VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold634 cpuregs\[23\]\[7\] VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold645 cpuregs\[21\]\[27\] VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold656 cpuregs\[23\]\[24\] VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 cpuregs\[13\]\[30\] VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09963_ net1150 _04735_ _04736_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__or3_1
Xhold678 cpuregs\[21\]\[29\] VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold689 cpuregs\[10\]\[20\] VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08914_ _04112_ _04114_ _04111_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__a21bo_1
XFILLER_131_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1010_A net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09894_ net1147 _04669_ _04670_ _04674_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a31o_1
XANTENNA__11144__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1301 count_instr\[23\] VGND VGND VPWR VPWR net2615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07899__A1 net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1312 genblk1.genblk1.pcpi_mul.rd\[14\] VGND VGND VPWR VPWR net2626 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__inv_2
Xhold1323 _00826_ VGND VGND VPWR VPWR net2637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12892__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10789__S net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1334 net182 VGND VGND VPWR VPWR net2648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout470_A _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1345 genblk1.genblk1.pcpi_mul.rd\[6\] VGND VGND VPWR VPWR net2659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout568_A net570 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1356 genblk1.genblk1.pcpi_mul.rdx\[56\] VGND VGND VPWR VPWR net2670 sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ _04122_ _04124_ _04117_ _04120_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__a211o_1
Xhold1367 genblk1.genblk1.pcpi_mul.rd\[0\] VGND VGND VPWR VPWR net2681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1378 genblk2.pcpi_div.divisor\[24\] VGND VGND VPWR VPWR net2692 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08259__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1389 genblk1.genblk1.pcpi_mul.rd\[34\] VGND VGND VPWR VPWR net2703 sky130_fd_sc_hd__dlygate4sd3_1
X_07727_ net794 _03245_ _03237_ net778 VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10655__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09879__A net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07658_ cpuregs\[18\]\[2\] net555 _03178_ net785 VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__o22a_1
X_07589_ reg_pc\[30\] decoded_imm\[30\] VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nand2_1
XANTENNA__10377__X _05082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_A net903 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_X net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
X_09328_ net1605 net282 net481 VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1252 VGND VGND VPWR VPWR picorv32_1252/HI eoi[10] sky130_fd_sc_hd__conb_1
XFILLER_167_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpicorv32_1263 VGND VGND VPWR VPWR picorv32_1263/HI eoi[21] sky130_fd_sc_hd__conb_1
Xpicorv32_1274 VGND VGND VPWR VPWR picorv32_1274/HI mem_addr[0] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1285 VGND VGND VPWR VPWR picorv32_1285/HI trace_data[7] sky130_fd_sc_hd__conb_1
XFILLER_21_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpicorv32_1296 VGND VGND VPWR VPWR picorv32_1296/HI trace_data[18] sky130_fd_sc_hd__conb_1
XFILLER_167_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09259_ net1513 net285 net491 VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__mux2_1
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12270_ net175 net174 _06611_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__and3_1
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11221_ cpuregs\[25\]\[24\] net640 net614 _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__o211a_1
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11152_ cpuregs\[14\]\[22\] cpuregs\[15\]\[22\] net682 VGND VGND VPWR VPWR _05830_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10103_ count_cycle\[38\] _04831_ count_cycle\[39\] VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__a21o_1
XFILLER_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11083_ cpuregs\[17\]\[20\] net624 net605 _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__o211a_1
XANTENNA_input31_A mem_rdata[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14911_ clknet_leaf_122_clk _01263_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_10034_ count_cycle\[13\] count_cycle\[14\] _04786_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__and3_1
XANTENNA__10699__S net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12883__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13075__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ clknet_leaf_41_clk _01194_ VGND VGND VPWR VPWR cpuregs\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14773_ clknet_leaf_162_clk _00028_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11985_ genblk2.pcpi_div.dividend\[8\] _06447_ net271 VGND VGND VPWR VPWR _01017_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output118_A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12635__B2 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10936_ cpuregs\[20\]\[16\] cpuregs\[21\]\[16\] net655 VGND VGND VPWR VPWR _05620_
+ sky130_fd_sc_hd__mux2_1
X_13724_ clknet_leaf_150_clk _00178_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10867_ net828 _05548_ _05550_ _05552_ net787 VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12419__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13655_ clknet_leaf_113_clk _00109_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12606_ net2759 net894 _02052_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__a21o_1
XANTENNA__13060__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13586_ net1325 VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_156_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ cpuregs\[9\]\[12\] net620 net604 _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__o211a_1
XFILLER_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12537_ genblk2.pcpi_div.divisor\[54\] _02024_ _05082_ VGND VGND VPWR VPWR _02025_
+ sky130_fd_sc_hd__mux2_1
X_15325_ clknet_leaf_35_clk _01665_ VGND VGND VPWR VPWR cpuregs\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15256_ clknet_leaf_49_clk _01597_ VGND VGND VPWR VPWR cpuregs\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07290__A2 net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12468_ net1169 _05100_ net718 VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_117_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11559__A net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11419_ _06088_ _06089_ net820 VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__mux2_1
X_14207_ clknet_leaf_176_clk _00661_ VGND VGND VPWR VPWR reg_pc\[15\] sky130_fd_sc_hd__dfxtp_1
X_15187_ clknet_leaf_179_clk _01536_ VGND VGND VPWR VPWR cpuregs\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07756__B net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12399_ net527 net1866 net471 VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__mux2_1
XANTENNA__11374__A1 net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14138_ clknet_leaf_126_clk _00592_ VGND VGND VPWR VPWR count_instr\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09319__A1 net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14069_ clknet_leaf_188_clk _00523_ VGND VGND VPWR VPWR cpuregs\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_06960_ genblk2.pcpi_div.dividend\[6\] net1125 _02538_ net949 VGND VGND VPWR VPWR
+ _02540_ sky130_fd_sc_hd__a31o_1
XFILLER_101_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07772__A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12874__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06891_ net1208 _02485_ _02487_ _02488_ _02446_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__o41a_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08630_ genblk1.genblk1.pcpi_mul.rd\[23\] genblk1.genblk1.pcpi_mul.next_rs2\[24\]
+ net1103 VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__nand3_1
XANTENNA__14378__Q net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08561_ genblk1.genblk1.pcpi_mul.next_rs2\[13\] net1090 _03940_ _03942_ VGND VGND
+ VPWR VPWR _03943_ sky130_fd_sc_hd__a22o_1
XANTENNA__11429__A2 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07512_ net1141 count_cycle\[56\] net979 _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__a211o_1
XANTENNA__09699__A decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08492_ _03881_ _03882_ _03878_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07443_ reg_pc\[20\] decoded_imm\[20\] VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nand2_1
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13051__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07374_ net7 _02694_ _02911_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__o21a_1
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09113_ net2291 net324 net506 VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__mux2_1
XANTENNA__11062__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_A net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1058_A net1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07947__A is_compare VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09638__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09044_ net334 net2267 net512 VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__mux2_1
XFILLER_164_958 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold420 cpuregs\[29\]\[16\] VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 cpuregs\[20\]\[13\] VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold442 cpuregs\[4\]\[16\] VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold453 cpuregs\[8\]\[10\] VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 cpuregs\[25\]\[5\] VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12999__S net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold475 cpuregs\[16\]\[18\] VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold486 cpuregs\[16\]\[6\] VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net903 VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__buf_2
Xhold497 cpuregs\[25\]\[18\] VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net913 VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__clkbuf_4
Xfanout922 net927 VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__buf_4
X_09946_ _04447_ _04721_ net1185 VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__mux2_1
Xfanout933 _03460_ VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1013_X net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout944 _00015_ VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12314__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09373__S net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout955 net957 VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__clkbuf_4
Xfanout966 net967 VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__clkbuf_4
Xfanout977 net979 VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_X net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1120 cpuregs\[3\]\[11\] VGND VGND VPWR VPWR net2434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09877_ net1146 _04658_ net1182 VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_5_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout988 net990 VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11408__S net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout999 net222 VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__buf_4
Xhold1131 cpuregs\[1\]\[14\] VGND VGND VPWR VPWR net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 cpuregs\[3\]\[30\] VGND VGND VPWR VPWR net2456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 net49 VGND VGND VPWR VPWR net2467 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _04166_ _04168_ _04161_ _04164_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__a211o_1
XFILLER_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1164 genblk1.genblk1.pcpi_mul.next_rs1\[35\] VGND VGND VPWR VPWR net2478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07741__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1175 genblk1.genblk1.pcpi_mul.next_rs1\[48\] VGND VGND VPWR VPWR net2489 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1186 cpuregs\[11\]\[26\] VGND VGND VPWR VPWR net2500 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ net886 _04108_ _04110_ net2682 net1193 VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__a32o_1
Xhold1197 genblk1.genblk1.pcpi_mul.next_rs1\[20\] VGND VGND VPWR VPWR net2511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12617__B2 net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_X net738 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11770_ net168 net131 net536 VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10721_ cpuregs\[27\]\[10\] net627 net594 _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__o211a_1
XANTENNA__10548__A net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13440_ _05031_ _05033_ _02342_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__o21a_1
X_10652_ cpuregs\[20\]\[8\] cpuregs\[21\]\[8\] net669 VGND VGND VPWR VPWR _05344_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13042__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13371_ _05009_ _05018_ _02281_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__o21a_1
X_10583_ net773 _05268_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__and3_1
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12322_ net1147 decoded_imm_j\[12\] net970 mem_rdata_q\[12\] VGND VGND VPWR VPWR
+ _06640_ sky130_fd_sc_hd__a22o_1
X_15110_ clknet_leaf_48_clk _01462_ VGND VGND VPWR VPWR cpuregs\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10800__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07857__A net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08452__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08305__X net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11379__A net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15041_ clknet_leaf_129_clk _01393_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_12253_ net3069 net377 net364 net2702 VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__a22o_1
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11204_ cpuregs\[14\]\[23\] cpuregs\[15\]\[23\] net661 VGND VGND VPWR VPWR _05881_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08221__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12184_ net751 _06584_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__nor2_1
XFILLER_96_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11135_ cpuregs\[16\]\[21\] net680 VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__or2_1
XFILLER_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09283__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input34_X net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11066_ net774 _05738_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__and3_1
XANTENNA__11318__S net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10017_ count_cycle\[7\] _04776_ count_cycle\[8\] VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__a21o_1
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07732__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14825_ clknet_leaf_32_clk _01177_ VGND VGND VPWR VPWR cpuregs\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13533__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13281__A1 net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14756_ clknet_leaf_122_clk _00041_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11968_ _06311_ _06327_ _06308_ _06310_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12657__B net913 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11561__B mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13707_ clknet_leaf_115_clk _00161_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06838__A2 net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_max_cap483_A _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10919_ cpuregs\[4\]\[16\] cpuregs\[5\]\[16\] net659 VGND VGND VPWR VPWR _05603_
+ sky130_fd_sc_hd__mux2_1
X_11899_ genblk2.pcpi_div.dividend\[27\] genblk2.pcpi_div.divisor\[27\] VGND VGND
+ VPWR VPWR _06370_ sky130_fd_sc_hd__and2b_1
X_14687_ clknet_leaf_155_clk _01072_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13638_ clknet_leaf_148_clk _00092_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13569_ net339 net2171 net411 VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__mux2_1
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15308_ clknet_leaf_19_clk _01648_ VGND VGND VPWR VPWR cpuregs\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07767__A net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07090_ net1121 genblk2.pcpi_div.quotient\[24\] _02650_ net952 VGND VGND VPWR VPWR
+ _02652_ sky130_fd_sc_hd__a31oi_1
XANTENNA__08215__X net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15239_ clknet_leaf_19_clk _01580_ VGND VGND VPWR VPWR cpuregs\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12544__B1 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08212__A1 _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09800_ _04584_ _04585_ _04587_ net984 VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__a22o_1
X_07992_ _03283_ _03503_ net770 VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07971__B1 net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09193__S net499 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09731_ decoded_imm_j\[9\] _04430_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__nand2_1
X_06943_ genblk2.pcpi_div.quotient\[0\] genblk2.pcpi_div.quotient\[1\] genblk2.pcpi_div.quotient\[2\]
+ genblk2.pcpi_div.quotient\[3\] VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_2_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10858__B1 net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09662_ net1187 _04423_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__or2_1
X_06874_ reg_sh\[3\] reg_sh\[2\] VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__or2_1
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07723__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08613_ genblk1.genblk1.pcpi_mul.next_rs2\[21\] net1102 _03984_ _03986_ VGND VGND
+ VPWR VPWR _03987_ sky130_fd_sc_hd__a22o_1
X_09593_ reg_pc\[2\] net878 _04423_ net848 VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__a22o_1
X_08544_ _03928_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__inv_2
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08475_ reg_pc\[31\] _03868_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout433_A net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07426_ count_cycle\[18\] net974 net844 _02960_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_114_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07357_ _02877_ _02892_ _02893_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout600_A _03153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout319_X net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09368__S net402 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08272__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13398__B _05926_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07288_ count_cycle\[9\] net971 net841 _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_96_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09027_ _03749_ net2326 net514 VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__mux2_1
XANTENNA__11338__A1 net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold250 cpuregs\[31\]\[10\] VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold261 net162 VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout590_X net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold272 cpuregs\[15\]\[29\] VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold283 cpuregs\[26\]\[30\] VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1715_A instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold294 cpuregs\[20\]\[28\] VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout730 _06244_ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__clkbuf_8
Xfanout741 net742 VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_123_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout752 net754 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__buf_2
X_09929_ net1127 _04446_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__and2_1
Xfanout763 _03877_ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__buf_1
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout855_X net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout774 _03170_ VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__clkbuf_8
Xfanout785 _03152_ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__buf_4
Xfanout796 net803 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__buf_4
X_12940_ net541 net2316 net454 VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__mux2_1
XANTENNA__07714__B1 net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12871_ mem_rdata_q\[8\] net31 net963 VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__mux2_1
XANTENNA__10977__S net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13248__D1 net1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14610_ clknet_leaf_106_clk _00996_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ genblk2.pcpi_div.divisor\[15\] genblk2.pcpi_div.dividend\[15\] VGND VGND
+ VPWR VPWR _06293_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08447__S net531 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15590_ clknet_leaf_36_clk _01926_ VGND VGND VPWR VPWR cpuregs\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__06756__A net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14541_ clknet_leaf_96_clk _00003_ VGND VGND VPWR VPWR is_sltiu_bltu_sltu sky130_fd_sc_hd__dfxtp_1
X_11753_ net1512 net106 net730 VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__mux2_1
XFILLER_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10704_ net839 _05391_ _05393_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__o21a_1
X_14472_ clknet_leaf_95_clk _00861_ VGND VGND VPWR VPWR instr_bltu sky130_fd_sc_hd__dfxtp_1
X_11684_ net1937 net586 net375 VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__mux2_1
X_10635_ net813 _05326_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__or2_1
X_13423_ net1188 net760 VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__or2_1
XFILLER_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09278__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_44_clk VGND VGND VPWR VPWR clkload109/Y sky130_fd_sc_hd__inv_8
X_13354_ _04998_ _04999_ _05001_ _02258_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__o211ai_1
XFILLER_154_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10566_ net789 _05255_ _05257_ _05259_ net777 VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_114_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12305_ mem_rdata_q\[21\] net559 _06631_ net532 VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__a211o_1
XFILLER_154_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13285_ _02201_ _02202_ _02206_ net395 net1029 VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__o32a_1
X_10497_ cpuregs\[22\]\[1\] cpuregs\[23\]\[1\] net688 VGND VGND VPWR VPWR _05196_
+ sky130_fd_sc_hd__mux2_1
X_12236_ net750 net2619 VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__nor2_1
X_15024_ clknet_leaf_139_clk net1365 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13528__S net416 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12167_ net2882 net380 net368 net2986 VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__a22o_1
XFILLER_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11118_ net810 _05794_ _05796_ net825 VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__o211a_1
XANTENNA__08211__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ net1003 net724 _06542_ net863 VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__a31o_1
X_11049_ _05717_ _05720_ _03171_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__o21a_1
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 mem_rdata[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_36_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14808_ clknet_leaf_78_clk _01160_ VGND VGND VPWR VPWR decoded_imm\[14\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__08357__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14739_ clknet_leaf_161_clk _01124_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08260_ reg_out\[7\] reg_next_pc\[7\] net921 VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__mux2_1
XFILLER_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07211_ _02751_ _02757_ _02759_ _02703_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__o22a_1
X_08191_ _03312_ net929 net966 VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__a21o_1
XFILLER_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11511__S net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09188__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07142_ net1050 _02384_ net1056 _02688_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__a31o_4
XANTENNA__07236__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07073_ genblk2.pcpi_div.dividend\[22\] net1121 _02635_ net949 VGND VGND VPWR VPWR
+ _02637_ sky130_fd_sc_hd__a31o_1
XANTENNA__07641__C1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10791__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13438__S net398 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11740__A1 net1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10543__A2 net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07975_ net1144 _03274_ _03487_ _03488_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout383_A net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09714_ _04507_ _04508_ net1149 _04506_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__a2bb2o_1
X_06926_ genblk2.pcpi_div.quotient\[0\] net1126 net2999 VGND VGND VPWR VPWR _02511_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06857_ mem_do_wdata net1232 cpu_state\[6\] _02453_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__and4b_1
X_09645_ reg_pc\[28\] net880 _04449_ net850 VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout550_A net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11482__A net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13173__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09576_ count_instr\[59\] count_instr\[58\] count_instr\[57\] _04408_ VGND VGND VPWR
+ VPWR _04413_ sky130_fd_sc_hd__and4_1
XANTENNA__08267__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13245__A1 net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06788_ net251 VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08527_ genblk1.genblk1.pcpi_mul.next_rs2\[8\] net1095 genblk1.genblk1.pcpi_mul.rd\[7\]
+ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1080_X net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout436_X net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A net821 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_X net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08458_ reg_out\[28\] alu_out_q\[28\] net1155 VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ net358 _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__nor2_1
X_08389_ net343 net2388 net529 VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout603_X net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10420_ net1088 cpu_state\[0\] VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__nor2_1
XANTENNA__09098__S net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10351_ net792 _05052_ _05054_ _05056_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_59_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12508__B1 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13070_ net572 net2160 net441 VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__mux2_1
X_10282_ _04923_ _04925_ _04926_ _04919_ _04918_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__a311o_1
XANTENNA__10519__C1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12021_ net861 _06348_ _06477_ _06476_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__a31o_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10534__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout571 _03761_ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout582 _03753_ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__buf_1
XANTENNA__13484__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12287__A2 net739 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout593 net596 VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_4
X_13972_ clknet_leaf_178_clk _00426_ VGND VGND VPWR VPWR cpuregs\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12923_ net294 net2438 net458 VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__mux2_1
XANTENNA__12692__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07163__A1 net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13083__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07163__B2 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15642_ clknet_leaf_12_clk _01978_ VGND VGND VPWR VPWR cpuregs\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13236__A1 net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12854_ net311 net2454 net461 VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_140_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11805_ genblk2.pcpi_div.dividend\[21\] genblk2.pcpi_div.divisor\[21\] VGND VGND
+ VPWR VPWR _06276_ sky130_fd_sc_hd__and2b_1
X_15573_ clknet_leaf_1_clk _01909_ VGND VGND VPWR VPWR cpuregs\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12785_ net1219 net2375 net2443 net908 net764 VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__a221o_1
X_14524_ clknet_leaf_69_clk _00913_ VGND VGND VPWR VPWR decoded_rd\[4\] sky130_fd_sc_hd__dfxtp_1
X_11736_ net1468 net1179 net729 VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__mux2_1
XFILLER_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14455_ clknet_leaf_64_clk _00844_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ is_sb_sh_sw mem_rdata_q\[7\] net745 VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__and3_1
XANTENNA__11331__S net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13406_ net570 _05964_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__nor2_1
XFILLER_127_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10618_ cpuregs\[25\]\[7\] net626 net608 _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__o211a_1
X_11598_ net741 _06196_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__nor2_1
X_14386_ clknet_leaf_85_clk _00807_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dfxtp_2
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10549_ net1078 _05242_ net855 VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__a21oi_1
X_13337_ _04992_ _04994_ _02251_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__o21a_1
XFILLER_115_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11970__A1 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13268_ net708 _02168_ _02189_ _02191_ net391 VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__a311o_1
XANTENNA__11567__A mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15007_ clknet_leaf_117_clk _01359_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12219_ genblk2.pcpi_div.quotient_msk\[23\] net273 net2766 VGND VGND VPWR VPWR _06602_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_166_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13199_ net1051 decoded_imm\[0\] net961 VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10190__B net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1708 genblk1.genblk1.pcpi_mul.next_rs2\[3\] VGND VGND VPWR VPWR net3022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1719 genblk2.pcpi_div.dividend\[28\] VGND VGND VPWR VPWR net3033 sky130_fd_sc_hd__dlygate4sd3_1
X_07760_ _03276_ _03277_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_127_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07780__A net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10289__A1 _04987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11486__B1 net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07691_ cpuregs\[30\]\[3\] cpuregs\[31\]\[3\] net677 VGND VGND VPWR VPWR _03211_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12683__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07154__A1 net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09430_ count_instr\[8\] count_instr\[7\] count_instr\[6\] _04313_ VGND VGND VPWR
+ VPWR _04318_ sky130_fd_sc_hd__and4_1
XFILLER_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14386__Q net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09361_ net1786 _03870_ net478 VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__mux2_1
X_08312_ _02369_ _02452_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__nor2_1
XFILLER_33_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09292_ net1799 net285 net487 VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__mux2_1
XFILLER_21_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07457__A2 net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09500__A _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08243_ net253 net941 _03702_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__a21o_1
XFILLER_165_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08174_ _03297_ _03664_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07125_ genblk2.pcpi_div.quotient\[30\] _02680_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__or2_1
XFILLER_134_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1040_A net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1138_A instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09646__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07090__B1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07056_ genblk2.pcpi_div.dividend\[19\] _02619_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__or2_1
Xoutput130 net130 VGND VGND VPWR VPWR mem_la_wstrb[0] sky130_fd_sc_hd__buf_2
XFILLER_115_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput141 net141 VGND VGND VPWR VPWR mem_wdata[15] sky130_fd_sc_hd__buf_2
Xoutput152 net152 VGND VGND VPWR VPWR mem_wdata[25] sky130_fd_sc_hd__buf_2
XANTENNA__13168__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput163 net163 VGND VGND VPWR VPWR mem_wdata[6] sky130_fd_sc_hd__buf_2
Xoutput174 net174 VGND VGND VPWR VPWR pcpi_insn[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput185 net185 VGND VGND VPWR VPWR pcpi_insn[22] sky130_fd_sc_hd__buf_2
XFILLER_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10516__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput196 net196 VGND VGND VPWR VPWR pcpi_insn[3] sky130_fd_sc_hd__buf_2
XFILLER_130_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11627__D mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12800__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07958_ net1180 net1051 net1178 net1049 VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__a22o_1
XANTENNA__09381__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06909_ net1066 _02475_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__and2_2
XFILLER_29_978 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout553_X net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12674__C1 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07889_ _03327_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__or2_1
XANTENNA__07145__A1 net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A net933 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07145__B2 net1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09628_ _03824_ reg_next_pc\[20\] net926 VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__mux2_2
XANTENNA__07696__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11229__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09559_ count_instr\[53\] count_instr\[52\] VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__and2_1
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout720_X net720 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_X net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12570_ genblk2.pcpi_div.divisor\[62\] _02049_ net874 VGND VGND VPWR VPWR _02050_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09842__B1 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11521_ mem_rdata_q\[14\] net3049 net740 VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__mux2_1
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07849__B net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11452_ cpuregs\[10\]\[30\] net689 VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__or2_1
X_14240_ clknet_leaf_26_clk _00694_ VGND VGND VPWR VPWR reg_next_pc\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10403_ net1162 _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__or2_1
XANTENNA__11939__X _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14171_ clknet_leaf_111_clk _00625_ VGND VGND VPWR VPWR count_instr\[42\] sky130_fd_sc_hd__dfxtp_1
X_11383_ _06053_ _06054_ net805 VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__mux2_1
XFILLER_125_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10755__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10334_ is_lui_auipc_jal _04880_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__or2_1
X_13122_ net308 net2360 net436 VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__mux2_1
XANTENNA__08460__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13078__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13053_ net1723 net76 net533 VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__mux2_1
XFILLER_127_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10265_ decoded_imm\[8\] net1033 VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__or2_1
XFILLER_87_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10507__A2 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12004_ _06299_ _06343_ _06345_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__nand3_1
XFILLER_3_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10196_ decoded_imm\[25\] net1002 VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__nor2_1
XFILLER_121_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11180__A2 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09291__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout390 _05097_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_161_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11468__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13955_ clknet_leaf_14_clk _00409_ VGND VGND VPWR VPWR cpuregs\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12649__C net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12906_ net404 net2005 net456 VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload7_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13209__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13886_ clknet_leaf_7_clk _00340_ VGND VGND VPWR VPWR cpuregs\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15625_ clknet_leaf_22_clk _01961_ VGND VGND VPWR VPWR cpuregs\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ net539 net2390 net459 VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13541__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15556_ clknet_leaf_54_clk _01892_ VGND VGND VPWR VPWR cpuregs\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07439__A2 net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12768_ net1219 genblk1.genblk1.pcpi_mul.next_rs1\[36\] net2432 net906 net763 VGND
+ VGND VPWR VPWR _01407_ sky130_fd_sc_hd__a221o_1
XANTENNA__12665__B net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14507_ clknet_leaf_92_clk _00896_ VGND VGND VPWR VPWR instr_ecall_ebreak sky130_fd_sc_hd__dfxtp_1
XANTENNA__08100__A3 net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11640__A0 decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11719_ net2710 _06236_ net547 VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__mux2_1
XANTENNA__07759__B net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15487_ clknet_leaf_35_clk _01823_ VGND VGND VPWR VPWR cpuregs\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12699_ net1217 net2527 net904 genblk1.genblk1.pcpi_mul.next_rs2\[63\] net714 VGND
+ VGND VPWR VPWR _01369_ sky130_fd_sc_hd__a221o_1
XANTENNA__10994__A2 decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput10 mem_rdata[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_4
X_14438_ clknet_leaf_64_clk net2981 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dfxtp_1
Xinput21 mem_rdata[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xinput32 mem_rdata[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10185__B net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13393__B1 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold805 cpuregs\[6\]\[31\] VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14369_ clknet_4_4_0_clk _00790_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dfxtp_2
Xhold816 cpuregs\[10\]\[28\] VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold827 cpuregs\[5\]\[16\] VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07775__A net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold838 cpuregs\[9\]\[15\] VGND VGND VPWR VPWR net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 cpuregs\[27\]\[29\] VGND VGND VPWR VPWR net2163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__A2 net1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08930_ genblk1.genblk1.pcpi_mul.rd\[3\] genblk1.genblk1.pcpi_mul.rd\[35\] net955
+ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__mux2_1
XANTENNA__11728__C net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08861_ _04189_ _04192_ _04194_ _04195_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__o211a_1
Xhold1505 genblk2.pcpi_div.quotient\[16\] VGND VGND VPWR VPWR net2819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1516 genblk1.genblk1.pcpi_mul.next_rs2\[12\] VGND VGND VPWR VPWR net2830 sky130_fd_sc_hd__dlygate4sd3_1
X_07812_ _03328_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nor2_1
XANTENNA__13448__A1 net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08792_ genblk1.genblk1.pcpi_mul.rd\[48\] genblk1.genblk1.pcpi_mul.rdx\[48\] VGND
+ VGND VPWR VPWR _04138_ sky130_fd_sc_hd__nand2_1
Xhold1527 count_cycle\[40\] VGND VGND VPWR VPWR net2841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 instr_jalr VGND VGND VPWR VPWR net2852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1549 genblk2.pcpi_div.quotient_msk\[14\] VGND VGND VPWR VPWR net2863 sky130_fd_sc_hd__dlygate4sd3_1
X_07743_ net835 _03257_ _03259_ _03261_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__a211o_1
XFILLER_65_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07674_ cpuregs\[4\]\[3\] net662 VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__or2_1
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09413_ _04305_ _04306_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__nor2_1
XFILLER_41_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout346_A _03802_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09344_ net1565 net347 net475 VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__mux2_1
XFILLER_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09275_ net1691 net350 net484 VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__mux2_1
XFILLER_166_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07669__B _03189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_A net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08226_ net1059 net1174 net1164 net942 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__a22o_1
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13384__B1 _05855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08157_ _03294_ _03649_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_91_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07108_ _02663_ _02664_ _02665_ _02666_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__o22ai_1
XANTENNA__09376__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08280__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08088_ net967 _03587_ _03338_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__o21ba_1
X_07039_ net1114 _02607_ genblk2.pcpi_div.quotient\[17\] VGND VGND VPWR VPWR _02608_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10050_ count_cycle\[20\] _04798_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__and2_1
XFILLER_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07366__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12530__S net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout935_X net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12111__A1 net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08315__B1 net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13740_ clknet_leaf_108_clk _00194_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_10952_ net772 _05627_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10985__S net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13671_ clknet_leaf_148_clk _00125_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10883_ cpuregs\[5\]\[15\] net621 net811 _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__o211a_1
X_15410_ clknet_leaf_4_clk _01749_ VGND VGND VPWR VPWR cpuregs\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ net2723 net888 _02060_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__a21o_1
XFILLER_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10425__A1 net1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15341_ clknet_leaf_166_clk _01681_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
X_12553_ genblk2.pcpi_div.divisor\[58\] _02036_ net874 VGND VGND VPWR VPWR _02037_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11504_ net1240 _06160_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__and2_1
XANTENNA__10830__D1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15272_ clknet_leaf_178_clk _01613_ VGND VGND VPWR VPWR cpuregs\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12484_ genblk2.pcpi_div.divisor\[43\] net870 VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__nor2_1
XANTENNA__13375__B1 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14223_ clknet_leaf_87_clk _00677_ VGND VGND VPWR VPWR reg_pc\[31\] sky130_fd_sc_hd__dfxtp_1
X_11435_ net1081 decoded_imm\[29\] VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__or2_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06770__Y _02378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09286__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07054__B1 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14154_ clknet_leaf_100_clk _00608_ VGND VGND VPWR VPWR count_instr\[25\] sky130_fd_sc_hd__dfxtp_1
X_11366_ cpuregs\[4\]\[28\] cpuregs\[5\]\[28\] net692 VGND VGND VPWR VPWR _06038_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output265_A net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13105_ net537 net2451 net435 VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__mux2_1
X_10317_ _04905_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__nand2_1
X_14085_ clknet_leaf_30_clk _00539_ VGND VGND VPWR VPWR cpuregs\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11297_ cpuregs\[1\]\[26\] net551 _05970_ net807 net836 VGND VGND VPWR VPWR _05971_
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ net1593 net89 net535 VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__mux2_1
X_10248_ net1051 decoded_imm\[0\] _04952_ _04950_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__a31o_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1130 net1132 VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__clkbuf_4
Xfanout1141 net1142 VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__buf_2
XANTENNA__13536__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12350__B2 mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1152 instr_jal VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11540__C_N net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10179_ instr_srl instr_srli _04883_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__or3_1
Xfanout1163 net239 VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__buf_4
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1174 net1175 VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__buf_4
Xfanout1185 net1186 VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1196 net1197 VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__buf_2
X_14987_ clknet_leaf_116_clk _01339_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13938_ clknet_leaf_26_clk _00392_ VGND VGND VPWR VPWR cpuregs\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13869_ clknet_leaf_49_clk _00323_ VGND VGND VPWR VPWR cpuregs\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15608_ clknet_leaf_1_clk _01944_ VGND VGND VPWR VPWR cpuregs\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_07390_ _02860_ _02864_ _02866_ _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__a211o_1
XANTENNA__08365__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10416__A1 net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15539_ clknet_leaf_3_clk _01875_ VGND VGND VPWR VPWR cpuregs\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07489__B decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08085__A2 net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09060_ _04273_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__nor2_4
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08011_ net967 _03349_ _03351_ net928 _03519_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__a221o_1
XFILLER_156_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold602 cpuregs\[29\]\[4\] VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 cpuregs\[8\]\[4\] VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 cpuregs\[6\]\[0\] VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 cpuregs\[2\]\[28\] VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15495__Q net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold646 cpuregs\[7\]\[13\] VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 cpuregs\[6\]\[17\] VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold668 cpuregs\[27\]\[6\] VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _04448_ _04449_ _04719_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__and3_1
Xhold679 cpuregs\[29\]\[23\] VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__dlygate4sd3_1
X_08913_ net1195 net2711 net888 _04233_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__a22o_1
X_09893_ net1147 _04671_ _04673_ net1184 VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__o31ai_1
XANTENNA__11144__A2 net859 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_A _03857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1302 _00606_ VGND VGND VPWR VPWR net2616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12341__B2 mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1313 genblk2.pcpi_div.divisor\[59\] VGND VGND VPWR VPWR net2627 sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ genblk1.genblk1.pcpi_mul.rd\[56\] genblk1.genblk1.pcpi_mul.rdx\[56\] VGND
+ VGND VPWR VPWR _04182_ sky130_fd_sc_hd__nand2_1
XANTENNA__10352__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07899__A2 _02404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06849__A net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1324 reg_next_pc\[9\] VGND VGND VPWR VPWR net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 genblk1.genblk1.pcpi_mul.rdx\[12\] VGND VGND VPWR VPWR net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 genblk1.genblk1.pcpi_mul.rd\[22\] VGND VGND VPWR VPWR net2660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 is_slli_srli_srai VGND VGND VPWR VPWR net2671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 genblk1.genblk1.pcpi_mul.rd\[42\] VGND VGND VPWR VPWR net2682 sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ genblk1.genblk1.pcpi_mul.rd\[45\] genblk1.genblk1.pcpi_mul.next_rs2\[46\]
+ net1090 VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout463_A net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1379 _01129_ VGND VGND VPWR VPWR net2693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07726_ net835 _03240_ _03242_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout630_A net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07657_ cpuregs\[19\]\[2\] net641 net601 VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout728_A _06244_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13181__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07588_ _03108_ _03111_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__or2_1
XANTENNA__08275__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09327_ net1743 net288 net482 VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1242 VGND VGND VPWR VPWR picorv32_1242/HI eoi[0] sky130_fd_sc_hd__conb_1
XANTENNA__11065__D1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08321__A_N net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1253 VGND VGND VPWR VPWR picorv32_1253/HI eoi[11] sky130_fd_sc_hd__conb_1
XANTENNA_fanout516_X net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1160_X net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1264 VGND VGND VPWR VPWR picorv32_1264/HI eoi[22] sky130_fd_sc_hd__conb_1
XFILLER_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpicorv32_1275 VGND VGND VPWR VPWR picorv32_1275/HI mem_addr[1] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1286 VGND VGND VPWR VPWR picorv32_1286/HI trace_data[8] sky130_fd_sc_hd__conb_1
XANTENNA__09895__A net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1297 VGND VGND VPWR VPWR picorv32_1297/HI trace_data[19] sky130_fd_sc_hd__conb_1
X_09258_ net1780 net289 net490 VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__mux2_1
XFILLER_167_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08209_ _03371_ _03688_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__nor2_1
X_09189_ net301 net1765 net498 VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__mux2_1
XFILLER_147_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11220_ cpuregs\[24\]\[24\] net699 VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__or2_1
XFILLER_153_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07587__A1 net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11151_ cpuregs\[12\]\[22\] cpuregs\[13\]\[22\] net682 VGND VGND VPWR VPWR _05829_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10102_ count_cycle\[38\] _04831_ _04833_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__o21a_1
XFILLER_161_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11082_ cpuregs\[16\]\[20\] net657 VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__or2_1
XFILLER_89_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10840__Y _05527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14910_ clknet_leaf_121_clk _01262_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_10033_ count_cycle\[13\] _04786_ count_cycle\[14\] VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__a21o_1
XFILLER_49_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07207__X _02756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input24_A mem_rdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14841_ clknet_leaf_1_clk _01193_ VGND VGND VPWR VPWR cpuregs\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ clknet_leaf_161_clk _00026_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_11984_ _06334_ _06446_ _06445_ net867 VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__a2bb2o_1
X_13723_ clknet_leaf_151_clk _00177_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10935_ _05606_ _05609_ _03171_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__o21a_1
XANTENNA__13091__S net442 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13654_ clknet_leaf_112_clk _00108_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10866_ cpuregs\[27\]\[14\] net625 net593 _05551_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__o211a_1
XFILLER_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12605_ net1199 genblk1.genblk1.pcpi_mul.next_rs2\[2\] net916 net1179 VGND VGND VPWR
+ VPWR _02052_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13585_ net278 net2431 net413 VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10797_ cpuregs\[8\]\[12\] net652 VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__or2_1
XFILLER_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15324_ clknet_leaf_16_clk _01664_ VGND VGND VPWR VPWR cpuregs\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12536_ net1158 _02023_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15255_ clknet_leaf_46_clk _01596_ VGND VGND VPWR VPWR cpuregs\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12467_ _06695_ net2571 net384 VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output92_A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14206_ clknet_leaf_176_clk _00660_ VGND VGND VPWR VPWR reg_pc\[14\] sky130_fd_sc_hd__dfxtp_2
X_11418_ cpuregs\[28\]\[29\] cpuregs\[29\]\[29\] net706 VGND VGND VPWR VPWR _06089_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15186_ clknet_leaf_24_clk _01535_ VGND VGND VPWR VPWR cpuregs\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12398_ net538 net1717 net472 VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__mux2_1
X_14137_ clknet_leaf_125_clk _00591_ VGND VGND VPWR VPWR count_instr\[8\] sky130_fd_sc_hd__dfxtp_1
X_11349_ cpuregs\[25\]\[27\] net639 net613 _06021_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__o211a_1
XFILLER_113_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14068_ clknet_leaf_185_clk _00522_ VGND VGND VPWR VPWR cpuregs\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12323__A1 decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07772__B net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13019_ net337 net2488 net444 VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__mux2_1
X_06890_ net1072 is_beq_bne_blt_bge_bltu_bgeu _02451_ _02380_ net1089 VGND VGND VPWR
+ VPWR _02488_ sky130_fd_sc_hd__a32o_1
XANTENNA__07735__D1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08560_ genblk1.genblk1.pcpi_mul.rd\[12\] genblk1.genblk1.pcpi_mul.rdx\[12\] VGND
+ VGND VPWR VPWR _03942_ sky130_fd_sc_hd__or2_1
XFILLER_35_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07511_ count_instr\[56\] net1133 net1137 count_instr\[24\] VGND VGND VPWR VPWR _03040_
+ sky130_fd_sc_hd__a22o_1
X_08491_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__inv_2
XFILLER_63_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07442_ reg_pc\[20\] decoded_imm\[20\] VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__or2_1
XFILLER_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07373_ net1054 _02797_ net938 VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_44_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09112_ net1835 net328 net504 VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__mux2_1
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09043_ net338 net2229 net512 VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__mux2_1
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08215__C1 net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold410 cpuregs\[6\]\[29\] VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 net161 VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10373__B is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6_0_clk_X clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold432 cpuregs\[24\]\[1\] VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 cpuregs\[16\]\[21\] VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold454 cpuregs\[22\]\[31\] VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A net1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold465 cpuregs\[14\]\[19\] VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__A2 net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold476 cpuregs\[28\]\[10\] VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1218_A net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold487 cpuregs\[21\]\[25\] VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout901 net902 VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__buf_2
Xhold498 cpuregs\[30\]\[17\] VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09945_ net1150 _04717_ _04718_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__a22o_1
Xfanout912 net913 VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__clkbuf_2
Xfanout923 net927 VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__buf_2
XANTENNA_fanout580_A _03753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout934 _03459_ VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__buf_2
Xfanout945 _00015_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__buf_4
XANTENNA__13176__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12314__B2 mem_rdata_q\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout956 net957 VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__clkbuf_4
Xfanout967 _02433_ VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__buf_4
X_09876_ _04441_ _04646_ _04657_ _04623_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__o22ai_1
XFILLER_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout978 net979 VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 cpuregs\[11\]\[19\] VGND VGND VPWR VPWR net2424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1006_X net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1121 genblk1.genblk1.pcpi_mul.pcpi_rd\[10\] VGND VGND VPWR VPWR net2435 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__clkbuf_2
XFILLER_100_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1132 reg_next_pc\[11\] VGND VGND VPWR VPWR net2446 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ genblk1.genblk1.pcpi_mul.rd\[53\] genblk1.genblk1.pcpi_mul.next_rs2\[54\]
+ net1102 VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__nand3_1
Xhold1143 cpuregs\[1\]\[26\] VGND VGND VPWR VPWR net2457 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_X net466 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1154 cpuregs\[5\]\[30\] VGND VGND VPWR VPWR net2468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1165 _01405_ VGND VGND VPWR VPWR net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 cpuregs\[9\]\[31\] VGND VGND VPWR VPWR net2490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 genblk1.genblk1.pcpi_mul.next_rs1\[34\] VGND VGND VPWR VPWR net2501 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _04109_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__inv_2
Xhold1198 reg_next_pc\[31\] VGND VGND VPWR VPWR net2512 sky130_fd_sc_hd__dlygate4sd3_1
X_07709_ reg_sh\[3\] reg_sh\[2\] VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _04050_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ cpuregs\[26\]\[10\] net668 VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__or2_1
XANTENNA__13205__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10548__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10651_ cpuregs\[22\]\[8\] cpuregs\[23\]\[8\] net668 VGND VGND VPWR VPWR _05343_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout800_X net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08018__B net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12250__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10582_ net827 _05271_ _05273_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__a211o_1
X_13370_ _05009_ _05018_ net961 VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12321_ decoded_imm\[13\] net743 _06632_ _06639_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__o22a_1
XANTENNA__07857__B net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_181_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15040_ clknet_leaf_129_clk net1329 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_170_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12252_ net2657 net377 net364 net2719 VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11203_ cpuregs\[12\]\[23\] cpuregs\[13\]\[23\] net662 VGND VGND VPWR VPWR _05880_
+ sky130_fd_sc_hd__mux2_1
X_12183_ net2529 net276 net2925 VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08221__A2 net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11134_ _05811_ _05812_ net798 VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__mux2_1
XANTENNA__08321__X _03749_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07980__A1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13086__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12305__A1 mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_196_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07980__B2 net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11065_ net831 _05741_ _05743_ _05745_ net792 VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__a2111o_1
XFILLER_95_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10016_ count_cycle\[7\] _04776_ _04778_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__o21a_1
XANTENNA_input27_X net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10867__A1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output130_A net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output228_A net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14824_ clknet_leaf_46_clk _01176_ VGND VGND VPWR VPWR cpuregs\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14755_ clknet_leaf_122_clk _00038_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ net3010 _06432_ net276 VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__mux2_1
XFILLER_32_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13706_ clknet_leaf_117_clk _00160_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11292__A1 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11561__C mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07496__B1 net979 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10918_ cpuregs\[6\]\[16\] cpuregs\[7\]\[16\] net659 VGND VGND VPWR VPWR _05602_
+ sky130_fd_sc_hd__mux2_1
X_14686_ clknet_leaf_156_clk _01071_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11898_ _06364_ _06367_ _06269_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__a21bo_1
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09237__A1 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13637_ clknet_leaf_145_clk _00091_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10849_ cpuregs\[1\]\[14\] net549 _05534_ net799 net826 VGND VGND VPWR VPWR _05535_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_119_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12241__B1 net372 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13568_ net343 net2358 net412 VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15307_ clknet_leaf_21_clk _01647_ VGND VGND VPWR VPWR cpuregs\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12519_ genblk2.pcpi_div.divisor\[50\] net872 VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__or2_1
XANTENNA__07767__B net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13499_ net1483 net356 net420 VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_149_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15238_ clknet_leaf_5_clk _01579_ VGND VGND VPWR VPWR cpuregs\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10193__B net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12544__A1 _02396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15169_ clknet_leaf_90_clk _01518_ VGND VGND VPWR VPWR mem_rdata_q\[20\] sky130_fd_sc_hd__dfxtp_2
X_07991_ net988 _03427_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__o21a_1
XFILLER_99_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11509__S net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07971__A1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09730_ decoded_imm_j\[9\] _04430_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__or2_1
X_06942_ _02521_ _02522_ _02524_ net949 VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09173__A0 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14389__Q net259 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ net1148 _04458_ _04459_ _04460_ _02380_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__a311o_1
X_06873_ instr_rdcycle net975 net1088 VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__o21a_1
XFILLER_39_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08612_ genblk1.genblk1.pcpi_mul.rd\[20\] genblk1.genblk1.pcpi_mul.rdx\[20\] VGND
+ VGND VPWR VPWR _03986_ sky130_fd_sc_hd__or2_1
X_09592_ _03752_ reg_next_pc\[2\] net923 VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__mux2_2
X_08543_ _03919_ _03922_ _03924_ _03926_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_46_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08474_ reg_out\[31\] alu_out_q\[31\] net1156 VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07425_ count_instr\[18\] net1136 net977 _02959_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__a211o_1
XANTENNA__07884__A_N net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1168_A net265 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07356_ _02878_ _02893_ _02892_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__a21bo_1
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07287_ net1139 count_cycle\[41\] net976 _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__a211o_1
XFILLER_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09026_ _03744_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__or2_1
XFILLER_108_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold240 cpuregs\[14\]\[26\] VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 cpuregs\[28\]\[13\] VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12803__S net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold262 cpuregs\[14\]\[18\] VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 cpuregs\[29\]\[6\] VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold284 cpuregs\[20\]\[20\] VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold295 cpuregs\[29\]\[3\] VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout962_A net965 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout720 _06673_ VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11419__S net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout742 _06164_ VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__buf_6
X_09928_ _04668_ _04703_ _04704_ _04687_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__a211o_1
XANTENNA__12104__A net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout753 net754 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__clkbuf_2
Xfanout764 _03877_ VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__buf_2
Xfanout775 _03170_ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__clkbuf_4
Xfanout786 _03152_ VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__buf_2
Xfanout797 net803 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__buf_2
XANTENNA__10849__B2 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_X net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09859_ _04621_ _04641_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__or2_1
XFILLER_46_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12870_ mem_rdata_q\[7\] net30 net962 VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__mux2_1
XANTENNA__13248__C1 _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11821_ genblk2.pcpi_div.dividend\[15\] genblk2.pcpi_div.divisor\[15\] VGND VGND
+ VPWR VPWR _06292_ sky130_fd_sc_hd__and2b_1
XFILLER_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14540_ clknet_leaf_96_clk net2655 VGND VGND VPWR VPWR is_slti_blt_slt sky130_fd_sc_hd__dfxtp_1
X_11752_ net2647 net105 net730 VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__mux2_1
XFILLER_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10703_ cpuregs\[1\]\[10\] net550 _05392_ net800 net828 VGND VGND VPWR VPWR _05393_
+ sky130_fd_sc_hd__a221o_1
X_14471_ clknet_leaf_95_clk _00860_ VGND VGND VPWR VPWR instr_bge sky130_fd_sc_hd__dfxtp_1
X_11683_ latched_rd\[1\] latched_rd\[0\] _04290_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__and3_1
XFILLER_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ net1000 net756 VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__or2_1
X_10634_ cpuregs\[14\]\[8\] cpuregs\[15\]\[8\] net664 VGND VGND VPWR VPWR _05326_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11026__B2 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06772__A net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11577__A2 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13353_ _05001_ _02258_ _04998_ _04999_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__a211o_1
X_10565_ cpuregs\[11\]\[6\] net629 net596 _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__o211a_1
XFILLER_154_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12304_ decoded_imm\[21\] net733 VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__and2_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07650__B1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13284_ reg_pc\[10\] net564 _02203_ _02205_ net391 VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__a2111o_1
X_10496_ cpuregs\[20\]\[1\] cpuregs\[21\]\[1\] net688 VGND VGND VPWR VPWR _05195_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15023_ clknet_leaf_140_clk _01375_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12526__B2 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12235_ genblk2.pcpi_div.quotient_msk\[31\] net275 net2618 VGND VGND VPWR VPWR _06610_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__09294__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07402__B1 _02938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12166_ net2791 net380 net368 net2882 VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__a22o_1
XFILLER_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07953__A1 net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11117_ net799 _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__or2_1
XFILLER_96_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12097_ net724 _06542_ net1003 VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__a21oi_1
XFILLER_77_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11048_ net792 _05724_ _05726_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__or4_1
Xinput8 mem_rdata[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07705__A1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07166__C1 net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13544__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14807_ clknet_leaf_77_clk _01159_ VGND VGND VPWR VPWR decoded_imm\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_91_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12999_ net1527 net280 net450 VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__mux2_1
XANTENNA__11265__A1 net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07469__B1 net1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14738_ clknet_leaf_165_clk net2770 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10188__B net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14669_ clknet_leaf_153_clk _01054_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07210_ net1139 count_cycle\[36\] count_cycle\[4\] net976 _02758_ VGND VGND VPWR
+ VPWR _02759_ sky130_fd_sc_hd__a221o_1
X_08190_ _03267_ _03673_ _03679_ VGND VGND VPWR VPWR alu_out\[28\] sky130_fd_sc_hd__a21o_1
XANTENNA__07778__A net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07141_ _02383_ net938 VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__nor2_2
XFILLER_119_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09993__A net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07072_ net1117 _02635_ genblk2.pcpi_div.dividend\[22\] VGND VGND VPWR VPWR _02636_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10528__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08197__A1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07974_ _03419_ _03425_ net989 VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__a21o_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09713_ _04427_ _04428_ _04488_ net1149 VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__a31o_1
X_06925_ genblk2.pcpi_div.quotient\[0\] net1126 genblk2.pcpi_div.quotient\[1\] VGND
+ VGND VPWR VPWR _02510_ sky130_fd_sc_hd__and3_1
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09644_ _03858_ reg_next_pc\[28\] net924 VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__mux2_2
XFILLER_56_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06856_ _02453_ _02458_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__nand2_1
XFILLER_82_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11482__B net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09575_ _04412_ net1238 _04411_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__and3b_1
XANTENNA__13245__A2 net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06787_ net1161 VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08526_ genblk1.genblk1.pcpi_mul.rd\[7\] genblk1.genblk1.pcpi_mul.next_rs2\[8\] net1095
+ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__nand3_1
XANTENNA__12453__B1 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08121__A1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08121__B2 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08457_ net293 net2458 net530 VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout710_A _02501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout429_X net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_A _03143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09379__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11702__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07408_ net9 net939 net936 VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08283__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08388_ _03800_ _03801_ net766 VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__mux2_2
XANTENNA__10826__B net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07339_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__nor2_1
XFILLER_109_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09621__B2 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10350_ cpuregs\[11\]\[31\] net638 net599 _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_59_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout798_X net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09009_ net337 net2009 net517 VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10281_ _04978_ _04982_ _04986_ _04928_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__a211o_1
X_12020_ _06294_ _06347_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__nand2_1
XANTENNA__13181__A1 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09408__A cpu_state\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout965_X net965 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11731__A2 _06242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout550 net551 VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__clkbuf_2
Xfanout561 net563 VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__buf_2
Xfanout572 _03761_ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__buf_1
XFILLER_93_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13971_ clknet_leaf_25_clk _00425_ VGND VGND VPWR VPWR cpuregs\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xfanout583 _03751_ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout594 net596 VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12922_ net297 net1793 net457 VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__mux2_1
XFILLER_74_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08458__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12692__B1 net903 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07163__A2 net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15641_ clknet_leaf_41_clk _01977_ VGND VGND VPWR VPWR cpuregs\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12853_ net313 net2429 net461 VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11804_ genblk2.pcpi_div.divisor\[21\] genblk2.pcpi_div.dividend\[21\] VGND VGND
+ VPWR VPWR _06275_ sky130_fd_sc_hd__and2b_1
X_15572_ clknet_leaf_194_clk _01908_ VGND VGND VPWR VPWR cpuregs\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12784_ net1219 genblk1.genblk1.pcpi_mul.next_rs1\[52\] net2375 net908 net764 VGND
+ VGND VPWR VPWR _01423_ sky130_fd_sc_hd__a221o_1
XANTENNA__08112__A1 net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14523_ clknet_leaf_69_clk _00912_ VGND VGND VPWR VPWR decoded_rd\[3\] sky130_fd_sc_hd__dfxtp_1
X_11735_ net1426 net1181 net727 VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__mux2_1
XANTENNA__09289__S net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14454_ clknet_leaf_55_clk _00843_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dfxtp_1
XANTENNA__10470__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11666_ mem_rdata_q\[20\] net745 _06223_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_4_14_0_clk_X clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12747__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13405_ _05024_ _05029_ _02311_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__a21oi_1
X_10617_ cpuregs\[24\]\[7\] net669 VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__or2_1
XANTENNA__12747__B2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14385_ clknet_leaf_84_clk _00806_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_12_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ is_alu_reg_imm _06181_ _06197_ net740 net2362 VGND VGND VPWR VPWR _00878_
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_12_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13336_ _04992_ _04994_ net960 VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__a21oi_1
X_10548_ net1078 decoded_imm\[5\] VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__or2_1
XFILLER_143_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13539__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13267_ net556 _02166_ _02190_ net564 reg_pc\[8\] VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__a32o_1
XANTENNA__12443__S net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10479_ cpuregs\[12\]\[1\] cpuregs\[13\]\[1\] net682 VGND VGND VPWR VPWR _05178_
+ sky130_fd_sc_hd__mux2_1
X_15006_ clknet_leaf_117_clk _01358_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_12218_ net748 net2809 VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__nor2_1
XANTENNA__11567__B mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13198_ net569 _05168_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_166_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12149_ genblk2.pcpi_div.quotient_msk\[8\] net382 net367 net2756 VGND VGND VPWR VPWR
+ _01050_ sky130_fd_sc_hd__a22o_1
Xhold1709 genblk1.genblk1.pcpi_mul.next_rs2\[31\] VGND VGND VPWR VPWR net3023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10898__S net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11583__A net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07780__B net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08368__S net529 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07690_ cpuregs\[28\]\[3\] cpuregs\[29\]\[3\] net677 VGND VGND VPWR VPWR _03210_
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07154__A2 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13227__A2 net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09360_ net1384 net287 net478 VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__mux2_1
X_08311_ _02486_ _03456_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__nor2_1
X_09291_ net2355 net289 net486 VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__mux2_1
XFILLER_21_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11522__S net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09199__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08242_ net252 net941 _03701_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__a21o_1
XFILLER_21_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15498__Q net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08173_ _03297_ _03664_ _03464_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09603__B2 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07124_ genblk2.pcpi_div.quotient\[29\] _02671_ net1123 VGND VGND VPWR VPWR _02680_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07922__A_N net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07055_ _02621_ _02620_ _02618_ net947 VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput120 net120 VGND VGND VPWR VPWR mem_la_wdata[30] sky130_fd_sc_hd__buf_2
Xoutput131 net131 VGND VGND VPWR VPWR mem_la_wstrb[1] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1033_A net1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13163__A1 _03870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput142 net142 VGND VGND VPWR VPWR mem_wdata[16] sky130_fd_sc_hd__buf_2
Xoutput153 net153 VGND VGND VPWR VPWR mem_wdata[26] sky130_fd_sc_hd__buf_2
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput164 net164 VGND VGND VPWR VPWR mem_wdata[7] sky130_fd_sc_hd__buf_2
Xoutput175 net175 VGND VGND VPWR VPWR pcpi_insn[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout493_A _04286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11174__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput186 net186 VGND VGND VPWR VPWR pcpi_insn[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput197 net197 VGND VGND VPWR VPWR pcpi_insn[4] sky130_fd_sc_hd__buf_2
XFILLER_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1200_A net1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07957_ net967 _03277_ net932 _03276_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout660_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13184__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _04884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06908_ net1316 net956 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.instr_any_mul
+ sky130_fd_sc_hd__or2_1
XANTENNA__08278__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07888_ _03324_ _03404_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07145__A2 net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14577__Q is_compare VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09627_ net3037 net877 _04440_ net847 VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__a22o_1
X_06839_ net1048 net1051 VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__or2_4
XFILLER_44_938 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout925_A net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09558_ net1237 _04400_ _04401_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__and3_1
XFILLER_52_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08509_ genblk1.genblk1.pcpi_mul.next_rs2\[5\] net1098 _03896_ _03898_ VGND VGND
+ VPWR VPWR _03899_ sky130_fd_sc_hd__a22o_1
XFILLER_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09489_ _04356_ _04357_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout713_X net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09842__A1 net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07302__C1 _02840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11520_ mem_rdata_q\[13\] net175 net740 VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11451_ cpuregs\[9\]\[30\] net637 net612 _06120_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__o211a_1
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10402_ net1163 net240 _05105_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__or3_1
X_14170_ clknet_leaf_125_clk _00624_ VGND VGND VPWR VPWR count_instr\[41\] sky130_fd_sc_hd__dfxtp_1
X_11382_ cpuregs\[30\]\[28\] cpuregs\[31\]\[28\] net690 VGND VGND VPWR VPWR _06054_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11952__A2 _02443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13121_ net313 net2343 net437 VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__mux2_1
X_10333_ net958 _05037_ _05038_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__and3_1
X_13052_ net1827 net75 net533 VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__mux2_1
X_10264_ _04948_ _04958_ _04959_ _04969_ _04947_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__o2111ai_1
XANTENNA__10291__B net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11165__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12003_ genblk2.pcpi_div.dividend\[11\] _06462_ net271 VGND VGND VPWR VPWR _01020_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08030__B1 net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10195_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__inv_2
XFILLER_79_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07881__A net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout380 net381 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__buf_2
XANTENNA__13094__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout391 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13954_ clknet_leaf_15_clk _00408_ VGND VGND VPWR VPWR cpuregs\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12905_ net409 net2117 net456 VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__mux2_1
XFILLER_47_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output210_A net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_194_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_194_clk sky130_fd_sc_hd__clkbuf_8
X_13885_ clknet_leaf_199_clk _00339_ VGND VGND VPWR VPWR cpuregs\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13209__A2 net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12836_ net542 net2448 net459 VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__mux2_1
X_15624_ clknet_leaf_31_clk _01960_ VGND VGND VPWR VPWR cpuregs\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_122_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ clknet_leaf_59_clk _01891_ VGND VGND VPWR VPWR cpuregs\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12767_ net1219 genblk1.genblk1.pcpi_mul.next_rs1\[35\] net2472 net907 net763 VGND
+ VGND VPWR VPWR _01406_ sky130_fd_sc_hd__a221o_1
XFILLER_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10979__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14506_ clknet_leaf_93_clk _00895_ VGND VGND VPWR VPWR instr_fence sky130_fd_sc_hd__dfxtp_1
XANTENNA__12665__C net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11718_ net29 net27 net28 _06227_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__and4b_1
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11640__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15486_ clknet_leaf_17_clk _01822_ VGND VGND VPWR VPWR cpuregs\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12698_ net1217 genblk1.genblk1.pcpi_mul.next_rs2\[63\] net904 net2956 net713 VGND
+ VGND VPWR VPWR _01368_ sky130_fd_sc_hd__a221o_1
X_14437_ clknet_leaf_64_clk net2637 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dfxtp_1
Xinput11 mem_rdata[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
X_11649_ decoded_imm_j\[14\] net6 net545 VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__mux2_1
Xinput22 mem_rdata[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_156_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput33 mem_ready VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
XANTENNA__13393__A1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14368_ clknet_leaf_172_clk _00789_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dfxtp_4
XFILLER_155_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold806 cpuregs\[8\]\[20\] VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 cpuregs\[18\]\[17\] VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ _04922_ _04984_ _04917_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__o21ai_1
Xhold828 cpuregs\[3\]\[10\] VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 cpuregs\[7\]\[18\] VGND VGND VPWR VPWR net2153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07775__B net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14299_ clknet_leaf_126_clk _00753_ VGND VGND VPWR VPWR count_cycle\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08860_ _04194_ _04195_ _04189_ _04192_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__a211o_1
XANTENNA__12901__S net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10903__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1506 genblk2.pcpi_div.quotient\[25\] VGND VGND VPWR VPWR net2820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07791__A net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07811_ net247 net1010 VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__nor2_1
Xhold1517 count_instr\[8\] VGND VGND VPWR VPWR net2831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08791_ net1196 net2913 net888 _04137_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__a22o_1
XFILLER_85_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13448__A2 net757 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1528 genblk1.genblk1.pcpi_mul.rd\[41\] VGND VGND VPWR VPWR net2842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1539 genblk2.pcpi_div.divisor\[11\] VGND VGND VPWR VPWR net2853 sky130_fd_sc_hd__dlygate4sd3_1
X_07742_ cpuregs\[18\]\[4\] net555 _03260_ net785 VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__o22a_1
XANTENNA__12202__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08324__A1 reg_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12120__A2 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10667__C1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07673_ cpuregs\[6\]\[3\] cpuregs\[7\]\[3\] net662 VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_185_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_185_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_80_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09412_ net3028 _04303_ net1231 VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07730__S net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09343_ net1557 net350 net475 VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__mux2_1
XFILLER_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13081__A0 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout339_A _03807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09274_ net1880 net354 net485 VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__mux2_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08225_ net1058 net1175 net238 net1055 VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__a22o_1
XFILLER_165_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1150_A net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A _04279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12187__A2 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13384__B2 is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08156_ _03294_ _03649_ net771 VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__o21ai_1
XFILLER_162_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06870__A net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08414__X _03823_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07107_ genblk2.pcpi_div.dividend\[27\] net1122 _02658_ net949 VGND VGND VPWR VPWR
+ _02666_ sky130_fd_sc_hd__a31o_1
XANTENNA__13179__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09229__Y _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10392__A net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08087_ _03337_ net930 VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nor2_1
XFILLER_106_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07038_ genblk2.pcpi_div.quotient\[16\] _02599_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__or2_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout875_A net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_X net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12811__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09392__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08989_ _02414_ net907 _04271_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout663_X net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11427__S net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12647__B1 net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12112__A net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10951_ net824 _05630_ _05632_ _05634_ net788 VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout830_X net830 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_176_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_176_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout928_X net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11951__A net873 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13670_ clknet_leaf_148_clk _00124_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10882_ cpuregs\[4\]\[15\] net659 VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__or2_1
X_12621_ net1193 genblk1.genblk1.pcpi_mul.next_rs2\[10\] net915 net1167 VGND VGND
+ VPWR VPWR _02060_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08079__B1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15340_ clknet_leaf_166_clk _01680_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_1
XANTENNA__10425__A2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12552_ net253 _02035_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11503_ net2542 _06158_ _06157_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__a21o_1
XFILLER_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15271_ clknet_leaf_25_clk _01612_ VGND VGND VPWR VPWR cpuregs\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12483_ _05103_ net715 net1165 VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09579__B1 net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14222_ clknet_leaf_67_clk _00676_ VGND VGND VPWR VPWR reg_pc\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13375__A1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11434_ _06078_ _06087_ _06104_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06780__A mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08324__X _03751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11398__A net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14770__Q genblk2.pcpi_div.pcpi_rd\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13089__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08251__A0 net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14153_ clknet_leaf_100_clk _00607_ VGND VGND VPWR VPWR count_instr\[24\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_100_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_8
X_11365_ cpuregs\[6\]\[28\] cpuregs\[7\]\[28\] net692 VGND VGND VPWR VPWR _06037_
+ sky130_fd_sc_hd__mux2_1
X_13104_ net544 net2310 net436 VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__mux2_1
X_10316_ decoded_imm\[24\] net1004 VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__or2_1
X_14084_ clknet_leaf_40_clk _00538_ VGND VGND VPWR VPWR cpuregs\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11296_ cpuregs\[2\]\[26\] cpuregs\[3\]\[26\] net702 VGND VGND VPWR VPWR _05970_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output258_A net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13035_ net1459 net86 net535 VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__mux2_1
XANTENNA__12886__A0 mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10247_ net1051 decoded_imm\[0\] _04951_ _04952_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__nand4_1
XFILLER_79_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1120 net1124 VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12350__A2 decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1131 net1132 VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1142 instr_rdcycleh VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__clkbuf_2
X_10178_ instr_srl instr_srli _04883_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__nor3_4
Xfanout1153 net1156 VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__buf_4
Xfanout1164 net238 VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__buf_4
Xfanout1175 net123 VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__buf_4
Xfanout1186 net1187 VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1197 net1198 VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__buf_2
XFILLER_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14986_ clknet_leaf_112_clk _01338_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_167_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_167_clk sky130_fd_sc_hd__clkbuf_8
X_13937_ clknet_leaf_176_clk _00391_ VGND VGND VPWR VPWR cpuregs\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13552__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13868_ clknet_leaf_53_clk _00322_ VGND VGND VPWR VPWR cpuregs\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15607_ clknet_leaf_0_clk _01943_ VGND VGND VPWR VPWR cpuregs\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12819_ net317 net2069 net465 VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__mux2_1
XFILLER_90_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13799_ clknet_leaf_71_clk _00253_ VGND VGND VPWR VPWR cpuregs\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ clknet_leaf_3_clk _01874_ VGND VGND VPWR VPWR cpuregs\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10196__B net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15469_ clknet_leaf_20_clk _01805_ VGND VGND VPWR VPWR cpuregs\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12169__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08010_ _03350_ net934 VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__nor2_1
XANTENNA__13366__A1 net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07786__A net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08234__X net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold603 cpuregs\[10\]\[30\] VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold614 cpuregs\[25\]\[8\] VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 cpuregs\[4\]\[25\] VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 cpuregs\[20\]\[1\] VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 genblk1.genblk1.pcpi_mul.next_rs1\[61\] VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold658 cpuregs\[6\]\[15\] VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _04448_ _04719_ _04449_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__a21oi_1
XFILLER_104_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold669 cpuregs\[16\]\[11\] VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08912_ _04090_ _04092_ _04089_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12877__A0 mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09892_ _04441_ _04442_ _04646_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__and3_1
XANTENNA__12341__A2 decoded_imm_j\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08843_ net1211 net2927 net900 _04181_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__a22o_1
Xhold1303 reg_next_pc\[15\] VGND VGND VPWR VPWR net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 genblk1.genblk1.pcpi_mul.rd\[10\] VGND VGND VPWR VPWR net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 reg_next_pc\[28\] VGND VGND VPWR VPWR net2639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout289_A _03860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1336 genblk1.genblk1.pcpi_mul.rd\[36\] VGND VGND VPWR VPWR net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1347 genblk2.pcpi_div.divisor\[9\] VGND VGND VPWR VPWR net2661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12629__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08774_ genblk1.genblk1.pcpi_mul.rd\[45\] genblk1.genblk1.pcpi_mul.next_rs2\[46\]
+ net1093 VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__and3_1
Xhold1358 _00924_ VGND VGND VPWR VPWR net2672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1369 genblk1.genblk1.pcpi_mul.rd\[26\] VGND VGND VPWR VPWR net2683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07725_ cpuregs\[11\]\[4\] net640 net601 _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_158_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_158_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout456_A _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11771__A _06245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13462__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_2_0_clk_X clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_A net1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07656_ cpuregs\[17\]\[2\] net641 net614 _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07587_ net1072 _03102_ _03103_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout623_A net624 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09326_ net1553 net291 net481 VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__mux2_1
XANTENNA__11604__A1 net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xpicorv32_1243 VGND VGND VPWR VPWR picorv32_1243/HI eoi[1] sky130_fd_sc_hd__conb_1
Xpicorv32_1254 VGND VGND VPWR VPWR picorv32_1254/HI eoi[12] sky130_fd_sc_hd__conb_1
XFILLER_138_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_1265 VGND VGND VPWR VPWR picorv32_1265/HI eoi[23] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1276 VGND VGND VPWR VPWR picorv32_1276/HI mem_la_addr[0] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07284__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10812__C1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09257_ net1679 net294 net490 VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1287 VGND VGND VPWR VPWR picorv32_1287/HI trace_data[9] sky130_fd_sc_hd__conb_1
XANTENNA__12806__S net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_X net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07284__B2 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1298 VGND VGND VPWR VPWR picorv32_1298/HI trace_data[20] sky130_fd_sc_hd__conb_1
XANTENNA_fanout1153_X net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11710__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_X net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08208_ _03394_ _03694_ net990 VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__a21o_1
XANTENNA__09387__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08291__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09188_ net307 net1570 net498 VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout992_A net993 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10834__B net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08233__A0 net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1738_A is_compare VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08139_ net966 _03326_ _03327_ net929 _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__a221o_1
XFILLER_135_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11150_ net840 _05825_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout780_X net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10101_ count_cycle\[38\] _04831_ net1206 VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12868__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11081_ _05759_ _05760_ net798 VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__mux2_1
XANTENNA__12541__S net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10032_ net3041 _04786_ _04788_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__o21a_1
XFILLER_88_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14840_ clknet_leaf_0_clk _01192_ VGND VGND VPWR VPWR cpuregs\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A mem_rdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14771_ clknet_leaf_164_clk _00025_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13293__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11983_ _06332_ _06333_ net862 VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_149_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_149_clk sky130_fd_sc_hd__clkbuf_8
X_13722_ clknet_leaf_151_clk _00176_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10934_ net788 _05613_ _05615_ _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__or4_1
XFILLER_72_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06775__A net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08319__X _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13653_ clknet_leaf_112_clk _00107_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10865_ cpuregs\[26\]\[14\] net664 VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__or2_1
X_12604_ net279 net2352 net469 VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__mux2_1
X_13584_ net283 net2441 net413 VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__mux2_1
X_10796_ net812 _05481_ _05483_ net826 VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15323_ clknet_leaf_43_clk _01663_ VGND VGND VPWR VPWR cpuregs\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12535_ _05113_ net719 VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__nand2_1
XFILLER_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15254_ clknet_leaf_72_clk _01595_ VGND VGND VPWR VPWR cpuregs\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12466_ genblk2.pcpi_div.divisor\[39\] _06694_ net868 VGND VGND VPWR VPWR _06695_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14205_ clknet_leaf_177_clk _00659_ VGND VGND VPWR VPWR reg_pc\[13\] sky130_fd_sc_hd__dfxtp_1
X_11417_ cpuregs\[30\]\[29\] cpuregs\[31\]\[29\] net706 VGND VGND VPWR VPWR _06088_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08224__B1 net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15185_ clknet_leaf_29_clk _01534_ VGND VGND VPWR VPWR cpuregs\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12397_ net541 net1942 net472 VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__mux2_1
XFILLER_141_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10031__B1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output85_A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09972__B1 net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14136_ clknet_leaf_125_clk _00590_ VGND VGND VPWR VPWR count_instr\[7\] sky130_fd_sc_hd__dfxtp_1
X_11348_ cpuregs\[24\]\[27\] net693 VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__or2_1
XANTENNA__10582__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13547__S net418 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12451__S net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14067_ clknet_leaf_176_clk _00521_ VGND VGND VPWR VPWR cpuregs\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11279_ net836 _05949_ _05951_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__a211o_1
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13018_ net341 net2152 net443 VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__mux2_1
XANTENNA__09724__B1 _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11531__A0 mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14969_ clknet_leaf_150_clk _01321_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_07510_ net17 net938 net937 VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08376__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08490_ _03878_ _03881_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__nor3_1
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07441_ net1074 _02966_ _02967_ _02974_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__a31o_1
XFILLER_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09996__A net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07372_ latched_is_lb latched_is_lh VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ net1725 net332 net504 VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__mux2_1
XANTENNA__11062__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13339__A1 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09042_ net342 net2403 net512 VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__mux2_1
XANTENNA__07947__C net933 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09000__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold400 cpuregs\[29\]\[17\] VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 cpuregs\[21\]\[17\] VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 net157 VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12562__A2 net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold433 cpuregs\[27\]\[10\] VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold444 cpuregs\[31\]\[14\] VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 cpuregs\[27\]\[15\] VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold466 cpuregs\[22\]\[28\] VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 net158 VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13457__S net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout902 net903 VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__clkbuf_2
X_09944_ net1150 _04719_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__nor2_1
Xhold488 cpuregs\[8\]\[12\] VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 cpuregs\[25\]\[15\] VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout913 _03875_ VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1113_A genblk2.pcpi_div.pcpi_ready VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout924 net925 VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__clkbuf_4
Xfanout935 _03459_ VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__buf_2
XANTENNA__12314__A2 decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout946 _00015_ VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input9_A mem_rdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout957 _02500_ VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__clkbuf_4
X_09875_ _04645_ _04441_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__nand2b_1
Xfanout968 _02432_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11522__A0 mem_rdata_q\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1100 cpuregs\[3\]\[22\] VGND VGND VPWR VPWR net2414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A _03761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout979 _02420_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 cpuregs\[5\]\[19\] VGND VGND VPWR VPWR net2425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1122 cpuregs\[17\]\[4\] VGND VGND VPWR VPWR net2436 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ genblk1.genblk1.pcpi_mul.rd\[53\] genblk1.genblk1.pcpi_mul.next_rs2\[54\]
+ net1102 VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__and3_1
Xhold1133 cpuregs\[9\]\[8\] VGND VGND VPWR VPWR net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 cpuregs\[18\]\[27\] VGND VGND VPWR VPWR net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 genblk1.genblk1.pcpi_mul.next_rs1\[49\] VGND VGND VPWR VPWR net2469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1166 genblk1.genblk1.pcpi_mul.next_rs1\[39\] VGND VGND VPWR VPWR net2480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 genblk1.genblk1.pcpi_mul.next_rs1\[57\] VGND VGND VPWR VPWR net2491 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _04101_ _04104_ _04106_ _04107_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__o211a_1
XFILLER_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1188 _01404_ VGND VGND VPWR VPWR net2502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13275__B1 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13192__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1199 cpuregs\[1\]\[9\] VGND VGND VPWR VPWR net2513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout459_X net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11705__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07708_ net987 _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nor2_1
XANTENNA__08286__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08688_ genblk1.genblk1.pcpi_mul.rd\[32\] genblk1.genblk1.pcpi_mul.rdx\[32\] VGND
+ VGND VPWR VPWR _04050_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13205__B _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07639_ cpuregs\[14\]\[2\] cpuregs\[15\]\[2\] net700 VGND VGND VPWR VPWR _03160_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10650_ net827 _05337_ _05339_ _05341_ net789 VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__a2111o_1
X_09309_ net1351 net354 net480 VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ cpuregs\[18\]\[6\] net553 _05274_ net780 VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__o22a_1
XANTENNA__11440__S net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12320_ net1147 decoded_imm_j\[13\] net970 mem_rdata_q\[13\] VGND VGND VPWR VPWR
+ _06639_ sky130_fd_sc_hd__a22o_1
XFILLER_167_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10800__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout995_X net995 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08206__B1 _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12251_ genblk2.pcpi_div.divisor\[14\] net377 net364 net2657 VGND VGND VPWR VPWR
+ _01120_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_151_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12002__B2 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11202_ net838 _05876_ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__o21a_1
XANTENNA__10013__B1 net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12182_ net751 _06583_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__nor2_1
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11133_ cpuregs\[22\]\[21\] cpuregs\[23\]\[21\] net680 VGND VGND VPWR VPWR _05812_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11064_ cpuregs\[27\]\[19\] net632 net597 _05744_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__o211a_1
XFILLER_89_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07717__C1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10015_ count_cycle\[7\] _04776_ net1204 VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07732__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14823_ clknet_leaf_39_clk _01175_ VGND VGND VPWR VPWR cpuregs\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12069__B2 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output123_A net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06940__B1 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06776__Y _02384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11966_ _06429_ _06431_ net868 VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__mux2_1
X_14754_ clknet_leaf_124_clk _00027_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12300__A decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13018__A0 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10917_ net1162 net853 _05600_ _05601_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__a22o_1
X_13705_ clknet_leaf_146_clk _00159_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_14685_ clknet_leaf_156_clk net2733 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11292__A2 net858 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11897_ _06364_ _06367_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__and2_1
XFILLER_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13636_ clknet_leaf_144_clk _00090_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10848_ cpuregs\[2\]\[14\] cpuregs\[3\]\[14\] net660 VGND VGND VPWR VPWR _05534_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08924__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13567_ net348 net2180 net411 VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__mux2_1
XANTENNA__12446__S net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10779_ cpuregs\[22\]\[12\] cpuregs\[23\]\[12\] net650 VGND VGND VPWR VPWR _05467_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15306_ clknet_leaf_21_clk _01646_ VGND VGND VPWR VPWR cpuregs\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12518_ _05110_ net718 net244 VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__a21bo_1
X_13498_ net1533 net404 net420 VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__mux2_1
XFILLER_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15237_ clknet_leaf_6_clk _01578_ VGND VGND VPWR VPWR cpuregs\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12449_ _02392_ _06681_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11201__C1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15168_ clknet_leaf_65_clk _01517_ VGND VGND VPWR VPWR mem_rdata_q\[19\] sky130_fd_sc_hd__dfxtp_2
XFILLER_153_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14119_ clknet_leaf_69_clk _00573_ VGND VGND VPWR VPWR cpuregs\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15099_ clknet_leaf_6_clk _01451_ VGND VGND VPWR VPWR cpuregs\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_07990_ net988 _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__nand2_1
X_06941_ genblk2.pcpi_div.quotient\[3\] _02523_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__xor2_1
XFILLER_140_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09660_ net1148 _04423_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__nor2_1
X_06872_ instr_rdcycle net975 VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__nor2_1
XANTENNA__10858__A2 net620 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07723__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08611_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__inv_2
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09591_ reg_pc\[1\] net878 _04422_ net848 VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__a22o_1
XANTENNA__11525__S net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08542_ _03924_ _03926_ _03919_ _03922_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_46_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07487__A1 net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08473_ net283 net2305 net530 VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__mux2_1
X_07424_ count_instr\[50\] net1132 net1140 count_cycle\[50\] VGND VGND VPWR VPWR _02959_
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07355_ reg_pc\[12\] decoded_imm\[12\] _02880_ _02877_ VGND VGND VPWR VPWR _02894_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout321_A _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout1063_A net1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout419_A net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07286_ count_instr\[41\] net1130 net1135 count_instr\[9\] VGND VGND VPWR VPWR _02830_
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09025_ _03743_ latched_rd\[1\] latched_rd\[0\] VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__or3b_4
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1230_A net1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08739__A1 net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09936__B1 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11767__Y _06245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold230 cpuregs\[14\]\[9\] VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 cpuregs\[22\]\[0\] VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 cpuregs\[13\]\[11\] VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 cpuregs\[23\]\[14\] VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13187__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold274 cpuregs\[12\]\[9\] VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 cpuregs\[20\]\[15\] VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold296 cpuregs\[14\]\[30\] VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10951__D1 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout710 _02501_ VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__buf_2
XFILLER_133_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout721 net723 VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__buf_2
X_09927_ _04444_ _04445_ net1127 VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__o21a_1
XANTENNA__12299__A1 mem_rdata_q\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout743 net744 VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_2
XFILLER_120_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout754 net755 VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__buf_2
XANTENNA_fanout955_A net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout765 _03877_ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__clkbuf_2
Xfanout776 net778 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__buf_4
Xfanout787 net788 VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10849__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09858_ decoded_imm_j\[17\] _04438_ _04439_ decoded_imm_j\[18\] VGND VGND VPWR VPWR
+ _04641_ sky130_fd_sc_hd__a22o_1
Xfanout798 net803 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__buf_4
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07714__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08809_ _04145_ _04148_ _04150_ _04151_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__o211a_1
X_09789_ _04434_ _04561_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06922__B1 net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ genblk2.pcpi_div.divisor\[16\] genblk2.pcpi_div.dividend\[16\] VGND VGND
+ VPWR VPWR _06291_ sky130_fd_sc_hd__xor2_1
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13216__A net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11751_ net1718 net104 net727 VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__mux2_1
XFILLER_121_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10702_ cpuregs\[2\]\[10\] cpuregs\[3\]\[10\] net673 VGND VGND VPWR VPWR _05392_
+ sky130_fd_sc_hd__mux2_1
X_14470_ clknet_leaf_95_clk _00859_ VGND VGND VPWR VPWR instr_blt sky130_fd_sc_hd__dfxtp_1
X_11682_ is_beq_bne_blt_bge_bltu_bgeu net548 _06233_ net1233 VGND VGND VPWR VPWR _00928_
+ sky130_fd_sc_hd__o211a_1
X_13421_ _04898_ _05026_ _05028_ _04897_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_153_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11026__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10633_ cpuregs\[12\]\[8\] cpuregs\[13\]\[8\] net665 VGND VGND VPWR VPWR _05325_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13352_ _02260_ _02261_ _02265_ net396 net1014 VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__o32a_1
XFILLER_139_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10564_ cpuregs\[10\]\[6\] net674 VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__or2_1
XANTENNA__10294__B net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10785__B2 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12303_ mem_rdata_q\[22\] net559 _06630_ net532 VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__a211o_1
XFILLER_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13283_ net1038 net752 _02204_ net708 VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__o211a_1
XANTENNA__07650__A1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10495_ net832 _05189_ _05191_ _05193_ net793 VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__a2111o_1
X_15022_ clknet_leaf_140_clk _01374_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12234_ net750 net2754 VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__nor2_1
XFILLER_154_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10537__A1 net830 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13097__S net442 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07402__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12165_ genblk2.pcpi_div.quotient_msk\[24\] net380 net368 net2791 VGND VGND VPWR
+ VPWR _01066_ sky130_fd_sc_hd__a22o_1
XANTENNA__10514__S net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11116_ cpuregs\[12\]\[21\] cpuregs\[13\]\[21\] net661 VGND VGND VPWR VPWR _05795_
+ sky130_fd_sc_hd__mux2_1
XFILLER_123_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12096_ net1005 _06536_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__or2_1
XANTENNA_output240_A net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10_0_clk_X clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11047_ cpuregs\[11\]\[19\] net632 net597 _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__o211a_1
XFILLER_49_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07166__B1 net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 mem_rdata[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14806_ clknet_leaf_77_clk _01158_ VGND VGND VPWR VPWR decoded_imm\[16\] sky130_fd_sc_hd__dfxtp_2
X_12998_ net1428 net284 net449 VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__mux2_1
XFILLER_45_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10469__B _05168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14737_ clknet_leaf_165_clk _01122_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11949_ genblk2.pcpi_div.dividend\[2\] _06417_ net277 VGND VGND VPWR VPWR _01011_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_71_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13560__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14668_ clknet_leaf_152_clk net2804 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07778__B net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13619_ clknet_leaf_31_clk _00074_ VGND VGND VPWR VPWR cpuregs\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14599_ clknet_leaf_115_clk _00985_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dfxtp_1
X_07140_ net1054 net1058 VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__nor2_2
XFILLER_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07071_ genblk2.pcpi_div.dividend\[21\] _02631_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__or2_1
XANTENNA__07641__A1 net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12904__S net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07794__A net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12503__B1_N net241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07973_ _03277_ _03284_ _03474_ _03276_ _03273_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__a311oi_2
X_09712_ _04427_ _04488_ _04428_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06924_ genblk2.pcpi_div.dividend\[0\] genblk2.pcpi_div.quotient\[0\] _02509_ VGND
+ VGND VPWR VPWR _00016_ sky130_fd_sc_hd__mux2_1
XANTENNA__12518__B1_N net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09643_ reg_pc\[27\] net879 _04448_ net849 VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__a22o_1
X_06855_ mem_do_rdata net1061 cpu_state\[6\] mem_do_wdata VGND VGND VPWR VPWR _02458_
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06857__B net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11255__S net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09574_ count_instr\[58\] count_instr\[57\] _04408_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__and3_1
XFILLER_55_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06786_ net240 VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_180_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ net892 _03910_ _03912_ net2659 net1201 VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_26_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12453__A1 net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13470__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08456_ _03853_ _03856_ net768 VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__mux2_2
XFILLER_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07407_ _02923_ _02930_ _02941_ _02942_ net991 VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__a311o_1
XANTENNA_clkbuf_leaf_195_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08387_ reg_pc\[14\] _03797_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__xor2_1
XANTENNA__10395__A net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07880__A1 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout703_A net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07338_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__nand2_1
XANTENNA__10767__A1 net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11964__B1 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09621__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12814__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07269_ _02811_ _02813_ net1060 VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1233_X net1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09395__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09008_ net342 net2056 net516 VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06840__C1 _02443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10280_ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__inv_2
XFILLER_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10519__B2 net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12115__A net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout860_X net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_6_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout540 _03769_ VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__buf_2
Xfanout551 _03198_ VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_45_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout562 net563 VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__buf_1
Xfanout573 _03761_ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__clkbuf_2
X_13970_ clknet_leaf_29_clk _00424_ VGND VGND VPWR VPWR cpuregs\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout584 _03751_ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__clkbuf_2
Xfanout595 net596 VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12141__B1 net372 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12921_ net301 net1956 net457 VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__mux2_1
XFILLER_100_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15640_ clknet_leaf_1_clk _01976_ VGND VGND VPWR VPWR cpuregs\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_148_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12852_ net316 net2057 net461 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__mux2_1
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _06270_ _06271_ _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__or3b_1
X_12783_ net1220 net2393 net2519 net908 net764 VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__a221o_1
X_15571_ clknet_leaf_3_clk _01907_ VGND VGND VPWR VPWR cpuregs\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12444__A1 net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08112__A2 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10455__B1 net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11734_ mem_do_wdata _02418_ _06238_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__and3_2
X_14522_ clknet_leaf_69_clk _00911_ VGND VGND VPWR VPWR decoded_rd\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07879__A net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08474__S net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08327__X _03753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14773__Q genblk2.pcpi_div.pcpi_rd\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14453_ clknet_leaf_64_clk _00842_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dfxtp_1
X_11665_ instr_jalr is_lb_lh_lw_lbu_lhu is_alu_reg_imm VGND VGND VPWR VPWR _06223_
+ sky130_fd_sc_hd__or3_2
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10616_ _05307_ _05308_ net814 VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__mux2_1
X_13404_ _05024_ _05029_ net958 VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11404__C1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14384_ clknet_leaf_84_clk _00805_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dfxtp_4
X_11596_ mem_rdata_q\[30\] _06196_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__or2_1
XFILLER_167_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13335_ _02245_ _02246_ _02250_ net396 net1018 VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__o32a_1
X_10547_ _05215_ _05224_ _05241_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__a21oi_2
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13266_ net1035 net752 VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__or2_1
X_10478_ _05174_ _05176_ net783 VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__a21o_1
XANTENNA__11168__D1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12217_ genblk2.pcpi_div.quotient_msk\[22\] net273 net2808 VGND VGND VPWR VPWR _06601_
+ sky130_fd_sc_hd__a21oi_1
X_15005_ clknet_leaf_118_clk net2846 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_124_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11567__C mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13197_ net2048 net281 net430 VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__mux2_1
XFILLER_151_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ net2909 net382 net366 net2920 VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_63_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13555__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12079_ genblk2.pcpi_div.dividend\[22\] _06527_ net273 VGND VGND VPWR VPWR _01031_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10199__B net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_08310_ net991 _03456_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__nor2_1
XFILLER_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08384__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09290_ net1818 net294 net486 VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__mux2_1
XANTENNA__07311__B1 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08241_ net251 net941 _03700_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__a21o_1
XFILLER_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08172_ _03442_ _03663_ net990 VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__mux2_1
XANTENNA__09603__A2 net882 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10749__B2 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07123_ net1124 _02678_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__nand2_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07054_ genblk2.pcpi_div.dividend\[19\] net1114 _02619_ net947 VGND VGND VPWR VPWR
+ _02621_ sky130_fd_sc_hd__a31o_1
Xoutput110 net110 VGND VGND VPWR VPWR mem_la_wdata[21] sky130_fd_sc_hd__buf_2
XFILLER_115_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput121 net121 VGND VGND VPWR VPWR mem_la_wdata[31] sky130_fd_sc_hd__buf_2
XFILLER_161_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput132 net132 VGND VGND VPWR VPWR mem_la_wstrb[2] sky130_fd_sc_hd__buf_2
Xoutput143 net143 VGND VGND VPWR VPWR mem_wdata[17] sky130_fd_sc_hd__buf_2
Xoutput154 net154 VGND VGND VPWR VPWR mem_wdata[27] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_81_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput165 net165 VGND VGND VPWR VPWR mem_wdata[8] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1026_A net1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput176 net176 VGND VGND VPWR VPWR pcpi_insn[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput187 net187 VGND VGND VPWR VPWR pcpi_insn[24] sky130_fd_sc_hd__buf_2
Xoutput198 net198 VGND VGND VPWR VPWR pcpi_insn[5] sky130_fd_sc_hd__buf_2
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout486_A _04288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13465__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07956_ _03278_ net930 VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__nor2_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06907_ genblk1.genblk1.pcpi_mul.instr_mulhsu genblk1.genblk1.pcpi_mul.instr_mulh
+ genblk1.genblk1.pcpi_mul.instr_mulhu VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__or3_1
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07887_ net1158 net1008 VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout274_X net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A net654 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06838_ net203 net1054 mem_wordsize\[0\] VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__a21o_1
X_09626_ _03819_ reg_next_pc\[19\] net922 VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__mux2_2
XFILLER_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09557_ count_instr\[52\] _04398_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_90_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11229__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_X net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06769_ net1181 VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout820_A net821 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12809__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_X net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net919 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11713__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
X_08508_ genblk1.genblk1.pcpi_mul.rd\[4\] genblk1.genblk1.pcpi_mul.rdx\[4\] VGND VGND
+ VPWR VPWR _03898_ sky130_fd_sc_hd__or2_1
XFILLER_102_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09488_ net2976 _04354_ net1239 VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08294__S net925 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08439_ _03841_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__nor2_1
XFILLER_157_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11450_ cpuregs\[8\]\[30\] net689 VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__or2_1
XANTENNA__12729__A2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10401_ net1163 _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__nor2_1
X_11381_ cpuregs\[28\]\[28\] cpuregs\[29\]\[28\] net690 VGND VGND VPWR VPWR _06053_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10853__A net797 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13120_ net318 net2259 net436 VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__mux2_1
X_10332_ _04891_ _05034_ _05035_ _05036_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__o211ai_1
XFILLER_118_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13051_ net1585 net74 net533 VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__mux2_1
X_10263_ _04966_ _04968_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__and2b_1
XFILLER_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12002_ _06461_ _06460_ _06458_ net862 VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10194_ _04898_ _04899_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__or2_1
XFILLER_120_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10912__A1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07881__B _02409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout370 _06578_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout381 net384 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_2
XFILLER_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout392 _04888_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_161_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13953_ clknet_leaf_41_clk _00407_ VGND VGND VPWR VPWR cpuregs\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10676__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12904_ net521 net2102 net456 VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__mux2_1
X_13884_ clknet_leaf_191_clk _00338_ VGND VGND VPWR VPWR cpuregs\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13209__A3 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15623_ clknet_leaf_45_clk _01959_ VGND VGND VPWR VPWR cpuregs\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12835_ net574 net2292 net462 VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output203_A net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__06784__Y _02392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_17_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ clknet_leaf_53_clk _01890_ VGND VGND VPWR VPWR cpuregs\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12766_ net1219 genblk1.genblk1.pcpi_mul.next_rs1\[34\] net2478 net907 net763 VGND
+ VGND VPWR VPWR _01405_ sky130_fd_sc_hd__a221o_1
XFILLER_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14505_ clknet_leaf_91_clk _00894_ VGND VGND VPWR VPWR instr_rdinstrh sky130_fd_sc_hd__dfxtp_1
X_11717_ is_alu_reg_imm _06235_ net547 VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__mux2_1
X_12697_ net1217 genblk1.genblk1.pcpi_mul.next_rs2\[62\] net904 net2945 net714 VGND
+ VGND VPWR VPWR _01367_ sky130_fd_sc_hd__a221o_1
X_15485_ clknet_leaf_42_clk _01821_ VGND VGND VPWR VPWR cpuregs\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14436_ clknet_leaf_89_clk net2613 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dfxtp_1
X_11648_ decoded_imm_j\[13\] net5 net545 VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__mux2_1
XANTENNA__08932__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput12 mem_rdata[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput23 mem_rdata[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xinput34 resetn VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
X_11579_ net2930 net740 net732 _06191_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__a22o_1
X_14367_ clknet_leaf_169_clk _00788_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dfxtp_2
Xhold807 cpuregs\[11\]\[10\] VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11578__B net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold818 mem_wordsize\[0\] VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13318_ _02230_ _02231_ _02235_ net395 net1022 VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__o32a_1
XFILLER_143_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold829 cpuregs\[1\]\[8\] VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_125_clk _00752_ VGND VGND VPWR VPWR count_cycle\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13249_ net1029 net758 VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11594__A mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07810_ net247 net1010 VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__and2_1
XANTENNA__07791__B net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08790_ _04135_ _04136_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__xnor2_1
Xhold1507 reg_next_pc\[5\] VGND VGND VPWR VPWR net2821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08379__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1518 count_instr\[45\] VGND VGND VPWR VPWR net2832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 genblk2.pcpi_div.quotient_msk\[28\] VGND VGND VPWR VPWR net2843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12105__B1 net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07741_ cpuregs\[19\]\[4\] net641 net601 VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__o21a_1
XFILLER_38_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07672_ decoded_imm_j\[2\] _02701_ _03192_ _02386_ _03190_ VGND VGND VPWR VPWR _06748_
+ sky130_fd_sc_hd__a221o_1
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09411_ count_instr\[2\] _04303_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__and2_1
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_09342_ net1692 net354 net476 VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__mux2_1
XANTENNA__08088__A1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09003__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09273_ net1804 net405 net485 VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__mux2_1
X_08224_ net1059 net1176 net1165 net942 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__a22o_1
XFILLER_147_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11769__A _06245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08155_ _03438_ _03648_ net990 VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout401_A _04293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12364__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06870__B net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1143_A net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11395__B2 net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07106_ net1122 _02658_ genblk2.pcpi_div.dividend\[27\] VGND VGND VPWR VPWR _02665_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_119_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08086_ _03344_ _03580_ _03586_ VGND VGND VPWR VPWR alu_out\[17\] sky130_fd_sc_hd__a21o_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07037_ net947 _02604_ _02605_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__or3_1
XFILLER_115_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07982__A net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_A net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08430__X _03836_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13195__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11708__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08289__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08988_ genblk1.genblk1.pcpi_mul.pcpi_wait_q net917 net1315 VGND VGND VPWR VPWR _04271_
+ sky130_fd_sc_hd__and3b_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07193__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07939_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__inv_2
XANTENNA__12647__B2 net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10950_ cpuregs\[27\]\[16\] net621 net591 _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__o211a_1
XFILLER_16_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09609_ reg_pc\[10\] net876 _04431_ net845 VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout823_X net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10881_ cpuregs\[6\]\[15\] cpuregs\[7\]\[15\] net659 VGND VGND VPWR VPWR _05566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13224__A net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12620_ net2668 net888 _02059_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ _05115_ net719 VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nand2_1
XANTENNA__11083__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11502_ net2542 _06159_ _06162_ _06157_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__a211o_1
X_12482_ net1165 _05103_ net715 VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__or3_1
X_15270_ clknet_leaf_25_clk _01611_ VGND VGND VPWR VPWR cpuregs\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14221_ clknet_leaf_66_clk _00675_ VGND VGND VPWR VPWR reg_pc\[29\] sky130_fd_sc_hd__dfxtp_1
X_11433_ net775 _06095_ _06103_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__and3_1
XANTENNA__07876__B net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10583__A net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14152_ clknet_leaf_100_clk net2616 VGND VGND VPWR VPWR count_instr\[23\] sky130_fd_sc_hd__dfxtp_1
X_11364_ _02397_ net860 _06036_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13103_ net572 net2183 net437 VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__mux2_1
X_10315_ _04907_ _05014_ _05017_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__o211a_1
X_14083_ clknet_leaf_14_clk _00537_ VGND VGND VPWR VPWR cpuregs\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11295_ _05967_ _05968_ net819 VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__mux2_1
XANTENNA__11138__B2 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13034_ net281 net2490 net446 VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_79_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10246_ net1047 decoded_imm\[1\] VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__or2_1
XANTENNA__12886__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10346__C1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06779__Y _02387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1110 net1111 VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__clkbuf_4
Xfanout1121 net1122 VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__buf_2
XFILLER_121_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1132 instr_rdinstrh VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__clkbuf_2
X_10177_ instr_sra instr_srai VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__or2_2
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1143 net1145 VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__clkbuf_4
Xfanout1154 net1156 VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__clkbuf_4
Xfanout1165 net237 VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__clkbuf_4
Xfanout1176 net122 VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12099__C1 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1187 decoder_trigger VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__clkbuf_4
X_14985_ clknet_leaf_108_clk _01337_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12797__X _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1198 net1205 VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_141_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13936_ clknet_leaf_76_clk _00390_ VGND VGND VPWR VPWR cpuregs\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08927__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07912__A_N net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13867_ clknet_leaf_68_clk _00321_ VGND VGND VPWR VPWR cpuregs\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11353__S net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15606_ clknet_leaf_10_clk _01942_ VGND VGND VPWR VPWR cpuregs\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13063__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12818_ net323 net2068 net464 VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__mux2_1
XFILLER_90_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13798_ clknet_leaf_33_clk _00252_ VGND VGND VPWR VPWR cpuregs\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ clknet_leaf_193_clk _01873_ VGND VGND VPWR VPWR cpuregs\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10416__A3 _05120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12749_ net2293 net897 _02108_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_139_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10821__B1 net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15468_ clknet_leaf_22_clk _01804_ VGND VGND VPWR VPWR cpuregs\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07786__B net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14419_ clknet_leaf_27_clk alu_out\[19\] VGND VGND VPWR VPWR alu_out_q\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13366__A2 net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15399_ clknet_leaf_17_clk _01738_ VGND VGND VPWR VPWR cpuregs\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08242__A1 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold604 cpuregs\[21\]\[4\] VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 cpuregs\[14\]\[5\] VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 count_instr\[63\] VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold637 cpuregs\[3\]\[18\] VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _01431_ VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 net178 VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _04732_ _04733_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12912__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_98_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08911_ net1200 net2662 net893 _04232_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__a22o_1
XANTENNA__12877__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09891_ _04657_ _04442_ _04438_ _04611_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__and4b_1
XANTENNA__11528__S net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08842_ _04179_ _04180_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__xnor2_1
Xhold1304 genblk2.pcpi_div.quotient\[31\] VGND VGND VPWR VPWR net2618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 genblk1.genblk1.pcpi_mul.next_rs2\[11\] VGND VGND VPWR VPWR net2629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1326 genblk1.genblk1.pcpi_mul.rdx\[48\] VGND VGND VPWR VPWR net2640 sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ genblk1.genblk1.pcpi_mul.next_rs2\[46\] net1090 genblk1.genblk1.pcpi_mul.rd\[45\]
+ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__a21o_1
Xhold1337 reg_next_pc\[3\] VGND VGND VPWR VPWR net2651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12629__B2 net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1348 genblk1.genblk1.pcpi_mul.rdx\[36\] VGND VGND VPWR VPWR net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 cpu_state\[0\] VGND VGND VPWR VPWR net2673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07724_ cpuregs\[10\]\[4\] net697 VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__or2_1
XFILLER_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ cpuregs\[16\]\[2\] net699 VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12359__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06865__B net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13054__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07586_ net1068 net994 _03109_ net1084 _03105_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__a221o_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09325_ net1788 net295 net481 VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__mux2_1
XFILLER_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpicorv32_1244 VGND VGND VPWR VPWR picorv32_1244/HI eoi[2] sky130_fd_sc_hd__conb_1
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_A _03148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1255 VGND VGND VPWR VPWR picorv32_1255/HI eoi[13] sky130_fd_sc_hd__conb_1
Xpicorv32_1266 VGND VGND VPWR VPWR picorv32_1266/HI eoi[24] sky130_fd_sc_hd__conb_1
X_09256_ net1421 net298 net491 VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1277 VGND VGND VPWR VPWR picorv32_1277/HI mem_la_addr[1] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06881__A _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1288 VGND VGND VPWR VPWR picorv32_1288/HI trace_data[10] sky130_fd_sc_hd__conb_1
Xpicorv32_1299 VGND VGND VPWR VPWR picorv32_1299/HI trace_data[21] sky130_fd_sc_hd__conb_1
X_08207_ _03372_ _03449_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__nand2_1
XANTENNA__12014__C1 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09187_ net309 net2241 net496 VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout404_X net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08138_ _03325_ net935 VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__nor2_1
XANTENNA__08233__A1 net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08069_ net770 _03570_ _03571_ _03565_ VGND VGND VPWR VPWR alu_out\[15\] sky130_fd_sc_hd__a31o_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12822__S net466 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07992__B1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10100_ _04831_ _04832_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__nor2_1
XFILLER_122_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11080_ cpuregs\[22\]\[20\] cpuregs\[23\]\[20\] net657 VGND VGND VPWR VPWR _05760_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout773_X net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11438__S net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10031_ count_cycle\[13\] _04786_ net1191 VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12123__A net995 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout940_X net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14770_ clknet_leaf_164_clk _00024_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ net1034 _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__xor2_1
XFILLER_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13293__B2 net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13721_ clknet_leaf_151_clk _00175_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10933_ cpuregs\[11\]\[16\] net621 net591 _05616_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__o211a_1
X_10864_ cpuregs\[25\]\[14\] net625 net607 _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__o211a_1
XANTENNA__13045__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13652_ clknet_leaf_116_clk _00106_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_12603_ net284 net2468 net469 VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__mux2_1
X_13583_ net286 net2168 net414 VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__mux2_1
X_10795_ net797 _05482_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__or2_1
XFILLER_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15322_ clknet_leaf_15_clk _01662_ VGND VGND VPWR VPWR cpuregs\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12534_ _02022_ net2690 net389 VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__mux2_1
XFILLER_158_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06791__A net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10584__Y _05278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14781__Q genblk2.pcpi_div.pcpi_rd\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15253_ clknet_leaf_47_clk _01594_ VGND VGND VPWR VPWR cpuregs\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12465_ net1169 _06693_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12556__B1 _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11359__B2 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14204_ clknet_leaf_177_clk _00658_ VGND VGND VPWR VPWR reg_pc\[12\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_117_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11416_ net795 _06082_ _06084_ _06086_ net778 VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__o41a_1
XANTENNA__08224__A1 net1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08224__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15184_ clknet_leaf_17_clk _01533_ VGND VGND VPWR VPWR cpuregs\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12396_ net571 net2032 net472 VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11347_ _06018_ _06019_ net806 VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__mux2_1
X_14135_ clknet_leaf_125_clk _00589_ VGND VGND VPWR VPWR count_instr\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12308__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output78_A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11278_ cpuregs\[18\]\[25\] net555 _05952_ net786 VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__o22a_1
X_14066_ clknet_leaf_26_clk _00520_ VGND VGND VPWR VPWR cpuregs\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09724__A1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13017_ net346 net2162 net444 VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__mux2_1
X_10229_ decoded_imm\[9\] net1031 VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__nand2_1
Xhold1 genblk1.genblk1.pcpi_mul.pcpi_wait VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13563__S net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14968_ clknet_leaf_151_clk _01320_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07414__X _02950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13919_ clknet_leaf_6_clk _00373_ VGND VGND VPWR VPWR cpuregs\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07499__C1 _03027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14899_ clknet_leaf_143_clk _01251_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_07440_ net358 _02968_ _02973_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13036__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11047__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07371_ _02907_ _02908_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__xor2_2
XANTENNA__12907__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09110_ net1912 net336 net504 VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__mux2_1
XANTENNA__12795__B1 net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07797__A net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09041_ net346 net2445 net512 VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__mux2_1
XFILLER_163_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07947__D net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12547__B1 net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08215__A1 net1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold401 cpuregs\[22\]\[5\] VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09412__B1 net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold412 cpuregs\[15\]\[26\] VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 cpuregs\[25\]\[2\] VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 genblk1.genblk1.pcpi_mul.pcpi_rd\[31\] VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 cpuregs\[12\]\[21\] VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold456 cpuregs\[10\]\[6\] VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__A1 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold467 cpuregs\[6\]\[12\] VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07736__S net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold478 cpuregs\[21\]\[6\] VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 cpuregs\[25\]\[20\] VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _04446_ _04447_ _04699_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__and3_1
Xfanout903 _03879_ VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout914 net919 VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__clkbuf_4
Xfanout925 net926 VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__buf_2
XANTENNA_fanout399_A _04293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout936 _02910_ VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__buf_2
Xfanout947 net948 VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__buf_2
XFILLER_58_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09874_ _04638_ _04644_ _04654_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__o21ai_1
Xfanout958 net959 VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10325__A2 net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout969 _02432_ VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__clkbuf_2
Xhold1101 cpuregs\[3\]\[1\] VGND VGND VPWR VPWR net2415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07037__A net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 cpuregs\[1\]\[18\] VGND VGND VPWR VPWR net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08825_ genblk1.genblk1.pcpi_mul.next_rs2\[54\] net1102 genblk1.genblk1.pcpi_mul.rd\[53\]
+ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__a21o_1
Xhold1123 cpuregs\[7\]\[22\] VGND VGND VPWR VPWR net2437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1134 cpuregs\[19\]\[5\] VGND VGND VPWR VPWR net2448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13473__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1145 cpuregs\[16\]\[0\] VGND VGND VPWR VPWR net2459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 _01419_ VGND VGND VPWR VPWR net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _01409_ VGND VGND VPWR VPWR net2481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1178 cpuregs\[19\]\[27\] VGND VGND VPWR VPWR net2492 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _04106_ _04107_ _04101_ _04104_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__a211o_1
XFILLER_39_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1189 cpuregs\[5\]\[28\] VGND VGND VPWR VPWR net2503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11286__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07707_ _03200_ _03209_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__a21oi_4
X_08687_ net1218 net2919 net905 _04049_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout733_A net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10398__A net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ cpuregs\[12\]\[2\] cpuregs\[13\]\[2\] net700 VGND VGND VPWR VPWR _03159_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11038__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07569_ count_instr\[28\] net1137 net978 _03093_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout900_A net903 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12817__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_X net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09308_ net1369 net406 net480 VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__mux2_1
XFILLER_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10580_ cpuregs\[19\]\[6\] net627 net594 VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__o21a_1
XFILLER_166_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12250__A2 net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1750_A decoded_imm_j\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10337__S net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09239_ net1469 net408 net489 VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__mux2_1
XFILLER_166_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12250_ net2677 net379 net364 net2728 VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__a22o_1
XFILLER_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08206__A1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08206__B2 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11201_ cpuregs\[1\]\[23\] net550 _05877_ net801 net829 VGND VGND VPWR VPWR _05878_
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout988_X net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11210__B1 net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12181_ genblk2.pcpi_div.quotient_msk\[4\] net276 net3011 VGND VGND VPWR VPWR _06583_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07414__C1 _02948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11132_ cpuregs\[20\]\[21\] cpuregs\[21\]\[21\] net657 VGND VGND VPWR VPWR _05811_
+ sky130_fd_sc_hd__mux2_1
Xhold990 cpuregs\[5\]\[6\] VGND VGND VPWR VPWR net2304 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09706__B2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11063_ cpuregs\[26\]\[19\] net680 VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__or2_1
XFILLER_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12710__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10014_ _04776_ _04777_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14822_ clknet_leaf_105_clk _01174_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08477__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06786__A net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14776__Q genblk2.pcpi_div.pcpi_rd\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1690 genblk1.genblk1.pcpi_mul.next_rs2\[10\] VGND VGND VPWR VPWR net3004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11277__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14753_ clknet_leaf_123_clk _00016_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11965_ net1041 _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_149_clk _00158_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_10916_ net1076 _05599_ net853 VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__a21oi_1
X_14684_ clknet_leaf_156_clk net2844 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_11896_ _06274_ _06276_ _06366_ _06365_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__o31a_1
XFILLER_60_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13635_ clknet_leaf_144_clk _00089_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10847_ net799 _05530_ _05532_ net838 VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__a211o_1
XFILLER_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13566_ net350 net2144 net411 VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__mux2_1
XANTENNA__12241__A2 net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10778_ net826 _05461_ _05463_ _05465_ net787 VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09101__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15305_ clknet_leaf_30_clk _01645_ VGND VGND VPWR VPWR cpuregs\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12517_ net244 net716 _05110_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__or3b_1
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13497_ net2165 net407 net420 VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__mux2_1
X_15236_ clknet_leaf_5_clk _01577_ VGND VGND VPWR VPWR cpuregs\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08940__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12448_ net1180 net1179 net1177 net717 VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13558__S net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09945__A1 net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15167_ clknet_leaf_64_clk _01516_ VGND VGND VPWR VPWR mem_rdata_q\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12462__S net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12544__A3 net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ net1645 net316 net361 VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__mux2_1
XFILLER_113_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11752__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14118_ clknet_leaf_30_clk _00572_ VGND VGND VPWR VPWR cpuregs\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11586__B mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15098_ clknet_leaf_18_clk _01450_ VGND VGND VPWR VPWR cpuregs\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06940_ genblk2.pcpi_div.quotient\[0\] genblk2.pcpi_div.quotient\[1\] genblk2.pcpi_div.quotient\[2\]
+ net1125 VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__o31a_1
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14049_ clknet_leaf_41_clk _00503_ VGND VGND VPWR VPWR cpuregs\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12701__B1 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06871_ net2654 instr_slti net2609 VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__or3_1
XFILLER_95_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08610_ genblk1.genblk1.pcpi_mul.rd\[20\] genblk1.genblk1.pcpi_mul.rdx\[20\] VGND
+ VGND VPWR VPWR _03984_ sky130_fd_sc_hd__nand2_1
XFILLER_55_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09590_ _03750_ reg_next_pc\[1\] net922 VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08541_ genblk1.genblk1.pcpi_mul.rd\[9\] genblk1.genblk1.pcpi_mul.next_rs2\[10\]
+ net1092 VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_46_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ net769 _03867_ _03868_ _03869_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__a31o_2
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07304__B decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07423_ net10 net939 net936 VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13322__A _02409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07354_ _02879_ _02881_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_21_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09011__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07285_ _02811_ _02828_ net1060 VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__o21a_1
X_09024_ net281 net2084 net519 VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09946__S net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13468__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold220 cpuregs\[20\]\[10\] VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12372__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold231 cpuregs\[20\]\[29\] VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 net53 VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold253 cpuregs\[30\]\[19\] VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 genblk1.genblk1.pcpi_mul.next_rs1\[27\] VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07411__A2 net1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold275 net187 VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 cpuregs\[31\]\[8\] VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout683_A net696 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout700 net701 VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__buf_2
XFILLER_160_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold297 cpuregs\[23\]\[13\] VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout711 _02083_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__clkbuf_4
Xfanout722 net723 VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09926_ _04664_ _04677_ _04686_ _04695_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__and4_1
Xfanout733 net735 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1011_X net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout744 net745 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout1109_X net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout755 net757 VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07990__A net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout766 _03747_ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__buf_4
XANTENNA_fanout850_A net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout777 net778 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__clkbuf_2
X_09857_ _04638_ _04639_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__nor2_1
XANTENNA__10703__C1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout471_X net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout788 net791 VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__buf_4
XANTENNA_fanout569_X net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout799 net803 VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__buf_2
X_08808_ _04150_ _04151_ _04145_ _04148_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__a211o_1
XANTENNA__08297__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13248__A1 net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09788_ _04561_ _04434_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__nand2b_1
X_08739_ net1197 net2924 net889 _04093_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__a22o_1
XANTENNA__12895__X _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07214__B decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11750_ net1508 net103 net728 VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__mux2_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10701_ _05389_ _05390_ net813 VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__mux2_1
X_11681_ _06171_ _06226_ net547 VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout903_X net903 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13420_ _04897_ _05028_ _05026_ _04898_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_153_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ net838 _05321_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__o21a_1
XFILLER_167_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12223__A2 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10563_ cpuregs\[9\]\[6\] net629 net609 _05256_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__o211a_1
X_13351_ net709 _02240_ _02262_ _02264_ net392 VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__a311o_1
XFILLER_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10785__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08045__B net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12302_ decoded_imm\[22\] net733 VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13282_ net1022 net758 VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__or2_1
XANTENNA__07650__A2 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10494_ cpuregs\[27\]\[1\] net636 net598 _05192_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__o211a_1
XFILLER_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15021_ clknet_leaf_122_clk _01373_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12233_ genblk2.pcpi_div.quotient_msk\[30\] net275 net2753 VGND VGND VPWR VPWR _06609_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07884__B net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12164_ genblk2.pcpi_div.quotient_msk\[23\] net380 net369 net2867 VGND VGND VPWR
+ VPWR _01065_ sky130_fd_sc_hd__a22o_1
XFILLER_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11115_ cpuregs\[14\]\[21\] cpuregs\[15\]\[21\] net661 VGND VGND VPWR VPWR _05794_
+ sky130_fd_sc_hd__mux2_1
X_12095_ _06379_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_X net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11046_ cpuregs\[10\]\[19\] net680 VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__or2_1
XANTENNA_output233_A net1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07166__A1 net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14805_ clknet_leaf_77_clk _01157_ VGND VGND VPWR VPWR decoded_imm\[17\] sky130_fd_sc_hd__dfxtp_2
X_12997_ net1638 net287 net449 VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ clknet_leaf_164_clk _01121_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07469__A2 net1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11948_ _06413_ _06414_ _06416_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08935__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ clknet_leaf_152_clk _01052_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11879_ _06292_ _06293_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__nand2b_1
XFILLER_20_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13618_ clknet_leaf_23_clk _00073_ VGND VGND VPWR VPWR cpuregs\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13411__A1 net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14598_ clknet_leaf_117_clk _00984_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07140__A net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13549_ net289 net2321 net417 VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__mux2_1
XFILLER_145_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11973__A1 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07070_ _02634_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__inv_2
XFILLER_134_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15219_ clknet_leaf_87_clk _00008_ VGND VGND VPWR VPWR cpu_state\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07794__B net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10705__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10528__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07972_ _03307_ net930 _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12920__S net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09711_ _04504_ _04505_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__xnor2_1
X_06923_ net1237 genblk1.genblk1.pcpi_mul.mul_finish VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__and2_2
XANTENNA__12686__C1 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08354__A0 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09642_ _03853_ reg_next_pc\[27\] net925 VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__mux2_2
X_06854_ instr_lbu _02456_ instr_lb net410 VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__or4b_1
XANTENNA__09006__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09573_ count_instr\[57\] _04408_ count_instr\[58\] VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a21o_1
X_06785_ net1174 VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__inv_2
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08524_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__inv_2
XANTENNA__09854__B1 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11661__A0 decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08455_ _03854_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nor2_1
XANTENNA__12367__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_A net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _03746_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07406_ _02923_ _02930_ _02941_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08386_ reg_out\[14\] alu_out_q\[14\] net1153 VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__mux2_1
XANTENNA__13402__A1 _02501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10395__B net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11413__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07337_ reg_pc\[13\] decoded_imm\[13\] VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__and2_1
XFILLER_164_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1059_X net1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10621__D1 net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07268_ net17 _02689_ _02694_ net31 _02812_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__o221a_1
XFILLER_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout898_A _03879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09007_ net346 net1705 net517 VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__mux2_1
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12508__A3 net720 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07199_ _02731_ _02733_ _02732_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10519__A2 net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12115__B net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09790__C1 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout530 _03746_ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__buf_4
Xfanout541 net544 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__clkbuf_2
Xfanout552 _03156_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__buf_4
X_09909_ _04664_ _04668_ _04677_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__a31o_1
Xfanout563 _06174_ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__buf_2
XANTENNA__12677__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout574 _03761_ VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__buf_1
XFILLER_101_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout585 _03751_ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkbuf_2
Xfanout596 _03153_ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__buf_2
X_12920_ net306 net2384 net458 VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__mux2_1
X_12851_ net321 net2260 net459 VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__mux2_1
XFILLER_15_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11802_ genblk2.pcpi_div.divisor\[22\] genblk2.pcpi_div.dividend\[22\] VGND VGND
+ VPWR VPWR _06273_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_107_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ clknet_leaf_3_clk _01906_ VGND VGND VPWR VPWR cpuregs\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12782_ net1220 net2264 net2393 net908 net765 VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__a221o_1
XANTENNA__12444__A2 net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14521_ clknet_leaf_69_clk _00910_ VGND VGND VPWR VPWR decoded_rd\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11733_ latched_rd\[4\] _06242_ _06243_ net1405 VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__a22o_1
XANTENNA__07879__B _02408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14452_ clknet_leaf_64_clk _00841_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11664_ decoded_imm_j\[3\] net16 net546 VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__mux2_1
XFILLER_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13403_ _02305_ _02306_ _02310_ net397 net1004 VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__o32a_1
X_10615_ cpuregs\[28\]\[7\] cpuregs\[29\]\[7\] net669 VGND VGND VPWR VPWR _05308_
+ sky130_fd_sc_hd__mux2_1
X_14383_ clknet_leaf_83_clk _00804_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dfxtp_2
X_11595_ mem_rdata_q\[30\] _06196_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ net708 _02225_ _02247_ _02249_ net391 VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__a311o_1
X_10546_ net772 _05232_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__and3_1
X_13265_ _02405_ net752 VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__nand2_1
XFILLER_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10477_ cpuregs\[1\]\[1\] net551 _05175_ net805 net832 VGND VGND VPWR VPWR _05176_
+ sky130_fd_sc_hd__a221o_1
X_15004_ clknet_leaf_145_clk _01356_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12216_ net748 _06600_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__nor2_1
X_13196_ net1981 net282 net430 VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12147_ net2833 net382 net371 net2909 VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__a22o_1
XFILLER_150_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12078_ net863 _06521_ _06522_ _06526_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__a31o_1
XANTENNA__12668__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07139__A1 _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11029_ net1075 decoded_imm\[18\] VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__or2_1
XANTENNA__11583__C net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07135__A net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10694__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13571__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10767__Y _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11643__A0 decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14719_ clknet_leaf_155_clk _01104_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08240_ net1170 net250 net941 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__mux2_1
XFILLER_166_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13396__B1 net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08171_ _03269_ _03662_ _03661_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__a21o_1
XANTENNA__12915__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10749__A2 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07122_ genblk2.pcpi_div.dividend\[27\] genblk2.pcpi_div.dividend\[26\] _02657_ _02677_
+ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__or4_1
XANTENNA__08253__X net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07053_ net1114 _02619_ genblk2.pcpi_div.dividend\[19\] VGND VGND VPWR VPWR _02620_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_93_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput100 net100 VGND VGND VPWR VPWR mem_la_wdata[12] sky130_fd_sc_hd__buf_2
XANTENNA__09509__B _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput111 net111 VGND VGND VPWR VPWR mem_la_wdata[22] sky130_fd_sc_hd__buf_2
Xoutput122 net1176 VGND VGND VPWR VPWR mem_la_wdata[3] sky130_fd_sc_hd__buf_2
Xoutput133 net133 VGND VGND VPWR VPWR mem_la_wstrb[3] sky130_fd_sc_hd__buf_2
XFILLER_115_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput144 net144 VGND VGND VPWR VPWR mem_wdata[18] sky130_fd_sc_hd__buf_2
XFILLER_114_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput155 net155 VGND VGND VPWR VPWR mem_wdata[28] sky130_fd_sc_hd__buf_2
Xoutput166 net166 VGND VGND VPWR VPWR mem_wdata[9] sky130_fd_sc_hd__buf_2
XFILLER_115_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput177 net177 VGND VGND VPWR VPWR pcpi_insn[15] sky130_fd_sc_hd__buf_2
XFILLER_99_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput188 net188 VGND VGND VPWR VPWR pcpi_insn[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput199 net199 VGND VGND VPWR VPWR pcpi_insn[6] sky130_fd_sc_hd__buf_2
XFILLER_130_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ net771 _03470_ _03471_ _03468_ VGND VGND VPWR VPWR alu_out\[1\] sky130_fd_sc_hd__a31o_1
XFILLER_130_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout381_A net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net483 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06906_ net2932 _02460_ _02467_ net1054 _02499_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__a221o_1
XFILLER_29_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07886_ net248 _02410_ _03403_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__o21ai_1
X_09625_ reg_pc\[18\] net877 _04439_ net847 VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__a22o_1
X_06837_ net1232 net2673 VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__and2_1
XFILLER_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13481__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07550__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09556_ count_instr\[52\] _04398_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__or2_1
X_06768_ net2561 VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__inv_2
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08507_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__inv_2
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09487_ count_instr\[27\] count_instr\[26\] _04352_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout434_X net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_X net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08438_ reg_pc\[24\] reg_pc\[23\] _03834_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__and3_1
X_08369_ reg_out\[11\] alu_out_q\[11\] net1153 VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout601_X net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12825__S net466 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10400_ net1164 _05104_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__or2_1
XFILLER_165_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11380_ net783 _06042_ _06051_ net778 VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__o211a_1
XFILLER_137_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10331_ _05035_ _05036_ _04891_ _05034_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__a211o_1
XANTENNA__09419__B net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12126__A net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10262_ _04944_ _04946_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__nor2_1
X_13050_ net1494 net73 net534 VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout970_X net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12001_ net1028 net723 _06459_ net862 VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__a31o_1
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11965__A net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10193_ decoded_imm\[26\] net1000 VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__nor2_1
XFILLER_132_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07654__S net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__buf_4
XFILLER_94_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13311__B1 net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout371 net372 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout382 net383 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_4
Xfanout393 _04888_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_4
X_13952_ clknet_leaf_2_clk _00406_ VGND VGND VPWR VPWR cpuregs\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_161_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12903_ net527 net2249 net455 VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13883_ clknet_leaf_196_clk _00337_ VGND VGND VPWR VPWR cpuregs\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07541__A1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15622_ clknet_leaf_36_clk _01958_ VGND VGND VPWR VPWR cpuregs\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12834_ net577 net2274 net459 VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__mux2_1
XANTENNA__06794__A net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14784__Q genblk2.pcpi_div.pcpi_rd\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15553_ clknet_leaf_50_clk _01889_ VGND VGND VPWR VPWR cpuregs\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12765_ net1215 genblk1.genblk1.pcpi_mul.next_rs1\[33\] net2501 net906 net762 VGND
+ VGND VPWR VPWR _01404_ sky130_fd_sc_hd__a221o_1
XFILLER_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14504_ clknet_leaf_91_clk _00893_ VGND VGND VPWR VPWR instr_rdinstr sky130_fd_sc_hd__dfxtp_2
XANTENNA__11205__A net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11716_ _06169_ _06226_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__nor2_1
XFILLER_15_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15484_ clknet_leaf_15_clk _01820_ VGND VGND VPWR VPWR cpuregs\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12696_ net1213 net2945 net901 net2963 net714 VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__a221o_1
XFILLER_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14435_ clknet_leaf_65_clk _00824_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dfxtp_1
X_11647_ decoded_imm_j\[12\] net4 net545 VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__mux2_1
Xinput13 mem_rdata[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
Xinput24 mem_rdata[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_167_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13451__A2_N _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14366_ clknet_leaf_170_clk _00787_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dfxtp_2
X_11578_ is_lb_lh_lw_lbu_lhu net747 VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__and2_1
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13317_ net556 _02211_ _02232_ _02234_ net391 VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__a311o_1
Xhold808 cpuregs\[26\]\[22\] VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold819 genblk1.genblk1.pcpi_mul.next_rs1\[12\] VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ net790 _05219_ _05221_ _05223_ net776 VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__o41a_1
XFILLER_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14297_ clknet_leaf_124_clk _00751_ VGND VGND VPWR VPWR count_cycle\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13248_ net1035 net758 _02173_ _02474_ net1064 VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__o2111a_1
XFILLER_124_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13566__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12470__S net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13179_ net1883 _03799_ net427 VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11594__B mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08309__A0 net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1508 genblk1.genblk1.pcpi_mul.pcpi_rd\[16\] VGND VGND VPWR VPWR net2822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_194_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1519 genblk2.pcpi_div.quotient_msk\[6\] VGND VGND VPWR VPWR net2833 sky130_fd_sc_hd__dlygate4sd3_1
X_07740_ cpuregs\[17\]\[4\] net641 net614 _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__o211a_1
XANTENNA__07136__Y _02690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10667__B2 net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07671_ _03191_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__inv_2
XANTENNA__10003__B net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09410_ net2558 _04302_ _04304_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__o21a_1
XANTENNA__08395__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09341_ net1790 net405 net476 VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09272_ net1703 net408 net485 VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__mux2_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13369__B1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08223_ net1058 net1176 net237 net1055 VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__a22o_1
XFILLER_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10954__A net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07048__B1 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13330__A net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08154_ _03590_ _03643_ _03647_ _03646_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__a31o_1
XFILLER_119_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11395__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07105_ net1123 genblk2.pcpi_div.quotient\[27\] _02661_ net952 VGND VGND VPWR VPWR
+ _02664_ sky130_fd_sc_hd__a31o_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08085_ _03345_ net932 net770 _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1136_A instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_147_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07036_ net1114 _02603_ genblk2.pcpi_div.dividend\[17\] VGND VGND VPWR VPWR _02605_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout596_A _03153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13476__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12344__B2 mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06879__A net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08987_ net1748 _04270_ net945 VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout384_X net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_102_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07938_ _03453_ _03454_ _03455_ _03392_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__a31o_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10658__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout551_X net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07869_ _03288_ _03301_ _03376_ _03379_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout930_A _03462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07523__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout649_X net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09608_ _03783_ reg_next_pc\[10\] net920 VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_104_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10880_ net240 net855 _05564_ _05565_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09539_ count_instr\[46\] _04387_ net1214 VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08079__A2 net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout816_X net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _02034_ net2631 net389 VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11501_ pcpi_timeout_counter\[1\] pcpi_timeout_counter\[0\] net2606 VGND VGND VPWR
+ VPWR _06162_ sky130_fd_sc_hd__o21a_1
XANTENNA__10830__A1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12481_ _06705_ _06706_ net2533 net386 VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__a2bb2o_1
X_14220_ clknet_leaf_67_clk _00674_ VGND VGND VPWR VPWR reg_pc\[28\] sky130_fd_sc_hd__dfxtp_1
X_11432_ net837 _06098_ _06100_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__a211o_1
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10043__C1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14151_ clknet_leaf_99_clk _00605_ VGND VGND VPWR VPWR count_instr\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11363_ net1081 _06034_ _06035_ net858 VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__a211o_1
XANTENNA__10594__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13102_ net575 net2405 net436 VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__mux2_1
X_10314_ _05003_ _05005_ _05019_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__or3_1
XFILLER_153_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14082_ clknet_leaf_18_clk _00536_ VGND VGND VPWR VPWR cpuregs\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11294_ cpuregs\[4\]\[26\] cpuregs\[5\]\[26\] net702 VGND VGND VPWR VPWR _05968_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11138__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12335__A1 decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08988__B net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12335__B2 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13033_ net282 net2342 net445 VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__mux2_1
XFILLER_112_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10245_ net1047 decoded_imm\[1\] VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_163_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06789__A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1100 net1109 VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__clkbuf_2
XFILLER_121_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14779__Q genblk2.pcpi_div.pcpi_rd\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1111 genblk2.pcpi_div.pcpi_ready VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10176_ net1207 _02478_ _04881_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__or3_1
Xfanout1122 net1123 VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__buf_2
Xfanout1133 net1134 VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__buf_2
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1144 net1145 VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__clkbuf_2
Xfanout1155 net1156 VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__buf_4
Xfanout1166 net236 VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__clkbuf_4
X_14984_ clknet_leaf_108_clk _01336_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1177 net119 VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__buf_4
Xfanout1188 net1189 VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1199 net1204 VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_141_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13935_ clknet_leaf_44_clk _00389_ VGND VGND VPWR VPWR cpuregs\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09503__A2 _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__A1 genblk2.pcpi_div.pcpi_rd\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11718__A_N net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13415__A net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkload5_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13866_ clknet_leaf_46_clk _00320_ VGND VGND VPWR VPWR cpuregs\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09104__S net505 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15605_ clknet_leaf_199_clk _01941_ VGND VGND VPWR VPWR cpuregs\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12817_ net327 net2307 net465 VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__mux2_1
XFILLER_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13797_ clknet_leaf_17_clk _00251_ VGND VGND VPWR VPWR cpuregs\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15536_ clknet_leaf_193_clk _01872_ VGND VGND VPWR VPWR cpuregs\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12748_ net1199 genblk1.genblk1.pcpi_mul.next_rs1\[23\] net916 net1005 VGND VGND
+ VPWR VPWR _02108_ sky130_fd_sc_hd__a22o_1
XANTENNA__08943__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15467_ clknet_leaf_29_clk _01803_ VGND VGND VPWR VPWR cpuregs\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ net1193 net2826 net886 net2938 net711 VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__a221o_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14418_ clknet_leaf_77_clk alu_out\[18\] VGND VGND VPWR VPWR alu_out_q\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13220__C1 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15398_ clknet_leaf_31_clk _01737_ VGND VGND VPWR VPWR cpuregs\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14349_ clknet_leaf_66_clk _06737_ VGND VGND VPWR VPWR reg_out\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold605 cpuregs\[4\]\[21\] VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 cpuregs\[20\]\[9\] VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09774__S net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold627 cpuregs\[25\]\[4\] VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold638 cpuregs\[15\]\[19\] VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 cpuregs\[25\]\[27\] VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12326__A1 decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08910_ _04068_ _04070_ _04067_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__a21bo_1
X_09890_ _04441_ _04646_ _04442_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_954 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08841_ _04173_ _04176_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__nand2_1
XFILLER_111_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1305 _06610_ VGND VGND VPWR VPWR net2619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1316 reg_next_pc\[2\] VGND VGND VPWR VPWR net2630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1327 genblk1.genblk1.pcpi_mul.rd\[56\] VGND VGND VPWR VPWR net2641 sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ net885 _04119_ _04121_ net2676 net1194 VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__a32o_1
XFILLER_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1338 genblk1.genblk1.pcpi_mul.rd\[50\] VGND VGND VPWR VPWR net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1349 genblk2.pcpi_div.running VGND VGND VPWR VPWR net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09803__A decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07723_ cpuregs\[9\]\[4\] net640 net614 _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__o211a_1
XFILLER_66_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07654_ _03173_ _03174_ net807 VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09014__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07887__A_N net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07585_ genblk1.genblk1.pcpi_mul.pcpi_rd\[29\] genblk2.pcpi_div.pcpi_rd\[29\] net1113
+ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1086_A net1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08138__B net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09324_ net1569 net299 net482 VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__mux2_1
XANTENNA__11065__A1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07269__B1 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12262__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpicorv32_1245 VGND VGND VPWR VPWR picorv32_1245/HI eoi[3] sky130_fd_sc_hd__conb_1
Xpicorv32_1256 VGND VGND VPWR VPWR picorv32_1256/HI eoi[14] sky130_fd_sc_hd__conb_1
Xpicorv32_1267 VGND VGND VPWR VPWR picorv32_1267/HI eoi[25] sky130_fd_sc_hd__conb_1
X_09255_ net1619 net302 net491 VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout511_A _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12375__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10812__B2 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1278 VGND VGND VPWR VPWR picorv32_1278/HI trace_data[0] sky130_fd_sc_hd__conb_1
XANTENNA_fanout609_A _03148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1289 VGND VGND VPWR VPWR picorv32_1289/HI trace_data[11] sky130_fd_sc_hd__conb_1
X_08206_ net966 _03367_ _03368_ net929 _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__a221o_1
XFILLER_147_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09186_ net315 net1987 net498 VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__mux2_1
X_08137_ _03465_ _03632_ _03625_ VGND VGND VPWR VPWR alu_out\[22\] sky130_fd_sc_hd__o21ai_2
XFILLER_162_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1041_X net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10040__A2 _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08068_ _03376_ _03569_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout880_A net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net979 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07019_ _02585_ _02586_ _02590_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__o21ai_1
XFILLER_150_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10030_ _04786_ _04787_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout766_X net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07744__A1 net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout933_X net933 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11981_ net1039 net1036 _06434_ net723 VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__o31a_1
XFILLER_57_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13720_ clknet_leaf_150_clk _00174_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10932_ cpuregs\[10\]\[16\] net655 VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__or2_1
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10500__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13651_ clknet_leaf_116_clk _00105_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_10863_ cpuregs\[24\]\[14\] net651 VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__or2_1
XFILLER_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12602_ net285 net2169 net469 VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__mux2_1
X_13582_ net289 net2484 net413 VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__mux2_1
XANTENNA__12253__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11056__B2 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10794_ cpuregs\[12\]\[12\] cpuregs\[13\]\[12\] net650 VGND VGND VPWR VPWR _05482_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15321_ clknet_leaf_14_clk _01661_ VGND VGND VPWR VPWR cpuregs\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_156_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10803__A1 net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12533_ genblk2.pcpi_div.divisor\[53\] _02021_ net872 VGND VGND VPWR VPWR _02022_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07887__B net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15252_ clknet_leaf_48_clk _01593_ VGND VGND VPWR VPWR cpuregs\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07680__B1 net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12464_ _05100_ net717 VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__nand2_1
XFILLER_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14203_ clknet_leaf_177_clk _00657_ VGND VGND VPWR VPWR reg_pc\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11359__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11415_ cpuregs\[11\]\[29\] net642 net602 _06085_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__o211a_1
X_15183_ clknet_leaf_32_clk _01532_ VGND VGND VPWR VPWR cpuregs\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08224__A2 net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12395_ net575 net2046 net472 VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14134_ clknet_leaf_127_clk _00588_ VGND VGND VPWR VPWR count_instr\[5\] sky130_fd_sc_hd__dfxtp_1
X_11346_ cpuregs\[30\]\[27\] cpuregs\[31\]\[27\] net694 VGND VGND VPWR VPWR _06019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07983__A1 net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12308__B2 mem_rdata_q\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14065_ clknet_leaf_179_clk _00519_ VGND VGND VPWR VPWR cpuregs\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11277_ cpuregs\[19\]\[25\] net642 net602 VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__o21a_1
X_13016_ net349 net2198 net443 VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__mux2_1
X_10228_ decoded_imm\[9\] net1031 VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__nor2_1
XANTENNA__07735__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10159_ _04869_ _04870_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__nor2_1
Xhold2 genblk1.genblk1.pcpi_mul.instr_mul VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08938__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14967_ clknet_leaf_151_clk _01319_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13284__A2 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13918_ clknet_leaf_18_clk _00372_ VGND VGND VPWR VPWR cpuregs\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_14898_ clknet_leaf_143_clk _01250_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_13849_ clknet_leaf_191_clk _00303_ VGND VGND VPWR VPWR cpuregs\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_138_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12244__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07370_ reg_pc\[14\] decoded_imm\[14\] _02895_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_44_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07797__B net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15519_ clknet_leaf_81_clk _01855_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dfxtp_1
XANTENNA__15292__CLK clknet_4_10_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09040_ net349 net2351 net512 VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__mux2_1
XFILLER_163_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12547__A1 net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08215__A2 _02384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12923__S net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold402 cpuregs\[10\]\[7\] VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 cpuregs\[4\]\[13\] VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 cpuregs\[4\]\[20\] VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 cpuregs\[22\]\[10\] VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08261__X net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold446 cpuregs\[8\]\[11\] VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 cpuregs\[15\]\[3\] VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 net173 VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09942_ _04445_ _04446_ _04691_ _04447_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__a31o_1
Xhold479 cpuregs\[7\]\[26\] VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 net905 VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__buf_2
XANTENNA__12224__A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09009__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout915 net919 VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__buf_2
Xfanout926 net927 VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout937 _02910_ VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__clkbuf_2
X_09873_ _04638_ _04644_ _04654_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__or3_1
Xfanout948 net949 VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07726__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_A _03857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout959 _02463_ VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__buf_4
XFILLER_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08824_ net896 _04163_ _04165_ net2610 net1203 VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__a32o_1
Xhold1102 cpuregs\[17\]\[1\] VGND VGND VPWR VPWR net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 cpuregs\[3\]\[19\] VGND VGND VPWR VPWR net2427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 cpuregs\[7\]\[27\] VGND VGND VPWR VPWR net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 cpuregs\[7\]\[17\] VGND VGND VPWR VPWR net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 cpuregs\[19\]\[1\] VGND VGND VPWR VPWR net2460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08755_ genblk1.genblk1.pcpi_mul.rd\[42\] genblk1.genblk1.pcpi_mul.next_rs2\[43\]
+ net1091 VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_68_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1157 cpuregs\[7\]\[23\] VGND VGND VPWR VPWR net2471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A _02118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1168 cpuregs\[1\]\[5\] VGND VGND VPWR VPWR net2482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1179 cpuregs\[18\]\[29\] VGND VGND VPWR VPWR net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11274__S net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07706_ net772 _03217_ _03225_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__and3_1
X_08686_ _04047_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12483__B1 net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_156_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ net835 _03146_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__a21o_1
XFILLER_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout726_A _06409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1089_X net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ count_instr\[60\] net1134 net1141 count_cycle\[60\] VGND VGND VPWR VPWR _03093_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06892__A net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09307_ net1357 _03782_ net480 VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout514_X net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07499_ net1067 net1006 _03028_ net1082 _03027_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__a221o_1
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09651__B2 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09238_ net1529 net520 net488 VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__mux2_1
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09169_ net541 net2224 net499 VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__mux2_1
XANTENNA__12833__S net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10549__B1 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11200_ cpuregs\[2\]\[23\] cpuregs\[3\]\[23\] net675 VGND VGND VPWR VPWR _05877_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_165_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09708__A decoded_imm_j\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07902__A_N net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12180_ net751 net2695 VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout883_X net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11131_ net824 _05805_ _05807_ _05809_ net788 VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_112_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold980 cpuregs\[11\]\[27\] VGND VGND VPWR VPWR net2294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold991 cpuregs\[18\]\[30\] VGND VGND VPWR VPWR net2305 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ cpuregs\[25\]\[19\] net632 net610 _05742_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__o211a_1
XANTENNA__15218__Q cpu_state\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12710__A1 net1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07717__B2 net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12710__B2 net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10013_ net2848 _04775_ net1223 VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07662__S net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input22_A mem_rdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14821_ clknet_leaf_82_clk _01173_ VGND VGND VPWR VPWR decoded_imm\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1680 instr_bgeu VGND VGND VPWR VPWR net2994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1691 instr_and VGND VGND VPWR VPWR net3005 sky130_fd_sc_hd__dlygate4sd3_1
X_14752_ clknet_leaf_152_clk _01137_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_ready
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_57_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11964_ net1043 _06423_ net726 VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__o21ai_1
X_13703_ clknet_leaf_147_clk _00157_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10915_ net1075 decoded_imm\[15\] VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__or2_1
X_14683_ clknet_leaf_153_clk _01068_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_11895_ _02359_ genblk2.pcpi_div.dividend\[20\] _06275_ VGND VGND VPWR VPWR _06366_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07350__C1 _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13634_ clknet_leaf_144_clk _00088_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10846_ cpuregs\[5\]\[14\] net623 net811 _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__o211a_1
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13565_ net355 net2301 net412 VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__mux2_1
X_10777_ cpuregs\[27\]\[12\] net619 net590 _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_136_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15304_ clknet_leaf_17_clk _01644_ VGND VGND VPWR VPWR cpuregs\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12516_ _02007_ _02008_ net2563 net385 VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_23_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13496_ net1943 net520 net420 VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__mux2_1
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15235_ clknet_leaf_20_clk _01576_ VGND VGND VPWR VPWR cpuregs\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12447_ _06680_ net2552 net383 VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__mux2_1
XANTENNA_output90_A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15166_ clknet_leaf_65_clk _01515_ VGND VGND VPWR VPWR mem_rdata_q\[17\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__11201__B2 net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12378_ net1342 net322 net361 VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__mux2_1
XFILLER_153_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14117_ clknet_leaf_37_clk _00571_ VGND VGND VPWR VPWR cpuregs\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07409__Y _02945_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11329_ cpuregs\[6\]\[27\] cpuregs\[7\]\[27\] net695 VGND VGND VPWR VPWR _06002_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11586__C mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12044__A net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15097_ clknet_leaf_6_clk _01449_ VGND VGND VPWR VPWR cpuregs\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14048_ clknet_leaf_1_clk _00502_ VGND VGND VPWR VPWR cpuregs\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13574__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06870_ net1152 net970 VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__or2_1
XANTENNA__10712__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08540_ genblk1.genblk1.pcpi_mul.rd\[9\] genblk1.genblk1.pcpi_mul.next_rs2\[10\]
+ net1091 VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__and3_1
XFILLER_82_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ net769 _03866_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__and2b_1
XFILLER_51_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12918__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10011__B net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07422_ _02953_ _02955_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__nand2_1
XFILLER_168_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07353_ reg_pc\[14\] decoded_imm\[14\] VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__xor2_1
XFILLER_149_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09633__B2 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07284_ net18 _02689_ _02694_ net32 _02812_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__o221a_1
X_09023_ net282 net2076 net518 VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__mux2_1
XANTENNA__11991__A2 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout307_A _03844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1049_A net1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold210 cpuregs\[12\]\[5\] VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold221 cpuregs\[12\]\[0\] VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 net147 VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold243 cpuregs\[28\]\[12\] VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold254 cpuregs\[21\]\[10\] VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _01397_ VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 cpuregs\[4\]\[29\] VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold287 cpuregs\[12\]\[4\] VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout701 net707 VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkbuf_4
Xhold298 cpuregs\[23\]\[23\] VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 _02083_ VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkbuf_2
X_09925_ net851 _04701_ _04702_ net881 net2910 VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__a32o_1
Xfanout723 _06409_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout734 net735 VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__buf_1
XANTENNA__13484__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout745 _06163_ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_A net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout756 net757 VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkbuf_4
Xfanout767 _03747_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__clkbuf_4
X_09856_ decoded_imm_j\[19\] _04440_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__nor2_1
XFILLER_112_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout778 _03169_ VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1004_X net1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout789 net791 VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07335__X _02876_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08807_ genblk1.genblk1.pcpi_mul.rd\[50\] genblk1.genblk1.pcpi_mul.next_rs2\[51\]
+ net1096 VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__nand3_1
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09787_ _02480_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__nand2_1
X_06999_ net1118 _02572_ net3025 VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout464_X net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12456__B1 net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08738_ _04091_ _04092_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__xnor2_1
X_08669_ genblk1.genblk1.pcpi_mul.next_rs2\[30\] net1106 genblk1.genblk1.pcpi_mul.rd\[29\]
+ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout631_X net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12828__S net466 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout729_X net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10700_ cpuregs\[4\]\[10\] cpuregs\[5\]\[10\] net666 VGND VGND VPWR VPWR _05390_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11680_ net2688 net737 net560 net2710 VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__a22o_1
XANTENNA__09202__S net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10631_ cpuregs\[1\]\[8\] net550 _05322_ net800 net827 VGND VGND VPWR VPWR _05323_
+ sky130_fd_sc_hd__a221o_1
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15501__Q net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13350_ net557 _02239_ _02263_ net565 reg_pc\[18\] VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__a32o_1
XANTENNA__11431__B2 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10562_ cpuregs\[8\]\[6\] net674 VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__or2_1
X_12301_ mem_rdata_q\[23\] net559 _06629_ net532 VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__a211o_1
XFILLER_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12563__S net390 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13281_ net1031 net753 net556 _02182_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_114_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10493_ cpuregs\[26\]\[1\] net691 VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__or2_1
XANTENNA__07650__A3 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15020_ clknet_leaf_122_clk net1492 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12232_ net750 _06608_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_131_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net2828 net378 net364 net2886 VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a22o_1
XFILLER_107_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08061__B net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11114_ _05790_ _05792_ net784 VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__a21o_1
X_12094_ _06267_ _06369_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__and2b_1
X_11045_ cpuregs\[9\]\[19\] net632 net610 _05725_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__o211a_1
XANTENNA__06797__A net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07166__A2 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input25_X net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output226_A net993 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14804_ clknet_leaf_77_clk _01156_ VGND VGND VPWR VPWR decoded_imm\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12996_ net1408 net292 net449 VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__mux2_1
X_14735_ clknet_leaf_164_clk _01120_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11947_ net873 _06323_ _06415_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_28_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11642__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13423__A net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14666_ clknet_leaf_152_clk _01051_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11878_ genblk2.pcpi_div.divisor\[14\] _02390_ _06348_ VGND VGND VPWR VPWR _06349_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__09112__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13617_ clknet_leaf_44_clk _00072_ VGND VGND VPWR VPWR cpuregs\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10829_ cpuregs\[27\]\[13\] net619 net590 _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__o211a_1
XFILLER_20_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14597_ clknet_leaf_115_clk _00983_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfxtp_1
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13411__A2 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13548_ net293 net2088 net417 VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__mux2_1
XANTENNA__08951__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13569__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13479_ net1742 net305 net426 VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__mux2_1
X_15218_ clknet_leaf_88_clk _00007_ VGND VGND VPWR VPWR cpu_state\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15149_ clknet_leaf_91_clk _01498_ VGND VGND VPWR VPWR mem_rdata_q\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10933__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07971_ net968 _03304_ net934 _03303_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__o22a_1
XFILLER_68_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09710_ _04494_ _04497_ _04493_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__o21a_1
XANTENNA__11489__A1 net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06922_ genblk2.pcpi_div.instr_rem net1370 _02509_ net1237 VGND VGND VPWR VPWR _00048_
+ sky130_fd_sc_hd__o31a_1
XFILLER_101_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08398__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12502__A net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09641_ reg_pc\[26\] net879 _04447_ net849 VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__a22o_1
X_06853_ instr_lhu instr_lw instr_lh VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_52_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09572_ count_instr\[57\] _04408_ _04410_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__o21a_1
X_06784_ net1176 VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__inv_2
XFILLER_83_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08523_ _03903_ _03906_ _03908_ _03909_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__o211a_1
XANTENNA__11110__B1 net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09854__A1 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08454_ reg_pc\[27\] reg_pc\[26\] _03847_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__and3_1
XANTENNA__11661__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09022__S net519 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07405_ _02939_ _02940_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__nand2_1
XFILLER_51_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08385_ net347 net2210 net528 VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__mux2_1
XFILLER_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout424_A net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1166_A net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10395__C net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08146__B net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07336_ net841 _02872_ _02873_ _02876_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__a31o_2
XANTENNA__13479__S net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12383__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07267_ _02367_ latched_is_lh net942 VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_59_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09006_ net349 net1488 net516 VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__mux2_1
XFILLER_152_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07198_ reg_pc\[4\] decoded_imm\[4\] VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout793_A net795 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10924__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09408__D net1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout960_A _02462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout520 net523 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkbuf_2
Xfanout531 _03746_ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout679_X net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout542 net544 VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09908_ _04442_ _04443_ net1127 VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__o21a_1
Xfanout553 _03156_ VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__buf_2
Xfanout564 net565 VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_2
Xfanout575 net576 VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12141__A2 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout586 net587 VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkbuf_2
Xfanout597 net600 VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkbuf_4
X_09839_ _04438_ _04611_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__or2_1
XFILLER_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout846_X net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12850_ net325 net2357 net461 VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__mux2_1
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11801_ genblk2.pcpi_div.divisor\[22\] genblk2.pcpi_div.dividend\[22\] VGND VGND
+ VPWR VPWR _06272_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_107_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ net1220 genblk1.genblk1.pcpi_mul.next_rs1\[49\] net2264 net909 net765 VGND
+ VGND VPWR VPWR _01420_ sky130_fd_sc_hd__a221o_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14520_ clknet_leaf_69_clk _00909_ VGND VGND VPWR VPWR decoded_rd\[0\] sky130_fd_sc_hd__dfxtp_1
X_11732_ latched_rd\[3\] _06242_ _06243_ net1613 VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__a22o_1
XANTENNA__10455__A2 net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11652__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14451_ clknet_4_11_0_clk _00840_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dfxtp_1
X_11663_ decoded_imm_j\[2\] net15 net546 VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13402_ _02501_ _02284_ _02307_ _02309_ net394 VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__a311o_1
XANTENNA__07608__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10614_ cpuregs\[30\]\[7\] cpuregs\[31\]\[7\] net669 VGND VGND VPWR VPWR _05307_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09867__S net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11404__A1 net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14382_ clknet_leaf_83_clk _00803_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dfxtp_2
XFILLER_167_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11594_ mem_rdata_q\[31\] mem_rdata_q\[29\] _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__or3_2
XFILLER_128_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13333_ net557 _02223_ _02248_ net564 reg_pc\[16\] VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__a32o_1
XANTENNA__07895__B net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10545_ net829 _05235_ _05237_ _05239_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__a211o_1
XFILLER_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_130_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_130_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13264_ net567 _05351_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__nor2_1
XFILLER_155_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10476_ cpuregs\[2\]\[1\] cpuregs\[3\]\[1\] net688 VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__mux2_1
X_15003_ clknet_leaf_146_clk net2929 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_12215_ net2810 net273 net2881 VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13195_ net1936 net287 net429 VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__mux2_1
X_12146_ net2529 net382 net371 net2833 VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ _06524_ _06525_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__nor2_1
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07139__A2 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09107__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12132__A2 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11028_ net772 _05701_ _05709_ _05693_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__a31oi_4
Xclkbuf_leaf_197_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_197_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07135__B net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08946__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12979_ net1563 net354 net448 VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__mux2_1
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14718_ clknet_leaf_156_clk _01103_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11643__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14649_ clknet_leaf_158_clk _01034_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12199__A2 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08170_ net252 net1002 _03292_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__a21o_1
XFILLER_119_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07121_ genblk2.pcpi_div.dividend\[29\] genblk2.pcpi_div.dividend\[28\] VGND VGND
+ VPWR VPWR _02677_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_121_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_121_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13148__A1 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07052_ genblk2.pcpi_div.dividend\[18\] genblk2.pcpi_div.dividend\[17\] _02603_ VGND
+ VGND VPWR VPWR _02619_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_93_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput101 net101 VGND VGND VPWR VPWR mem_la_wdata[13] sky130_fd_sc_hd__buf_2
XFILLER_161_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput112 net112 VGND VGND VPWR VPWR mem_la_wdata[23] sky130_fd_sc_hd__buf_2
Xoutput123 net1174 VGND VGND VPWR VPWR mem_la_wdata[4] sky130_fd_sc_hd__buf_2
Xoutput134 net134 VGND VGND VPWR VPWR mem_valid sky130_fd_sc_hd__buf_2
Xoutput145 net145 VGND VGND VPWR VPWR mem_wdata[19] sky130_fd_sc_hd__buf_2
XFILLER_114_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput156 net156 VGND VGND VPWR VPWR mem_wdata[29] sky130_fd_sc_hd__buf_2
Xoutput167 net167 VGND VGND VPWR VPWR mem_wstrb[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput178 net178 VGND VGND VPWR VPWR pcpi_insn[16] sky130_fd_sc_hd__buf_2
Xoutput189 net189 VGND VGND VPWR VPWR pcpi_insn[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13328__A _04987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12659__B1 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07954_ net1144 _02377_ _03469_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__or3_1
XANTENNA__12232__A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09017__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06905_ instr_lhu instr_lh net410 VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__o21a_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_188_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_188_clk sky130_fd_sc_hd__clkbuf_8
X_07885_ _03334_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__nand2_1
XFILLER_29_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout374_A net376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09624_ _03816_ reg_next_pc\[18\] net922 VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__mux2_2
X_06836_ _02440_ _02439_ net1232 VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__and3b_1
XFILLER_44_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09555_ _04398_ _04399_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__nor2_1
X_06767_ net2615 VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__inv_2
XANTENNA__12378__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11282__S net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_941 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08506_ genblk1.genblk1.pcpi_mul.rd\[4\] genblk1.genblk1.pcpi_mul.rdx\[4\] VGND VGND
+ VPWR VPWR _03896_ sky130_fd_sc_hd__nand2_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09486_ _04354_ _04355_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__nor2_1
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08437_ reg_pc\[23\] _03834_ reg_pc\[24\] VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1071_X net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A _03143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1169_X net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08368_ net405 net2156 net529 VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__mux2_1
XFILLER_20_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08263__A0 net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07319_ _02792_ _02795_ _02808_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__a211o_1
X_08299_ net1000 _03733_ net982 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_112_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_165_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10330_ net1188 decoded_imm\[31\] VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__nand2_1
XFILLER_125_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12126__B net995 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout796_X net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12841__S net460 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10261_ _04945_ _04947_ _04966_ _04946_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__a211o_1
XFILLER_106_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12000_ net723 _06459_ net1028 VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_148_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10192_ decoded_imm\[26\] net1000 VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__and2_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout350 net351 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_2
Xfanout361 net363 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09515__B1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout372 _06578_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13951_ clknet_leaf_2_clk _00405_ VGND VGND VPWR VPWR cpuregs\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xfanout383 net384 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_179_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_179_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout394 _04888_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11322__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12902_ net538 net2038 net455 VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10676__A2 net628 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13882_ clknet_leaf_196_clk _00336_ VGND VGND VPWR VPWR cpuregs\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15621_ clknet_leaf_49_clk _01957_ VGND VGND VPWR VPWR cpuregs\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12833_ net581 net2203 net462 VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__mux2_1
XFILLER_28_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ net1215 net2337 net2521 net906 net762 VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__a221o_1
X_15552_ clknet_leaf_57_clk _01888_ VGND VGND VPWR VPWR cpuregs\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14503_ clknet_leaf_91_clk _00892_ VGND VGND VPWR VPWR instr_rdcycleh sky130_fd_sc_hd__dfxtp_2
X_11715_ net2118 net280 net376 VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__mux2_1
XFILLER_159_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15483_ clknet_leaf_12_clk _01819_ VGND VGND VPWR VPWR cpuregs\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12695_ net1213 genblk1.genblk1.pcpi_mul.next_rs2\[60\] net901 net2958 net714 VGND
+ VGND VPWR VPWR _01365_ sky130_fd_sc_hd__a221o_1
XFILLER_159_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14434_ clknet_leaf_91_clk _00823_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11646_ decoded_imm_j\[10\] net24 net545 VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__mux2_1
Xinput14 mem_rdata[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_128_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 mem_rdata[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
X_14365_ clknet_leaf_171_clk _00786_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_103_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_8
X_11577_ net2904 net740 _06190_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__a22o_1
XFILLER_156_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13316_ net708 _02210_ _02233_ net564 reg_pc\[14\] VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__a32o_1
X_10528_ cpuregs\[11\]\[5\] net630 net595 _05222_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__o211a_1
Xhold809 cpuregs\[4\]\[11\] VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08006__S net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14296_ clknet_leaf_123_clk _00750_ VGND VGND VPWR VPWR count_cycle\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12889__A0 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13247_ net1040 net752 VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__or2_1
XFILLER_108_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10459_ cpuregs\[28\]\[0\] cpuregs\[29\]\[0\] net684 VGND VGND VPWR VPWR _05159_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13178_ net1806 net351 net427 VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__mux2_1
XANTENNA__11367__S net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12129_ _06260_ _06386_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__and2_1
XFILLER_2_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12052__A net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1509 genblk1.genblk1.pcpi_mul.next_rs2\[21\] VGND VGND VPWR VPWR net2823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13302__A1 decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11313__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13582__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10667__A2 net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07670_ _02475_ _02476_ net1066 VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09340_ net1798 _03782_ net475 VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__mux2_1
XANTENNA__12813__A0 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09271_ net2012 net520 net484 VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__mux2_1
XANTENNA__07296__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12926__S net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07296__B2 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08222_ net1056 net1177 net236 net942 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__a22o_1
XANTENNA__13369__B2 net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06924__S _02509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09300__S net482 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13330__B _05637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08153_ _03608_ _03626_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__nor2_1
XANTENNA__12041__B2 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07104_ net1122 _02661_ net2854 VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__a21oi_1
X_08084_ _03347_ _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07035_ genblk2.pcpi_div.dividend\[17\] net1114 _02603_ VGND VGND VPWR VPWR _02604_
+ sky130_fd_sc_hd__and3_1
XFILLER_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1129_A decoded_imm_j\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12344__A2 decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout491_A _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06879__B _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08986_ genblk1.genblk1.pcpi_mul.rd\[31\] genblk1.genblk1.pcpi_mul.rd\[63\] net957
+ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__mux2_1
X_07937_ instr_bne _03389_ _03452_ is_slti_blt_slt _03391_ VGND VGND VPWR VPWR _03455_
+ sky130_fd_sc_hd__a221oi_1
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11304__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout756_A net757 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_X net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13492__S net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07868_ _03285_ _03306_ _03383_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__or4_1
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06819_ instr_xori instr_addi instr_blt instr_bne VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__or4_1
X_09607_ reg_pc\[9\] net876 _04430_ net845 VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__a22o_1
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07799_ net1169 net1036 VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__nor2_1
XFILLER_73_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout923_A net927 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09538_ _04387_ _04388_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__nor2_1
XANTENNA__10210__A decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09469_ count_instr\[21\] count_instr\[20\] count_instr\[19\] _04338_ VGND VGND VPWR
+ VPWR _04344_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout711_X net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11083__A2 net624 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12836__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11740__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout809_X net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ net2861 net2850 _06157_ _06161_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__a211o_1
XFILLER_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12480_ net870 _06703_ _06704_ net386 VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__a31o_1
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09210__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11431_ cpuregs\[18\]\[29\] net555 _06101_ net786 VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__o22a_1
XANTENNA__08236__A0 net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14150_ clknet_leaf_97_clk _00604_ VGND VGND VPWR VPWR count_instr\[21\] sky130_fd_sc_hd__dfxtp_1
X_11362_ net1081 decoded_imm\[27\] VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nor2_1
XFILLER_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13101_ net579 net2461 net437 VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__mux2_1
X_10313_ _05007_ _05016_ _05018_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__or3b_1
XANTENNA__12571__S net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ clknet_leaf_41_clk _00535_ VGND VGND VPWR VPWR cpuregs\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11293_ cpuregs\[6\]\[26\] cpuregs\[7\]\[26\] net702 VGND VGND VPWR VPWR _05967_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13032_ net287 net2313 net446 VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__mux2_1
XANTENNA__12335__A2 net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10244_ net1047 decoded_imm\[1\] VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__and2_1
XFILLER_152_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10346__A1 net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_163_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1101 net1102 VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__buf_2
Xfanout1112 genblk2.pcpi_div.pcpi_ready VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__buf_4
X_10175_ net1088 _04880_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__nor2_1
Xfanout1123 net1124 VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__buf_2
Xfanout1134 instr_rdinstrh VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__buf_2
XFILLER_78_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1145 instr_sub VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__clkbuf_4
XFILLER_113_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1156 latched_stalu VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12099__A1 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1167 net266 VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__clkbuf_4
X_14983_ clknet_leaf_108_clk _01335_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1178 net1179 VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__buf_4
Xfanout1189 net227 VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__buf_4
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13934_ clknet_leaf_39_clk _00388_ VGND VGND VPWR VPWR cpuregs\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07253__X _02799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13415__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13865_ clknet_leaf_48_clk _00319_ VGND VGND VPWR VPWR cpuregs\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15604_ clknet_leaf_197_clk _01940_ VGND VGND VPWR VPWR cpuregs\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12816_ net331 net1872 net463 VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__mux2_1
XFILLER_90_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13796_ clknet_leaf_44_clk _00250_ VGND VGND VPWR VPWR cpuregs\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15535_ clknet_leaf_181_clk _01871_ VGND VGND VPWR VPWR cpuregs\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__06901__B_N is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12747_ net1191 net1328 net2392 net897 _02107_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__a221o_1
XFILLER_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11650__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10821__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12678_ net1193 net2938 net886 net2975 net711 VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__a221o_1
X_15466_ clknet_leaf_18_clk _01802_ VGND VGND VPWR VPWR cpuregs\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_139_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10774__B net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09120__S net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11629_ mem_rdata_q\[23\] mem_rdata_q\[22\] mem_rdata_q\[20\] mem_rdata_q\[21\] VGND
+ VGND VPWR VPWR _06216_ sky130_fd_sc_hd__or4b_1
XANTENNA__08227__B1 net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14417_ clknet_leaf_26_clk alu_out\[17\] VGND VGND VPWR VPWR alu_out_q\[17\] sky130_fd_sc_hd__dfxtp_1
X_15397_ clknet_leaf_45_clk _01736_ VGND VGND VPWR VPWR cpuregs\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14348_ clknet_leaf_68_clk _06736_ VGND VGND VPWR VPWR reg_out\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold606 cpuregs\[25\]\[10\] VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 cpuregs\[24\]\[23\] VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13577__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold628 cpuregs\[4\]\[5\] VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ clknet_leaf_98_clk _00733_ VGND VGND VPWR VPWR count_cycle\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold639 cpuregs\[10\]\[2\] VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10990__D1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09727__B1 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12326__A2 net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11534__A0 mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08840_ _04177_ _04178_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nand2_1
XFILLER_112_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14412__D alu_out\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10742__D1 net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1306 cpuregs\[16\]\[29\] VGND VGND VPWR VPWR net2620 sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__inv_2
Xhold1317 genblk2.pcpi_div.divisor\[56\] VGND VGND VPWR VPWR net2631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1328 reg_next_pc\[14\] VGND VGND VPWR VPWR net2642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1339 genblk2.pcpi_div.divisor\[51\] VGND VGND VPWR VPWR net2653 sky130_fd_sc_hd__dlygate4sd3_1
X_07722_ cpuregs\[8\]\[4\] net697 VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_69_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08259__X net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07653_ cpuregs\[22\]\[2\] cpuregs\[23\]\[2\] net701 VGND VGND VPWR VPWR _03174_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07584_ count_cycle\[29\] net973 net843 _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09323_ net1410 net303 net482 VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__mux2_1
XFILLER_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout337_A _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1246 VGND VGND VPWR VPWR picorv32_1246/HI eoi[4] sky130_fd_sc_hd__conb_1
XANTENNA_fanout1079_A cpu_state\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09254_ net1660 _03844_ net491 VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1257 VGND VGND VPWR VPWR picorv32_1257/HI eoi[15] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_32_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10812__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1268 VGND VGND VPWR VPWR picorv32_1268/HI eoi[26] sky130_fd_sc_hd__conb_1
Xpicorv32_1279 VGND VGND VPWR VPWR picorv32_1279/HI trace_data[1] sky130_fd_sc_hd__conb_1
XANTENNA__09030__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08205_ _03366_ net935 VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__nor2_1
XFILLER_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12014__A1 net1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08218__B1 net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09185_ net317 net2112 net497 VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout504_A _04279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08136_ _03323_ _03631_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07441__A1 net1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08067_ _03376_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__or2_1
XFILLER_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout1034_X net1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07485__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07018_ _02588_ _02589_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__or2_1
XANTENNA__11525__A0 mem_rdata_q\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10879__A2 _05563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08969_ net1731 _04261_ net945 VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__mux2_1
XANTENNA__06952__B1 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_X net759 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11735__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11980_ genblk2.pcpi_div.dividend\[7\] _06443_ net271 VGND VGND VPWR VPWR _01016_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10931_ cpuregs\[9\]\[16\] net621 net605 _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout926_X net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15504__Q net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__15731__A net1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10862_ _05546_ _05547_ net813 VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__mux2_1
X_13650_ clknet_leaf_116_clk _00104_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12601_ net291 net2503 net469 VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__mux2_1
X_13581_ net293 net2372 net413 VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__mux2_1
XFILLER_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11056__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12566__S net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10793_ cpuregs\[14\]\[12\] cpuregs\[15\]\[12\] net652 VGND VGND VPWR VPWR _05481_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15320_ clknet_leaf_40_clk _01660_ VGND VGND VPWR VPWR cpuregs\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12532_ net248 _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_193_clk_A clknet_4_0_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12463_ _06692_ net2546 net383 VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__mux2_1
X_15251_ clknet_leaf_34_clk _01592_ VGND VGND VPWR VPWR cpuregs\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13202__B1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11414_ cpuregs\[10\]\[29\] net702 VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__or2_1
XANTENNA__12556__A2 net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14202_ clknet_leaf_177_clk _00656_ VGND VGND VPWR VPWR reg_pc\[10\] sky130_fd_sc_hd__dfxtp_2
X_15182_ clknet_leaf_35_clk _01531_ VGND VGND VPWR VPWR cpuregs\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_117_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12394_ net579 net1828 net473 VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14133_ clknet_leaf_127_clk _00587_ VGND VGND VPWR VPWR count_instr\[4\] sky130_fd_sc_hd__dfxtp_1
X_11345_ cpuregs\[28\]\[27\] cpuregs\[29\]\[27\] net694 VGND VGND VPWR VPWR _06018_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13505__A1 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14064_ clknet_leaf_76_clk _00518_ VGND VGND VPWR VPWR cpuregs\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11516__A0 mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11276_ cpuregs\[17\]\[25\] net642 net615 _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__o211a_1
XFILLER_141_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output256_A net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13015_ net352 net2269 net443 VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__mux2_1
X_10227_ _04931_ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10158_ count_cycle\[58\] _04868_ net1239 VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13269__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 cpuregs\[0\]\[25\] VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11645__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10089_ _04825_ net1228 _04824_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__and3b_1
X_14966_ clknet_leaf_149_clk _01318_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09115__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13917_ clknet_leaf_7_clk _00371_ VGND VGND VPWR VPWR cpuregs\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07499__A1 net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07499__B2 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14897_ clknet_leaf_143_clk _01249_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08160__A2 net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_146_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13848_ clknet_leaf_188_clk _00302_ VGND VGND VPWR VPWR cpuregs\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08954__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11047__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13779_ clknet_leaf_22_clk _00233_ VGND VGND VPWR VPWR cpuregs\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15518_ clknet_leaf_79_clk _01854_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
X_15449_ clknet_leaf_15_clk _01788_ VGND VGND VPWR VPWR cpuregs\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10007__B1 net1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold403 cpuregs\[4\]\[6\] VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 cpuregs\[20\]\[11\] VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold425 cpuregs\[30\]\[7\] VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 cpuregs\[31\]\[5\] VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 net155 VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13100__S net438 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold458 cpuregs\[29\]\[28\] VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 cpuregs\[2\]\[19\] VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _04715_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout905 _03879_ VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout916 net919 VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__clkbuf_4
Xfanout927 _03708_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__clkbuf_4
X_09872_ _04651_ _04653_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__and2_1
XANTENNA__07187__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout938 net939 VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__buf_2
Xfanout949 _02509_ VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1103 cpuregs\[17\]\[5\] VGND VGND VPWR VPWR net2417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08823_ _04164_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__inv_2
Xhold1114 cpuregs\[13\]\[19\] VGND VGND VPWR VPWR net2428 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10730__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1125 cpuregs\[17\]\[6\] VGND VGND VPWR VPWR net2439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 cpuregs\[18\]\[19\] VGND VGND VPWR VPWR net2450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08754_ genblk1.genblk1.pcpi_mul.next_rs2\[43\] net1091 genblk1.genblk1.pcpi_mul.rd\[42\]
+ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__a21o_1
Xhold1147 cpuregs\[11\]\[2\] VGND VGND VPWR VPWR net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 genblk1.genblk1.pcpi_mul.next_rs1\[36\] VGND VGND VPWR VPWR net2472 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1169 genblk1.genblk1.pcpi_mul.pcpi_rd\[18\] VGND VGND VPWR VPWR net2483 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ net829 _03220_ _03222_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__a211o_1
XANTENNA__11286__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08685_ _04041_ _04044_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_92_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1196_A net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07636_ _03149_ net785 _03155_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__or3_1
XANTENNA__10494__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12386__S net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07567_ net21 net939 net937 VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_81_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11038__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13432__B1 net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09306_ net1530 net522 net480 VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout719_A net720 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07498_ genblk1.genblk1.pcpi_mul.pcpi_rd\[23\] genblk2.pcpi_div.pcpi_rd\[23\] net1112
+ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__mux2_1
XANTENNA__09651__A2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09237_ net1958 net524 net488 VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout507_X net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09168_ net571 net2341 net496 VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__mux2_1
XANTENNA__10549__A1 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout990_A _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07414__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08119_ _03615_ _03616_ _03607_ VGND VGND VPWR VPWR alu_out\[20\] sky130_fd_sc_hd__a21o_1
XFILLER_108_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11210__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10634__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09099_ net1650 net543 net507 VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07414__B2 net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13010__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11130_ cpuregs\[27\]\[21\] net632 net591 _05808_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__o211a_1
XFILLER_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold970 cpuregs\[9\]\[19\] VGND VGND VPWR VPWR net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 cpuregs\[19\]\[30\] VGND VGND VPWR VPWR net2295 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold992 cpuregs\[19\]\[16\] VGND VGND VPWR VPWR net2306 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ cpuregs\[24\]\[19\] net681 VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__or2_1
XFILLER_135_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07717__A2 net551 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10012_ count_cycle\[4\] count_cycle\[5\] count_cycle\[6\] _04771_ VGND VGND VPWR
+ VPWR _04776_ sky130_fd_sc_hd__and4_1
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14820_ clknet_leaf_82_clk _01172_ VGND VGND VPWR VPWR decoded_imm\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input15_A mem_rdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1670 decoded_imm_j\[8\] VGND VGND VPWR VPWR net2984 sky130_fd_sc_hd__dlygate4sd3_1
X_14751_ clknet_leaf_153_clk net2174 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[30\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1681 genblk1.genblk1.pcpi_mul.rd\[51\] VGND VGND VPWR VPWR net2995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11277__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11963_ _06327_ _06428_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__xnor2_1
Xhold1692 genblk1.genblk1.pcpi_mul.next_rs2\[40\] VGND VGND VPWR VPWR net3006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11131__D1 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_83_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_158_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ clknet_leaf_119_clk _00156_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10485__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11682__C1 net1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10914_ _05572_ _05581_ _05598_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__a21oi_4
X_14682_ clknet_leaf_153_clk _01067_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11894_ _06271_ _06272_ _06270_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__o21ba_1
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10845_ cpuregs\[4\]\[14\] net660 VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__or2_1
X_13633_ clknet_leaf_119_clk _00087_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10776_ cpuregs\[26\]\[12\] net650 VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__or2_1
X_13564_ net405 net2192 net412 VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__mux2_1
XANTENNA__07102__B1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15303_ clknet_leaf_31_clk _01643_ VGND VGND VPWR VPWR cpuregs\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12515_ net870 _02005_ _02006_ net385 VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_23_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13495_ net1657 net526 net420 VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15234_ clknet_leaf_181_clk _01575_ VGND VGND VPWR VPWR cpuregs\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12446_ genblk2.pcpi_div.divisor\[34\] _06679_ net868 VGND VGND VPWR VPWR _06680_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15165_ clknet_leaf_65_clk _01514_ VGND VGND VPWR VPWR mem_rdata_q\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11201__A2 net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12377_ net1809 net325 net362 VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__mux2_1
XANTENNA_output83_A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11328_ net253 net857 _06000_ _06001_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__a22o_1
X_14116_ clknet_leaf_44_clk _00570_ VGND VGND VPWR VPWR cpuregs\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15096_ clknet_leaf_19_clk _01448_ VGND VGND VPWR VPWR cpuregs\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14047_ clknet_leaf_0_clk _00501_ VGND VGND VPWR VPWR cpuregs\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_11259_ cpuregs\[2\]\[25\] net699 VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__or2_1
XANTENNA__08949__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12060__A net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14949_ clknet_leaf_33_clk _01301_ VGND VGND VPWR VPWR cpuregs\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08470_ reg_pc\[30\] _03863_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__nand2_1
XFILLER_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07421_ _02953_ _02955_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__or2_1
X_07352_ _02890_ _02891_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__or2_1
XANTENNA__09633__A2 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11976__B1 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07283_ _02807_ _02809_ _02824_ _02826_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__a31o_1
X_09022_ net287 net1838 net519 VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__mux2_1
XFILLER_129_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10962__B net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold200 cpuregs\[20\]\[17\] VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold211 cpuregs\[23\]\[16\] VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 cpuregs\[29\]\[5\] VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold233 cpuregs\[26\]\[8\] VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 cpuregs\[16\]\[2\] VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 cpuregs\[24\]\[26\] VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 cpuregs\[28\]\[15\] VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold277 cpuregs\[22\]\[21\] VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 cpuregs\[22\]\[23\] VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 decoded_rd\[3\] VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net705 VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__clkbuf_4
X_09924_ net1184 _04445_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__or2_1
Xfanout713 _02083_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkbuf_4
Xfanout724 net725 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1111_A genblk2.pcpi_div.pcpi_ready VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1209_A _02378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout735 _06164_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__buf_2
XANTENNA__12153__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout746 net747 VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07616__X _03137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input7_A mem_rdata[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout757 _04885_ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__buf_2
X_09855_ decoded_imm_j\[19\] _04440_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__and2_1
Xfanout768 _03747_ VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__buf_4
XANTENNA_fanout571_A _03761_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10703__B2 net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout779 net782 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__buf_4
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout669_A net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08806_ genblk1.genblk1.pcpi_mul.next_rs2\[51\] net1096 genblk1.genblk1.pcpi_mul.rd\[50\]
+ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__a21o_1
X_06998_ genblk2.pcpi_div.dividend\[11\] _02569_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__or2_1
X_09786_ _04567_ _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__xor2_1
XANTENNA__07064__A net1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06922__A3 _02509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08737_ _04085_ _04088_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__nand2_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10202__B net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_A net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_X net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10467__B1 net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08668_ net904 _04031_ _04033_ net2577 net1217 VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__a32o_1
X_07619_ net1080 decoded_imm_j\[15\] _03138_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10629__S net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08599_ genblk1.genblk1.pcpi_mul.rd\[18\] genblk1.genblk1.pcpi_mul.next_rs2\[19\]
+ net1097 VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout624_X net624 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10219__B1 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13005__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10630_ cpuregs\[2\]\[8\] cpuregs\[3\]\[8\] net674 VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10561_ net815 _05252_ _05254_ net829 VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__o211a_1
XANTENNA__11431__A2 net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12844__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ decoded_imm\[23\] net733 VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__and2_1
XFILLER_167_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13280_ net567 _05421_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__nor2_1
X_10492_ cpuregs\[25\]\[1\] net636 net612 _05190_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout993_X net993 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231_ net2732 net274 net2985 VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_131_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11195__B2 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12162_ net2810 net378 net365 net2828 VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_15_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08060__A1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10942__B2 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11113_ cpuregs\[1\]\[21\] net549 _05791_ net804 net825 VGND VGND VPWR VPWR _05792_
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12093_ genblk2.pcpi_div.dividend\[24\] _06539_ net273 VGND VGND VPWR VPWR _01033_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12144__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11044_ cpuregs\[8\]\[19\] net680 VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__or2_1
XFILLER_89_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11352__D1 net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ clknet_leaf_77_clk _01155_ VGND VGND VPWR VPWR decoded_imm\[19\] sky130_fd_sc_hd__dfxtp_2
XANTENNA_input18_X net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12995_ net1672 net296 net450 VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_56_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_output219_A net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14734_ clknet_leaf_164_clk _01119_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_24_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11946_ _06317_ _06318_ _06319_ _06322_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__a211o_1
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13423__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14665_ clknet_leaf_152_clk net2757 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11877_ _06294_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__or2_1
X_13616_ clknet_leaf_13_clk _00071_ VGND VGND VPWR VPWR cpuregs\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_10828_ cpuregs\[26\]\[13\] net650 VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__or2_1
X_14596_ clknet_leaf_159_clk _00982_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11958__B1 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13547_ net297 net1686 net418 VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_158_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10759_ net800 _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__or2_1
XFILLER_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13478_ net1551 net308 net424 VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__mux2_1
X_15217_ clknet_leaf_86_clk _00006_ VGND VGND VPWR VPWR cpu_state\[2\] sky130_fd_sc_hd__dfxtp_1
X_12429_ net2709 _06666_ _06667_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__o21ai_1
XFILLER_127_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07149__A net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08051__A1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15148_ clknet_leaf_80_clk _06750_ VGND VGND VPWR VPWR reg_sh\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13585__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07970_ _03273_ net932 _03480_ _03484_ VGND VGND VPWR VPWR alu_out\[3\] sky130_fd_sc_hd__a211o_1
X_15079_ clknet_leaf_102_clk net1962 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_06921_ genblk2.pcpi_div.instr_div genblk2.pcpi_div.instr_divu VGND VGND VPWR VPWR
+ _02509_ sky130_fd_sc_hd__or2_2
XANTENNA__11489__A2 _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06852_ mem_do_rdata net1208 _02454_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__nor3_1
X_09640_ _03850_ reg_next_pc\[26\] net924 VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__mux2_2
XFILLER_83_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14420__D alu_out\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09571_ count_instr\[57\] _04408_ net1215 VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_06783_ genblk2.pcpi_div.dividend\[6\] VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__inv_2
XFILLER_71_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_47_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
X_08522_ _03908_ _03909_ _03903_ _03906_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__a211o_1
XANTENNA__10449__B1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08267__X net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09303__S net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08453_ reg_pc\[26\] _03847_ reg_pc\[27\] VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07404_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__or2_1
X_08384_ _03795_ _03798_ net766 VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_98_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07335_ net1071 _02867_ _02868_ _02875_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_98_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10973__A net791 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A _02357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1159_A net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07266_ latched_is_lb _02799_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__and2_2
X_09005_ net352 net1802 net516 VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__mux2_1
XFILLER_164_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07197_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__inv_2
XFILLER_145_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11177__A1 net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout786_A _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13495__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09790__A1 net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09790__B2 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__06898__A net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout510 _04278_ VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout521 net522 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout532 _06620_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__buf_2
X_09907_ _04684_ _04685_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__nor2_1
XANTENNA__12677__A1 net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout543 net544 VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout953_A _02508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout554 _03156_ VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__buf_4
Xfanout565 net566 VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkbuf_4
Xfanout576 _03756_ VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__buf_1
X_09838_ _04438_ _04611_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__nand2_1
Xfanout587 _03749_ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10213__A decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout598 net600 VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12839__S net460 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09769_ _04543_ _04549_ _04558_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_38_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout839_X net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11743__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11800_ genblk2.pcpi_div.dividend\[23\] genblk2.pcpi_div.divisor\[23\] VGND VGND
+ VPWR VPWR _06271_ sky130_fd_sc_hd__and2b_1
XFILLER_73_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ net1220 genblk1.genblk1.pcpi_mul.next_rs1\[48\] net2469 net908 net765 VGND
+ VGND VPWR VPWR _01419_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09213__S net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11731_ latched_rd\[2\] _06242_ _06243_ net1406 VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14450_ clknet_leaf_55_clk _00839_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dfxtp_1
XFILLER_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11662_ decoded_imm_j\[1\] net14 net546 VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__mux2_1
XFILLER_23_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13401_ net558 _02285_ _02308_ net566 reg_pc\[24\] VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__a32o_1
X_10613_ net827 _05301_ _05303_ _05305_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__a211o_1
X_11593_ mem_rdata_q\[28\] mem_rdata_q\[27\] mem_rdata_q\[26\] mem_rdata_q\[25\] VGND
+ VGND VPWR VPWR _06195_ sky130_fd_sc_hd__or4_1
X_14381_ clknet_leaf_128_clk _00802_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dfxtp_4
XANTENNA__12574__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13332_ net1020 net754 VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__or2_1
X_10544_ cpuregs\[18\]\[5\] net552 _05238_ net781 VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__o22a_1
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13263_ net959 _04973_ _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__and3_1
X_10475_ net806 _05171_ _05173_ net839 VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__a211o_1
XANTENNA__11168__A1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15002_ clknet_leaf_147_clk _01354_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12214_ net748 net2762 VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__nor2_1
X_13194_ net2246 net290 net430 VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__mux2_1
XFILLER_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12145_ genblk2.pcpi_div.quotient_msk\[4\] net382 net371 net2529 VGND VGND VPWR VPWR
+ _01046_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12076_ net1008 net724 _06523_ net863 VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__a31o_1
XANTENNA__12668__B2 genblk1.genblk1.pcpi_mul.next_rs2\[32\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11027_ net822 _05704_ _05706_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__a211o_1
XANTENNA__07544__B1 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_92_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11653__S net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12978_ net1622 net406 net448 VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_61_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09123__S net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14717_ clknet_leaf_156_clk _01102_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_11929_ _06393_ _06398_ _06399_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__nor3_1
XFILLER_60_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07151__B net975 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14648_ clknet_leaf_160_clk _01033_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08962__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14579_ clknet_leaf_69_clk _00965_ VGND VGND VPWR VPWR latched_rd\[0\] sky130_fd_sc_hd__dfxtp_2
X_07120_ _02675_ _02676_ _02674_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10603__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07051_ genblk2.pcpi_div.quotient\[19\] _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14415__D alu_out\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput102 net102 VGND VGND VPWR VPWR mem_la_wdata[14] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR mem_la_wdata[24] sky130_fd_sc_hd__buf_2
Xoutput124 net1173 VGND VGND VPWR VPWR mem_la_wdata[5] sky130_fd_sc_hd__buf_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput135 net135 VGND VGND VPWR VPWR mem_wdata[0] sky130_fd_sc_hd__buf_2
Xoutput146 net146 VGND VGND VPWR VPWR mem_wdata[1] sky130_fd_sc_hd__buf_2
Xoutput157 net157 VGND VGND VPWR VPWR mem_wdata[2] sky130_fd_sc_hd__buf_2
Xoutput168 net168 VGND VGND VPWR VPWR mem_wstrb[1] sky130_fd_sc_hd__buf_2
Xoutput179 net179 VGND VGND VPWR VPWR pcpi_insn[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12513__A net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07953_ net1143 _02377_ _03469_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11316__D1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12659__B2 net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06904_ _02496_ _02497_ _02498_ _02494_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_50_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07884_ net247 net1010 VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__and2b_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09623_ reg_pc\[17\] net877 _04438_ net847 VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__a22o_1
XFILLER_95_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06835_ instr_ecall_ebreak pcpi_timeout VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__nor2_1
XFILLER_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09554_ net2954 _04396_ net1230 VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__o21ai_1
X_06766_ net2582 VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__inv_2
XFILLER_71_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09033__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08505_ net1199 net2872 net894 _03895_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__a22o_1
X_09485_ net3066 _04352_ net1239 VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout534_A _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10842__B1 net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08436_ reg_out\[24\] alu_out_q\[24\] net1156 VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__mux2_1
XFILLER_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08367_ _03783_ _03784_ net766 VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__mux2_2
XANTENNA__12394__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10907__S net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout701_A net707 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_X net1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07318_ _02824_ _02835_ _02848_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__or3_1
XFILLER_164_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08298_ reg_out\[26\] reg_next_pc\[26\] net924 VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__mux2_1
XFILLER_165_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07249_ _02790_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__or2_1
XFILLER_164_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10208__A decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1231_X net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08015__A1 net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10260_ _04937_ _04939_ _04943_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__or3_1
XANTENNA__08460__X _03860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11738__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09763__A1 net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ decoded_imm\[27\] net998 VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__or2_1
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09208__S net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_X net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout340 _03807_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__buf_1
XFILLER_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout351 net353 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_2
Xfanout362 net363 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_8
XANTENNA__15734__A net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout373 net374 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__buf_4
X_13950_ clknet_leaf_11_clk _00404_ VGND VGND VPWR VPWR cpuregs\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout384 net390 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_2
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout395 net398 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12901_ net543 net2323 net456 VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__mux2_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13881_ clknet_leaf_191_clk _00335_ VGND VGND VPWR VPWR cpuregs\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10878__A net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ clknet_leaf_53_clk _01956_ VGND VGND VPWR VPWR cpuregs\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12832_ net584 net2460 net461 VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__mux2_1
X_15551_ clknet_leaf_58_clk _01887_ VGND VGND VPWR VPWR cpuregs\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12763_ net1216 genblk1.genblk1.pcpi_mul.next_rs1\[31\] net2337 net907 net762 VGND
+ VGND VPWR VPWR _01402_ sky130_fd_sc_hd__a221o_1
X_14502_ clknet_leaf_91_clk _00891_ VGND VGND VPWR VPWR instr_rdcycle sky130_fd_sc_hd__dfxtp_1
XFILLER_43_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11714_ net2096 net282 net376 VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__mux2_1
X_15482_ clknet_leaf_42_clk _01818_ VGND VGND VPWR VPWR cpuregs\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12694_ net1212 net2958 net901 net2969 net714 VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__a221o_1
XFILLER_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14433_ clknet_leaf_91_clk net2555 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dfxtp_1
X_11645_ decoded_imm_j\[9\] net22 net545 VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__mux2_1
XFILLER_30_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 mem_rdata[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14364_ clknet_leaf_136_clk _00785_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_2
Xinput26 mem_rdata[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11576_ net741 _06188_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__nor2_1
XFILLER_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13315_ net1014 net758 VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__or2_1
X_10527_ cpuregs\[10\]\[5\] net675 VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__or2_1
X_14295_ clknet_leaf_123_clk _00749_ VGND VGND VPWR VPWR count_cycle\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13246_ _04943_ _04962_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__xnor2_1
X_10458_ net834 _05153_ _05155_ _05157_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__a211o_1
XANTENNA__12889__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11648__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177_ net1566 net357 net427 VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__mux2_1
X_10389_ _05086_ _05088_ _05091_ _05093_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__or4_1
XFILLER_124_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09118__S net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12128_ net993 net725 _06567_ net864 VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__a31o_1
XANTENNA__13302__A2 net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12059_ net721 _06508_ net1011 VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__a21o_1
XANTENNA__08957__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11383__S net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11077__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10300__B net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09270_ net1948 net524 net484 VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09690__B1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08221_ net1056 net1177 net236 net1055 VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__a22o_1
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13103__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08152_ _03326_ _03644_ _03645_ _03643_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__a22o_1
XANTENNA__08245__A1 net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07103_ _02658_ _02659_ _02661_ _02662_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08083_ net1143 _03342_ _03581_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__o31a_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12942__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07034_ genblk2.pcpi_div.dividend\[16\] _02596_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__or2_1
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout1024_A net1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09028__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08985_ net1496 _04269_ net946 VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__mux2_1
XANTENNA__10760__C1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_A _04288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07936_ _02413_ _02365_ _03451_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__mux2_1
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12389__S net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net654 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07867_ _03275_ _03279_ _03384_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__or3_1
XANTENNA__06895__B is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11293__S net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09606_ _03778_ reg_next_pc\[9\] net927 VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__mux2_2
XANTENNA__13057__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06818_ instr_beq instr_jal instr_rdcycle instr_srai VGND VGND VPWR VPWR _02423_
+ sky130_fd_sc_hd__or4_1
XFILLER_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07798_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09537_ net2832 _04386_ net1227 VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__o21ai_1
XFILLER_25_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10210__B net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_A net919 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_X net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ _04342_ _04343_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__nor2_1
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09681__B1 _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08419_ net321 net2475 net528 VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout704_X net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09399_ net199 net189 net191 net188 VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__or4b_1
XFILLER_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13013__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08236__A1 net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11430_ cpuregs\[19\]\[29\] net644 net602 VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__o21a_1
XFILLER_138_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10043__A1 _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11361_ net774 _06025_ _06033_ _06017_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__a31oi_4
XANTENNA__11240__B1 net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12852__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15729__A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10594__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10312_ _04911_ _04912_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__nor2_1
X_13100_ net584 net2507 net438 VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__mux2_1
XFILLER_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08190__X alu_out\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14080_ clknet_leaf_2_clk _00534_ VGND VGND VPWR VPWR cpuregs\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11292_ net252 net858 _05965_ _05966_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__a22o_1
XFILLER_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13031_ net289 net2273 net446 VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__mux2_1
X_10243_ decoded_imm\[2\] net1045 VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__nand2_1
XANTENNA__10372__S _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12740__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10174_ net1068 net958 VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__or2_1
Xfanout1102 net1104 VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__buf_2
Xfanout1113 genblk2.pcpi_div.pcpi_ready VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__buf_2
Xfanout1124 net1125 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1135 net1136 VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__buf_2
Xfanout1146 net1147 VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__buf_2
X_14982_ clknet_leaf_108_clk _01334_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1157 net259 VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__clkbuf_4
Xfanout1168 net265 VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__buf_4
XFILLER_93_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1179 net108 VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__buf_4
XFILLER_87_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13933_ clknet_leaf_49_clk _00387_ VGND VGND VPWR VPWR cpuregs\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13864_ clknet_leaf_57_clk _00318_ VGND VGND VPWR VPWR cpuregs\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13048__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10401__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15603_ clknet_leaf_196_clk _01939_ VGND VGND VPWR VPWR cpuregs\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12815_ net335 net1971 net463 VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__mux2_1
X_13795_ clknet_leaf_16_clk _00249_ VGND VGND VPWR VPWR cpuregs\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15534_ clknet_leaf_182_clk _01870_ VGND VGND VPWR VPWR cpuregs\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12746_ _02411_ net911 VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__nor2_1
XFILLER_31_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15465_ clknet_leaf_31_clk _01801_ VGND VGND VPWR VPWR cpuregs\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_12677_ net1197 genblk1.genblk1.pcpi_mul.next_rs2\[42\] net887 net2942 net711 VGND
+ VGND VPWR VPWR _01347_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_139_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08227__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14416_ clknet_leaf_175_clk alu_out\[16\] VGND VGND VPWR VPWR alu_out_q\[16\] sky130_fd_sc_hd__dfxtp_1
X_11628_ instr_rdcycleh net738 _06214_ _06215_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__a22o_1
XANTENNA__08227__B2 net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15396_ clknet_leaf_37_clk _01735_ VGND VGND VPWR VPWR cpuregs\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14347_ clknet_leaf_67_clk _06735_ VGND VGND VPWR VPWR reg_out\[27\] sky130_fd_sc_hd__dfxtp_1
X_11559_ net747 _06180_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__and2_1
XFILLER_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold607 cpuregs\[2\]\[9\] VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 cpuregs\[29\]\[26\] VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 cpuregs\[15\]\[8\] VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14278_ clknet_leaf_98_clk _00732_ VGND VGND VPWR VPWR count_cycle\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09727__A1 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13229_ _02151_ _02153_ _02157_ net396 net1044 VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__o32a_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07157__A reg_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1307 genblk1.genblk1.pcpi_mul.rdx\[20\] VGND VGND VPWR VPWR net2621 sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ genblk1.genblk1.pcpi_mul.next_rs2\[45\] net1090 _04116_ _04118_ VGND VGND
+ VPWR VPWR _04120_ sky130_fd_sc_hd__and4_1
Xhold1318 genblk1.genblk1.pcpi_mul.rd\[18\] VGND VGND VPWR VPWR net2632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1329 net192 VGND VGND VPWR VPWR net2643 sky130_fd_sc_hd__dlygate4sd3_1
X_07721_ _03238_ _03239_ net819 VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__mux2_1
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13039__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07652_ cpuregs\[20\]\[2\] cpuregs\[21\]\[2\] net697 VGND VGND VPWR VPWR _03173_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07583_ net1141 count_cycle\[61\] net978 _03106_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__a211o_1
XANTENNA__13444__D1 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12937__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09322_ net1624 net307 net481 VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__mux2_1
XFILLER_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12262__A2 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08275__X net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09311__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07620__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11470__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpicorv32_1247 VGND VGND VPWR VPWR picorv32_1247/HI eoi[5] sky130_fd_sc_hd__conb_1
X_09253_ net1602 net308 net490 VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1258 VGND VGND VPWR VPWR picorv32_1258/HI eoi[16] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_32_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1269 VGND VGND VPWR VPWR picorv32_1269/HI eoi[27] sky130_fd_sc_hd__conb_1
XFILLER_22_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11142__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08204_ _03370_ net933 _03687_ _03691_ VGND VGND VPWR VPWR alu_out\[30\] sky130_fd_sc_hd__a211o_1
XANTENNA__08218__A1 net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09184_ net322 net2014 net497 VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__mux2_1
XANTENNA__12014__A2 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08218__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09415__B1 net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08135_ _03629_ _03630_ net1144 VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__mux2_1
XANTENNA__09966__B2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_A net1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07977__B1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08066_ _03567_ _03568_ net988 VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__mux2_1
XFILLER_150_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07017_ net1115 genblk2.pcpi_div.quotient\[14\] _02587_ net950 VGND VGND VPWR VPWR
+ _02589_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout699_A net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1027_X net1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10205__B net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10920__S net811 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08968_ genblk1.genblk1.pcpi_mul.rd\[22\] genblk1.genblk1.pcpi_mul.rd\[54\] net956
+ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__mux2_1
XFILLER_69_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07919_ _03376_ _03379_ _03436_ _03410_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__a31oi_4
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout654_X net654 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08899_ net1192 net2649 net885 _04226_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13008__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10930_ cpuregs\[8\]\[16\] net657 VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__or2_1
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10861_ cpuregs\[28\]\[14\] cpuregs\[29\]\[14\] net664 VGND VGND VPWR VPWR _05547_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12847__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_X net821 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_X net919 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11751__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12600_ net293 net2353 net469 VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__mux2_1
XFILLER_140_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13580_ net297 net2251 net414 VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__mux2_1
XANTENNA__12253__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10792_ net838 _05477_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__o21a_1
XFILLER_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09221__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11461__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12531_ _05112_ net719 VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__nand2_1
XFILLER_157_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15250_ clknet_leaf_32_clk _01591_ VGND VGND VPWR VPWR cpuregs\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12462_ genblk2.pcpi_div.divisor\[38\] _06691_ net869 VGND VGND VPWR VPWR _06692_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13202__A1 net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13202__B2 net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14201_ clknet_leaf_173_clk _00655_ VGND VGND VPWR VPWR reg_pc\[9\] sky130_fd_sc_hd__dfxtp_1
X_11413_ cpuregs\[9\]\[29\] net643 net615 _06083_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__o211a_1
XANTENNA__09957__B2 net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12582__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15181_ clknet_leaf_37_clk _01530_ VGND VGND VPWR VPWR cpuregs\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12393_ _03751_ net2063 net473 VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__mux2_1
XANTENNA__11764__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07968__B1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14132_ clknet_leaf_127_clk _00586_ VGND VGND VPWR VPWR count_instr\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11344_ net783 _06007_ _06016_ net778 VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__o211a_1
XFILLER_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14063_ clknet_leaf_44_clk _00517_ VGND VGND VPWR VPWR cpuregs\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11275_ cpuregs\[16\]\[25\] net705 VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__or2_1
XFILLER_134_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13014_ net356 net1984 net443 VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__mux2_1
X_10226_ decoded_imm\[10\] net1029 VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__or2_1
XANTENNA_output249_A net249 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10157_ count_cycle\[58\] _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13269__B2 net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold4 cpuregs\[0\]\[30\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08300__S net925 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10088_ count_cycle\[32\] count_cycle\[33\] _04821_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__and3_1
X_14965_ clknet_leaf_149_clk _01317_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12330__B decoded_imm_j\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13916_ clknet_leaf_19_clk _00370_ VGND VGND VPWR VPWR cpuregs\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07499__A2 net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14896_ clknet_leaf_140_clk _01248_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09893__B1 net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13847_ clknet_leaf_182_clk _00301_ VGND VGND VPWR VPWR cpuregs\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11661__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13442__A net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12244__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13778_ clknet_leaf_23_clk _00232_ VGND VGND VPWR VPWR cpuregs\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09131__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15517_ clknet_leaf_81_clk _01853_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dfxtp_1
XFILLER_31_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12729_ net1331 net883 _02098_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__a21o_1
XANTENNA__12058__A net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15448_ clknet_leaf_12_clk _01787_ VGND VGND VPWR VPWR cpuregs\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08970__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15379_ clknet_leaf_1_clk _01718_ VGND VGND VPWR VPWR cpuregs\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12952__A0 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold404 net142 VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 cpuregs\[2\]\[18\] VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold426 decoded_rd\[0\] VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 cpuregs\[29\]\[31\] VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 cpuregs\[25\]\[13\] VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold459 cpuregs\[21\]\[9\] VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14423__D alu_out\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09940_ _04705_ _04708_ _04706_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12704__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout906 net907 VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout917 net918 VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__buf_2
XFILLER_124_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09871_ net1128 _04441_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__or2_1
Xfanout928 _03463_ VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07187__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout939 _02693_ VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__buf_2
X_08822_ genblk1.genblk1.pcpi_mul.next_rs2\[53\] net1102 _04160_ _04162_ VGND VGND
+ VPWR VPWR _04164_ sky130_fd_sc_hd__and4_1
Xhold1104 cpuregs\[1\]\[27\] VGND VGND VPWR VPWR net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 cpuregs\[19\]\[22\] VGND VGND VPWR VPWR net2429 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09306__S net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1126 cpuregs\[18\]\[4\] VGND VGND VPWR VPWR net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 cpuregs\[11\]\[6\] VGND VGND VPWR VPWR net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net886 _04103_ _04105_ net2842 net1193 VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__a32o_1
Xhold1148 cpuregs\[9\]\[18\] VGND VGND VPWR VPWR net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _01406_ VGND VGND VPWR VPWR net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07704_ cpuregs\[18\]\[3\] net552 _03223_ net781 VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__o22a_1
X_08684_ _04045_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__nand2_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07635_ net623 net788 VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__nand2_4
XFILLER_26_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout447_A net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07566_ _03086_ _03089_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__nand2_1
XANTENNA__13432__A1 net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12235__A2 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09041__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09305_ net1349 net525 net480 VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__mux2_1
X_07497_ count_cycle\[23\] net973 net843 _03026_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout614_A net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09236_ net1637 net539 net488 VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__mux2_1
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13498__S net420 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout402_X net402 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09167_ net576 net2050 net496 VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__mux2_1
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11746__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10549__A2 _05242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08118_ _03330_ _03614_ net771 VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_151_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07414__A2 net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09098_ net1918 net574 net507 VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__mux2_1
XFILLER_163_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08049_ _03288_ _03553_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__or2_1
XFILLER_150_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold960 cpuregs\[19\]\[3\] VGND VGND VPWR VPWR net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 cpuregs\[2\]\[31\] VGND VGND VPWR VPWR net2285 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11060_ _05739_ _05740_ net816 VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__mux2_1
Xhold982 reg_next_pc\[20\] VGND VGND VPWR VPWR net2296 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold993 cpuregs\[6\]\[19\] VGND VGND VPWR VPWR net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout771_X net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11746__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10011_ _04775_ net1223 _04774_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09216__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1660 count_instr\[13\] VGND VGND VPWR VPWR net2974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1671 genblk2.pcpi_div.quotient\[29\] VGND VGND VPWR VPWR net2985 sky130_fd_sc_hd__dlygate4sd3_1
X_14750_ clknet_leaf_153_clk _01135_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1682 count_cycle\[24\] VGND VGND VPWR VPWR net2996 sky130_fd_sc_hd__dlygate4sd3_1
X_11962_ _06309_ _06311_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__nor2_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1693 genblk1.genblk1.pcpi_mul.next_rs2\[34\] VGND VGND VPWR VPWR net3007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09740__A net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13701_ clknet_leaf_112_clk _00155_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_10913_ net772 _05589_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_158_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ clknet_leaf_153_clk net2792 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12577__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _06274_ _06277_ _06278_ _06362_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__or4bb_1
XFILLER_72_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13632_ clknet_leaf_120_clk _00086_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10844_ cpuregs\[6\]\[14\] cpuregs\[7\]\[14\] net660 VGND VGND VPWR VPWR _05530_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13563_ net407 net2282 net412 VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__mux2_1
X_10775_ cpuregs\[25\]\[12\] net619 net604 _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ clknet_leaf_44_clk _01642_ VGND VGND VPWR VPWR cpuregs\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_136_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12514_ genblk2.pcpi_div.divisor\[49\] net870 VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13494_ net2188 net537 net420 VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__mux2_1
XFILLER_12_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15233_ clknet_leaf_180_clk _01574_ VGND VGND VPWR VPWR cpuregs\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12445_ net1177 _06678_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10825__S net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11737__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15164_ clknet_leaf_64_clk _01513_ VGND VGND VPWR VPWR mem_rdata_q\[15\] sky130_fd_sc_hd__dfxtp_2
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12376_ net1391 net328 net360 VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__mux2_1
XFILLER_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ clknet_leaf_13_clk _00569_ VGND VGND VPWR VPWR cpuregs\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11327_ net1083 _05999_ net857 VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__a21oi_1
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15095_ clknet_leaf_4_clk _01447_ VGND VGND VPWR VPWR cpuregs\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_97_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14046_ clknet_leaf_10_clk _00500_ VGND VGND VPWR VPWR cpuregs\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output76_A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09915__A net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12698__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11258_ cpuregs\[1\]\[25\] net642 net615 _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11656__S net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10209_ decoded_imm\[17\] net1017 VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__nand2_1
XFILLER_122_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11189_ cpuregs\[22\]\[23\] cpuregs\[23\]\[23\] net675 VGND VGND VPWR VPWR _05866_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08118__B1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14948_ clknet_leaf_72_clk _01300_ VGND VGND VPWR VPWR cpuregs\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08965__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14879_ clknet_leaf_35_clk _01231_ VGND VGND VPWR VPWR cpuregs\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11391__S net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07420_ _02942_ _02939_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_63_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12217__A2 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07892__A2 net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07351_ net1071 _02882_ _02883_ _02888_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__a31o_1
XANTENNA__15160__Q mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07282_ net1071 _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__nand2_1
XFILLER_136_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09021_ net289 net1662 net519 VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__mux2_1
XFILLER_163_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13111__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold201 cpuregs\[13\]\[18\] VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 cpuregs\[13\]\[2\] VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 cpuregs\[28\]\[0\] VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14504__Q instr_rdinstr VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold234 cpuregs\[22\]\[11\] VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 cpuregs\[14\]\[31\] VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12950__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold256 cpuregs\[2\]\[24\] VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold267 cpuregs\[14\]\[0\] VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 cpuregs\[29\]\[22\] VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ net985 _04697_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__o21ai_1
Xfanout703 net704 VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__buf_2
Xhold289 cpuregs\[31\]\[7\] VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 _02083_ VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12689__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout397_A net398 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout725 _06409_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_74_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13350__B1 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout736 net738 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13347__A net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout747 _06163_ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkbuf_2
X_09854_ net847 _04636_ _04637_ net877 net2420 VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__a32o_1
XFILLER_58_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout758 _04884_ VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__buf_2
XFILLER_113_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout769 _03747_ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1104_A net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09036__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10703__A2 net550 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08805_ net889 _04147_ _04149_ net2870 net1197 VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__a32o_1
X_09785_ _04571_ _04573_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__and2_1
XANTENNA__07580__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06997_ net948 _02570_ _02571_ _02568_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout564_A net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08109__B1 net933 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_192_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08736_ _04089_ _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__nand2_1
XANTENNA__11113__C1 net825 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11664__A0 decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08667_ _04032_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__inv_2
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12397__S net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_A net830 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07618_ net1080 decoded_imm_j\[15\] _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__o21a_1
XFILLER_121_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08598_ genblk1.genblk1.pcpi_mul.next_rs2\[19\] net1097 genblk1.genblk1.pcpi_mul.rd\[18\]
+ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__a21o_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07080__A net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10219__A1 decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11416__B1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10219__B2 decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07549_ _03058_ _03061_ _03073_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07096__B1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10560_ net801 _05253_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09219_ net1592 net314 net494 VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__mux2_1
XANTENNA__10645__S net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10491_ cpuregs\[24\]\[1\] net683 VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__or2_1
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13021__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12230_ net750 net2807 VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07399__A1 genblk2.pcpi_div.pcpi_rd\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout986_X net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11195__A2 net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12860__S net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12161_ net2794 net384 net365 net2810 VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_145_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10942__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11112_ cpuregs\[2\]\[21\] cpuregs\[3\]\[21\] net685 VGND VGND VPWR VPWR _05791_
+ sky130_fd_sc_hd__mux2_1
X_12092_ _06538_ _06537_ _06535_ net863 VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold790 cpuregs\[19\]\[29\] VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13257__A _02404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13341__B1 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11043_ net804 _05721_ _05723_ net831 VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__o211a_1
XFILLER_150_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07571__A1 genblk2.pcpi_div.pcpi_rd\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_14802_ clknet_leaf_75_clk _01154_ VGND VGND VPWR VPWR decoded_imm\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12994_ net2547 net300 net450 VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__mux2_1
Xhold1490 _01053_ VGND VGND VPWR VPWR net2804 sky130_fd_sc_hd__dlygate4sd3_1
X_14733_ clknet_leaf_163_clk net2678 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14451__CLK clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11945_ net1046 _02443_ net726 net866 VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__a31o_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11505__A _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14664_ clknet_leaf_152_clk _01049_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11876_ _06296_ _06297_ _06346_ _06295_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__a31o_1
XANTENNA__11407__B1 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13615_ clknet_leaf_11_clk _00070_ VGND VGND VPWR VPWR cpuregs\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_10827_ cpuregs\[25\]\[13\] net619 net604 _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__o211a_1
X_14595_ clknet_leaf_159_clk _00981_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07087__B1 net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13546_ net301 net1868 net418 VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__mux2_1
X_10758_ cpuregs\[12\]\[11\] cpuregs\[13\]\[11\] net651 VGND VGND VPWR VPWR _05447_
+ sky130_fd_sc_hd__mux2_1
XFILLER_146_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13477_ net1420 net312 net425 VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__mux2_1
X_10689_ _05378_ _05379_ net800 VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__mux2_1
XANTENNA__12907__A0 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15216_ clknet_leaf_87_clk _00005_ VGND VGND VPWR VPWR cpu_state\[1\] sky130_fd_sc_hd__dfxtp_1
X_12428_ net2709 _06666_ net917 VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__a21oi_1
X_15147_ clknet_leaf_80_clk _06749_ VGND VGND VPWR VPWR reg_sh\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07149__B _02387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12359_ net1636 net584 net362 VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__mux2_1
XFILLER_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15078_ clknet_leaf_102_clk _01430_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06920_ genblk2.pcpi_div.instr_div genblk2.pcpi_div.instr_divu VGND VGND VPWR VPWR
+ _02508_ sky130_fd_sc_hd__nor2_1
X_14029_ clknet_leaf_50_clk _00483_ VGND VGND VPWR VPWR cpuregs\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_06851_ net1061 _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09570_ _04408_ _04409_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__nor2_1
X_06782_ genblk2.pcpi_div.dividend\[14\] VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__inv_2
XFILLER_83_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08521_ genblk1.genblk1.pcpi_mul.rd\[6\] genblk1.genblk1.pcpi_mul.next_rs2\[7\] net1097
+ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__nand3_1
XANTENNA__10449__A1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11646__A0 decoded_imm_j\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11110__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13106__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08452_ reg_out\[27\] alu_out_q\[27\] net1155 VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__mux2_1
XFILLER_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07403_ reg_pc\[17\] decoded_imm\[17\] VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__nand2_1
XFILLER_168_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12945__S net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08383_ _03796_ _03797_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07334_ net1063 net1026 _02874_ net1077 _02870_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__a221o_1
XANTENNA__08283__X net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10621__A1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07265_ _02792_ _02795_ _02808_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout1054_A mem_wordsize\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09004_ net356 net1760 net516 VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__mux2_1
X_07196_ reg_pc\[4\] decoded_imm\[4\] VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__nand2_1
XFILLER_133_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12374__A1 _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1221_A net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10924__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07250__B1 net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout500 net501 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__buf_4
XANTENNA_fanout681_A net696 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout511 _04278_ VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__buf_4
XANTENNA_fanout779_A net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11296__S net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout522 net523 VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__clkbuf_2
X_09906_ net1127 _04444_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__nor2_1
Xfanout533 net534 VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__buf_4
Xfanout544 _03766_ VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__clkbuf_2
Xfanout555 _03156_ VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__clkbuf_4
Xfanout566 _05080_ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__buf_2
Xfanout577 _03756_ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__clkbuf_2
X_09837_ _04615_ _04620_ net984 VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__a21o_1
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout588 _03749_ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10213__B net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_A _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout599 net600 VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout567_X net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09768_ _04556_ _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__and2_1
XANTENNA__07362__X _02901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08719_ _04076_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__inv_2
XANTENNA__07803__A net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09699_ decoded_imm_j\[6\] _04427_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13016__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11730_ latched_rd\[1\] _06242_ _06243_ net1465 VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11661_ decoded_imm_j\[11\] net13 net545 VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__mux2_1
XANTENNA__12855__S net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13400_ _02411_ net760 VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__nand2_1
X_10612_ cpuregs\[18\]\[7\] net553 _05304_ net780 VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__o22a_1
X_14380_ clknet_leaf_79_clk _00801_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dfxtp_4
X_11592_ mem_rdata_q\[29\] mem_rdata_q\[28\] VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__nor2_1
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08805__B2 net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13331_ net1010 net759 VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__or2_1
XANTENNA__10612__B2 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10543_ cpuregs\[19\]\[5\] net631 net595 VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__o21a_1
XFILLER_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13262_ _04940_ _04963_ _04971_ _04936_ _04937_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__a221o_1
XFILLER_155_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10474_ cpuregs\[5\]\[1\] net636 net817 _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__o211a_1
XFILLER_136_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15001_ clknet_leaf_147_clk net2916 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_12213_ genblk2.pcpi_div.quotient_msk\[20\] net270 net2761 VGND VGND VPWR VPWR _06599_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__12590__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13193_ net2158 net295 net429 VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__mux2_1
X_12144_ net2858 net383 net371 net2966 VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12117__A1 net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12075_ net724 _06523_ net1008 VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10404__A net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input30_X net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11026_ cpuregs\[18\]\[18\] net552 _05707_ net779 VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__o22a_1
XANTENNA_output231_A net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07272__X _02817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12977_ net1695 _03782_ net447 VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__mux2_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13309__A2_N _05527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14716_ clknet_leaf_156_clk _01101_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_11928_ _06392_ _06394_ _06395_ _06397_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__or4_1
X_14647_ clknet_leaf_161_clk _01032_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11859_ genblk2.pcpi_div.dividend\[7\] genblk2.pcpi_div.divisor\[7\] VGND VGND VPWR
+ VPWR _06330_ sky130_fd_sc_hd__nand2b_1
XFILLER_14_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14578_ clknet_leaf_93_clk _00964_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
XANTENNA__13250__C1 net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13529_ net520 net1443 net416 VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__mux2_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12066__A net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07050_ genblk2.pcpi_div.quotient\[18\] _02610_ net1116 VGND VGND VPWR VPWR _02617_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_11_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput103 net103 VGND VGND VPWR VPWR mem_la_wdata[15] sky130_fd_sc_hd__buf_2
Xoutput114 net114 VGND VGND VPWR VPWR mem_la_wdata[25] sky130_fd_sc_hd__buf_2
Xoutput125 net125 VGND VGND VPWR VPWR mem_la_wdata[6] sky130_fd_sc_hd__buf_2
Xoutput136 net136 VGND VGND VPWR VPWR mem_wdata[10] sky130_fd_sc_hd__buf_2
Xoutput147 net147 VGND VGND VPWR VPWR mem_wdata[20] sky130_fd_sc_hd__buf_2
XFILLER_142_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput158 net158 VGND VGND VPWR VPWR mem_wdata[30] sky130_fd_sc_hd__buf_2
Xoutput169 net169 VGND VGND VPWR VPWR mem_wstrb[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14431__D alu_out\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07952_ _03285_ _03422_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06903_ _02451_ _02486_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__nor2_1
XFILLER_56_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07883_ _03340_ _03398_ _03400_ _03336_ _03399_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__o221a_1
XFILLER_96_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09622_ _03811_ reg_next_pc\[17\] net922 VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__mux2_4
X_06834_ _02437_ _02438_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__and2b_1
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09314__S net479 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09553_ count_instr\[51\] count_instr\[50\] _04395_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__and3_1
X_06765_ net2584 VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__inv_2
XFILLER_71_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08504_ _03893_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09484_ count_instr\[26\] _04352_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__and2_1
XFILLER_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10842__A1 net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08435_ net311 net2406 net530 VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout527_A _03774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ reg_pc\[10\] _03780_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__xor2_1
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07317_ _02851_ _02856_ _02858_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__or3_1
X_08297_ net1002 _03732_ net982 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__mux2_1
XFILLER_20_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1057_X net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07248_ _02791_ _02793_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__or2_1
XFILLER_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout896_A net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12347__B2 mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07179_ net1062 _02719_ _02729_ net1082 _02722_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a221o_1
XFILLER_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout1224_X net1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10190_ decoded_imm\[28\] net996 VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__xor2_1
XFILLER_2_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10224__A decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout330 _03818_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_2
Xfanout341 _03807_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_2
Xfanout352 net353 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_2
Xfanout363 _06662_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__buf_4
XANTENNA_fanout851_X net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout374 net376 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_109_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11322__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout385 net388 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_2
XANTENNA_fanout949_X net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout396 net398 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_2
X_12900_ net571 net1967 net457 VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__mux2_1
XFILLER_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11754__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13880_ clknet_leaf_186_clk _00334_ VGND VGND VPWR VPWR cpuregs\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10878__B decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09224__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12831_ net587 net2308 net461 VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__mux2_1
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11086__A1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15550_ clknet_leaf_35_clk _01886_ VGND VGND VPWR VPWR cpuregs\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12762_ net1216 net1836 net2477 net907 _03876_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__a221o_1
X_14501_ clknet_leaf_93_clk _00890_ VGND VGND VPWR VPWR instr_srai sky130_fd_sc_hd__dfxtp_1
XFILLER_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11713_ net2163 net288 net375 VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__mux2_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15481_ clknet_leaf_9_clk _01817_ VGND VGND VPWR VPWR cpuregs\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12585__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12693_ net1211 genblk1.genblk1.pcpi_mul.next_rs2\[58\] net901 net2900 net713 VGND
+ VGND VPWR VPWR _01363_ sky130_fd_sc_hd__a221o_1
XFILLER_159_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14432_ clknet_leaf_100_clk _00821_ VGND VGND VPWR VPWR pcpi_timeout sky130_fd_sc_hd__dfxtp_1
XFILLER_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11644_ net2984 net21 net545 VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__mux2_1
X_14363_ clknet_leaf_133_clk _00784_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_1
Xinput16 mem_rdata[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xwire731 _06219_ VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__clkbuf_1
X_11575_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__inv_2
Xinput27 mem_rdata[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13314_ _02406_ net758 VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__nand2_1
X_10526_ cpuregs\[9\]\[5\] net630 net609 _05220_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__o211a_1
X_14294_ clknet_leaf_123_clk _00748_ VGND VGND VPWR VPWR count_cycle\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13245_ net1040 net396 _02171_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__o21ba_1
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10833__S net797 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10457_ cpuregs\[16\]\[0\] net554 _05156_ net784 VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__o22a_1
XANTENNA__08303__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13176_ net1755 net404 net428 VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10388_ _05089_ _05090_ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__or3_1
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12127_ net725 _06567_ net993 VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__a21oi_1
X_12058_ net1011 net721 _06508_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__nand3_1
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07517__A1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11664__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11009_ cpuregs\[11\]\[18\] net618 net589 _05690_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__o211a_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09134__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08973__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08220_ net1059 net1178 net1167 net942 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__a22o_1
XANTENNA__12026__B1 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11412__B net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08151_ _03626_ _03642_ _03628_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__o21ai_1
X_07102_ genblk2.pcpi_div.quotient\[26\] _02660_ net952 VGND VGND VPWR VPWR _02662_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08082_ net1161 _02407_ _03582_ net1143 VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12329__A1 decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12329__B2 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07033_ _02597_ _02598_ _02602_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10743__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09309__S net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11001__A1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07205__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07337__B decoded_imm\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08984_ genblk1.genblk1.pcpi_mul.rd\[30\] genblk1.genblk1.pcpi_mul.rd\[62\] net957
+ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__mux2_1
XFILLER_102_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07935_ _02366_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout477_A _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13355__A net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07866_ _03283_ _03318_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__or2_1
XANTENNA__10512__B1 net858 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09605_ reg_pc\[8\] net876 _04429_ net846 VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__a22o_1
XANTENNA__09044__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06817_ instr_slli instr_sb instr_lw instr_jalr VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout644_A net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07797_ net1169 net1035 VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nand2_1
XFILLER_25_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09536_ count_instr\[45\] count_instr\[44\] count_instr\[43\] _04382_ VGND VGND VPWR
+ VPWR _04387_ sky130_fd_sc_hd__and4_1
XANTENNA__12265__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ net2997 _04340_ net1229 VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_84_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10918__S net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net812 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1174_X net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11603__A net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12017__B1 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08418_ _03824_ _03825_ net768 VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__mux2_4
X_09398_ net190 net194 net192 net195 VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__or4_1
XFILLER_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08349_ reg_out\[7\] alu_out_q\[7\] net1153 VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__mux2_1
XANTENNA__10579__B1 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11360_ net833 _06028_ _06030_ _06032_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__a211o_1
XFILLER_164_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10311_ _04911_ _05010_ _05016_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__or3_1
XANTENNA__11749__S net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10653__S net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11291_ net1083 decoded_imm\[25\] _05133_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__o21a_1
X_13030_ net296 net2334 net445 VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__mux2_1
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09219__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10242_ decoded_imm\[3\] net1044 VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__and2_2
XFILLER_133_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12740__B2 net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10173_ net1068 net958 VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__nor2_2
XANTENNA__07247__B decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1103 net1104 VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__buf_2
Xfanout1114 net1116 VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__buf_2
Xfanout1125 net1126 VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09743__A decoded_imm_j\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1136 instr_rdinstr VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__buf_2
XFILLER_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1147 net1148 VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__clkbuf_2
X_14981_ clknet_leaf_107_clk _01333_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[28\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1158 net249 VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__buf_4
XFILLER_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1169 net1170 VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__buf_4
X_13932_ clknet_leaf_46_clk _00386_ VGND VGND VPWR VPWR cpuregs\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13863_ clknet_leaf_72_clk _00317_ VGND VGND VPWR VPWR cpuregs\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15602_ clknet_leaf_198_clk _01938_ VGND VGND VPWR VPWR cpuregs\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12814_ net338 net2189 net463 VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__mux2_1
XANTENNA__12256__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13794_ clknet_leaf_14_clk _00248_ VGND VGND VPWR VPWR cpuregs\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10806__A1 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15533_ clknet_leaf_20_clk _01869_ VGND VGND VPWR VPWR cpuregs\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12745_ net1328 net897 _02106_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__a21o_1
XFILLER_31_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12609__A _02392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ clknet_leaf_45_clk _01800_ VGND VGND VPWR VPWR cpuregs\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12676_ net1195 net2942 net888 net3006 net711 VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_139_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12328__B decoded_imm_j\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ clknet_leaf_176_clk alu_out\[15\] VGND VGND VPWR VPWR alu_out_q\[15\] sky130_fd_sc_hd__dfxtp_1
X_11627_ mem_rdata_q\[26\] _06204_ _06205_ mem_rdata_q\[27\] VGND VGND VPWR VPWR _06215_
+ sky130_fd_sc_hd__and4b_1
XANTENNA__08227__A2 net1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15395_ clknet_leaf_49_clk _01734_ VGND VGND VPWR VPWR cpuregs\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13220__A2 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07435__B1 net1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14346_ clknet_leaf_68_clk _06734_ VGND VGND VPWR VPWR reg_out\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11558_ mem_rdata_q\[14\] _06179_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__nor2_1
XANTENNA__11231__B2 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold608 cpuregs\[5\]\[7\] VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11659__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09196__Y _04286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10509_ net119 net860 _05206_ _03190_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__o22a_1
X_14277_ clknet_leaf_98_clk _00731_ VGND VGND VPWR VPWR count_cycle\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold619 cpuregs\[21\]\[14\] VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ net991 _02480_ _02487_ instr_jalr _06149_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__a221o_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13228_ reg_pc\[3\] net565 _02155_ _02156_ net392 VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__a221o_1
X_13159_ net1832 net300 net433 VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08968__S net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1308 genblk1.genblk1.pcpi_mul.rd\[32\] VGND VGND VPWR VPWR net2622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1319 genblk1.genblk1.pcpi_mul.next_rs2\[17\] VGND VGND VPWR VPWR net2633 sky130_fd_sc_hd__dlygate4sd3_1
X_07720_ cpuregs\[12\]\[4\] cpuregs\[13\]\[4\] net698 VGND VGND VPWR VPWR _03239_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11298__A1 net840 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08163__A1 net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07651_ _03162_ _03167_ _03171_ _03158_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__o211a_1
XANTENNA__15163__Q mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12247__B1 net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07582_ count_instr\[61\] net1133 net1137 count_instr\[29\] VGND VGND VPWR VPWR _03106_
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07901__A net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09321_ net1931 net310 net481 VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07620__B decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09252_ net1481 net312 net490 VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1248 VGND VGND VPWR VPWR picorv32_1248/HI eoi[6] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_32_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpicorv32_1259 VGND VGND VPWR VPWR picorv32_1259/HI eoi[17] sky130_fd_sc_hd__conb_1
X_08203_ _03372_ _03689_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__o21a_1
XFILLER_21_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08218__A2 net1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09183_ net326 net1783 net497 VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__mux2_1
XANTENNA__12953__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08134_ _03334_ _03619_ _03404_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_117_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08291__X net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08065_ _03378_ _03560_ _03377_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__o21ba_1
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1134_A instr_rdinstrh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07016_ net1115 _02587_ genblk2.pcpi_div.quotient\[14\] VGND VGND VPWR VPWR _02588_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__09039__S net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout594_A net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08967_ net2300 _04260_ net945 VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout382_X net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A _05134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07918_ net1163 _02406_ _03288_ _03433_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__o221ai_4
X_08898_ _03936_ _03938_ _03935_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__a21bo_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07849_ net1188 net1157 VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout647_X net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10860_ cpuregs\[30\]\[14\] cpuregs\[31\]\[14\] net664 VGND VGND VPWR VPWR _05546_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12238__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07811__A net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09519_ _04376_ net1226 _04375_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__and3b_1
XFILLER_25_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout814_X net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10791_ cpuregs\[1\]\[12\] net549 _05478_ net797 net823 VGND VGND VPWR VPWR _05479_
+ sky130_fd_sc_hd__a221o_1
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13024__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12530_ _02019_ net2653 net385 VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__mux2_1
XFILLER_157_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12461_ net1171 _06690_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__xor2_1
XFILLER_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13202__A2 net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14200_ clknet_leaf_173_clk _00654_ VGND VGND VPWR VPWR reg_pc\[8\] sky130_fd_sc_hd__dfxtp_1
X_11412_ cpuregs\[8\]\[29\] net704 VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__or2_1
XANTENNA__11213__A1 net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15180_ clknet_leaf_65_clk _01529_ VGND VGND VPWR VPWR mem_rdata_q\[31\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__09957__A2 net880 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12392_ net588 net1990 net474 VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__mux2_1
X_14131_ clknet_leaf_127_clk _00585_ VGND VGND VPWR VPWR count_instr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11343_ net793 _06011_ _06013_ _06015_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_134_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10972__B1 net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14062_ clknet_leaf_39_clk _00516_ VGND VGND VPWR VPWR cpuregs\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_11274_ _05947_ _05948_ net820 VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__mux2_1
XFILLER_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13013_ net403 net2134 net444 VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__mux2_1
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10225_ decoded_imm\[10\] net1029 VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__nand2_1
XANTENNA__07692__S net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10156_ _04868_ net1238 _04866_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__and3b_1
XANTENNA__12611__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 cpuregs\[0\]\[2\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10412__A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10087_ count_cycle\[32\] _04821_ count_cycle\[33\] VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__a21o_1
X_14964_ clknet_leaf_147_clk _01316_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13915_ clknet_leaf_5_clk _00369_ VGND VGND VPWR VPWR cpuregs\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14895_ clknet_leaf_140_clk _01247_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkload3_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13846_ clknet_leaf_187_clk _00300_ VGND VGND VPWR VPWR cpuregs\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13777_ clknet_leaf_22_clk _00231_ VGND VGND VPWR VPWR cpuregs\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10989_ cpuregs\[27\]\[17\] net617 net589 _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__o211a_1
XANTENNA__09645__B2 net850 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11243__A net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15516_ clknet_leaf_79_clk _01852_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07656__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12728_ net1190 genblk1.genblk1.pcpi_mul.next_rs1\[13\] net914 net1023 VGND VGND
+ VPWR VPWR _02098_ sky130_fd_sc_hd__a22o_1
XFILLER_148_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12058__B net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ net1212 genblk1.genblk1.pcpi_mul.next_rs2\[29\] net917 net255 VGND VGND VPWR
+ VPWR _02079_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15447_ clknet_leaf_41_clk _01786_ VGND VGND VPWR VPWR cpuregs\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12401__A0 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15378_ clknet_leaf_4_clk _01717_ VGND VGND VPWR VPWR cpuregs\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold405 cpuregs\[20\]\[26\] VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ clknet_leaf_171_clk _06747_ VGND VGND VPWR VPWR reg_out\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12074__A net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold416 cpuregs\[8\]\[3\] VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 cpuregs\[8\]\[17\] VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10963__B1 net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold438 cpuregs\[16\]\[16\] VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 cpuregs\[31\]\[17\] VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15158__Q mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12704__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout907 net910 VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__buf_2
X_09870_ _04651_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__inv_2
Xfanout918 net919 VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__buf_2
Xfanout929 _03463_ VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__buf_2
XFILLER_140_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07455__X _02988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08821_ genblk1.genblk1.pcpi_mul.next_rs2\[53\] net1102 _04160_ _04162_ VGND VGND
+ VPWR VPWR _04163_ sky130_fd_sc_hd__a22o_1
XANTENNA__06800__A net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1105 cpuregs\[1\]\[31\] VGND VGND VPWR VPWR net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13109__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1116 genblk1.genblk1.pcpi_mul.pcpi_rd\[13\] VGND VGND VPWR VPWR net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 cpuregs\[17\]\[30\] VGND VGND VPWR VPWR net2441 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _04104_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__inv_2
XFILLER_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1138 cpuregs\[18\]\[11\] VGND VGND VPWR VPWR net2452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__B1 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1149 cpuregs\[7\]\[28\] VGND VGND VPWR VPWR net2463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07703_ cpuregs\[19\]\[3\] net630 net595 VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__o21a_1
X_08683_ genblk1.genblk1.pcpi_mul.next_rs2\[32\] net1107 genblk1.genblk1.pcpi_mul.rd\[31\]
+ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__a21o_1
XANTENNA__12948__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07634_ cpuregs\[3\]\[2\] net640 net601 _03154_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__o211a_1
XANTENNA__11691__A1 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09322__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07565_ _03086_ _03089_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout342_A _03807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13432__A2 _04883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_A net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09304_ net1478 net540 net479 VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__mux2_1
XANTENNA__11153__A net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07496_ count_instr\[23\] net1137 net979 _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__a211o_1
XFILLER_167_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09235_ net1715 net543 net491 VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__mux2_1
XFILLER_22_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout607_A net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09558__A net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09166_ net580 net1774 net499 VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__mux2_1
XFILLER_163_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08117_ _03330_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09097_ net1889 net577 net504 VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08048_ _03434_ _03552_ net988 VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__mux2_1
Xhold950 genblk1.genblk1.pcpi_mul.next_rs1\[50\] VGND VGND VPWR VPWR net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout597_X net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold961 cpuregs\[8\]\[19\] VGND VGND VPWR VPWR net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A net979 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold972 genblk1.genblk1.pcpi_mul.next_rs1\[56\] VGND VGND VPWR VPWR net2286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold983 cpuregs\[1\]\[6\] VGND VGND VPWR VPWR net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 cpuregs\[19\]\[0\] VGND VGND VPWR VPWR net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_134_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12171__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10010_ count_cycle\[4\] count_cycle\[5\] _04771_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__and3_1
X_09999_ count_cycle\[0\] count_cycle\[1\] net1231 VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13019__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__A decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1650 genblk2.pcpi_div.divisor\[2\] VGND VGND VPWR VPWR net2964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1661 genblk1.genblk1.pcpi_mul.next_rs2\[42\] VGND VGND VPWR VPWR net2975 sky130_fd_sc_hd__dlygate4sd3_1
X_11961_ genblk2.pcpi_div.dividend\[4\] _06427_ net276 VGND VGND VPWR VPWR _01013_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout931_X net931 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1672 genblk2.pcpi_div.quotient_msk\[27\] VGND VGND VPWR VPWR net2986 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12858__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1683 count_instr\[20\] VGND VGND VPWR VPWR net2997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11762__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1694 mem_do_rdata VGND VGND VPWR VPWR net3008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13700_ clknet_leaf_107_clk _00154_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rdx\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_10912_ net822 _05592_ _05594_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a211o_1
XANTENNA__11682__A1 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14680_ clknet_leaf_153_clk net2868 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11892_ _06278_ _06362_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_158_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07350__A2 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09232__S net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13631_ clknet_leaf_120_clk _00085_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10843_ net1163 net854 _05528_ _05529_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__a22o_1
XANTENNA__09627__B2 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_143_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13562_ net520 net2232 net412 VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__mux2_1
X_10774_ cpuregs\[24\]\[12\] net650 VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__or2_1
XFILLER_44_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12513_ net1160 _05109_ net715 VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__or3_1
X_15301_ clknet_leaf_36_clk _01641_ VGND VGND VPWR VPWR cpuregs\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10642__C1 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12593__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13493_ net1856 net544 net419 VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_160_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_160_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_23_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15232_ clknet_leaf_20_clk _01573_ VGND VGND VPWR VPWR cpuregs\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12444_ net1180 net1178 net717 VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__o21ai_1
XFILLER_154_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15163_ clknet_leaf_65_clk _01512_ VGND VGND VPWR VPWR mem_rdata_q\[14\] sky130_fd_sc_hd__dfxtp_4
XFILLER_138_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12375_ net1388 net332 net360 VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__mux2_1
XANTENNA__10407__A net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11002__S net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14114_ clknet_leaf_11_clk _00568_ VGND VGND VPWR VPWR cpuregs\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11326_ net1083 decoded_imm\[26\] VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__or2_1
X_15094_ clknet_leaf_4_clk _01446_ VGND VGND VPWR VPWR cpuregs\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_152_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14045_ clknet_leaf_199_clk _00499_ VGND VGND VPWR VPWR cpuregs\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11257_ cpuregs\[0\]\[25\] net702 VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__or2_1
XFILLER_69_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10208_ decoded_imm\[17\] net1017 VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__nor2_1
XANTENNA_output69_A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11188_ net835 _05860_ _05862_ _05864_ net792 VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__a2111o_1
XFILLER_121_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10139_ _04856_ _04857_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__nor2_1
XFILLER_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14947_ clknet_leaf_35_clk _01299_ VGND VGND VPWR VPWR cpuregs\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11122__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09866__A1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11673__A1 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12870__A0 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14878_ clknet_leaf_17_clk _01230_ VGND VGND VPWR VPWR cpuregs\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09142__S net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13829_ clknet_leaf_23_clk _00283_ VGND VGND VPWR VPWR cpuregs\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07350_ net1063 net1024 _02889_ net1077 _02885_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__a221o_1
XFILLER_148_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07281_ _02807_ _02809_ _02824_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_151_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_151_clk sky130_fd_sc_hd__clkbuf_8
X_09020_ net296 net2090 net518 VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__mux2_1
XFILLER_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11420__B net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold202 cpuregs\[4\]\[26\] VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 cpuregs\[30\]\[31\] VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold224 cpuregs\[20\]\[23\] VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 cpuregs\[13\]\[6\] VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11627__A_N mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold246 cpuregs\[14\]\[25\] VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 cpuregs\[26\]\[26\] VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 genblk1.genblk1.pcpi_mul.next_rs1\[62\] VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 net58 VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10751__S net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09922_ net1150 _04698_ _04699_ net1184 VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__o31a_1
XANTENNA__12532__A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout704 net705 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__buf_2
XANTENNA__06801__Y _02409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout715 net716 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__clkbuf_2
Xfanout726 _06409_ VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__buf_2
XANTENNA__13350__A1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09317__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout737 net738 VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09853_ net1182 _04439_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__or2_1
XANTENNA__13347__B _05710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout748 net749 VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__buf_2
XANTENNA_fanout292_A _03860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout759 _04884_ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08804_ _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__inv_2
X_09784_ _04556_ _04572_ _04568_ _04547_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__o2bb2a_1
X_06996_ net1118 _02569_ genblk2.pcpi_div.dividend\[11\] VGND VGND VPWR VPWR _02571_
+ sky130_fd_sc_hd__a21oi_1
X_08735_ genblk1.genblk1.pcpi_mul.next_rs2\[40\] net1094 genblk1.genblk1.pcpi_mul.rd\[39\]
+ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout557_A _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13363__A net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07632__Y _03153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08666_ genblk1.genblk1.pcpi_mul.next_rs2\[29\] net1106 _04028_ _04030_ VGND VGND
+ VPWR VPWR _04032_ sky130_fd_sc_hd__and4_1
XANTENNA__11664__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09052__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07617_ net986 decoded_imm_j\[11\] VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__or2_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08597_ net890 _03971_ _03973_ net2838 net1196 VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__a32o_1
XANTENNA__08176__B net935 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_X net1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11416__A1 net795 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10219__A2 net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07548_ _03058_ _03061_ _03073_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_153_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08293__A0 net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout512_X net512 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_142_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_142_clk sky130_fd_sc_hd__clkbuf_8
X_07479_ _02993_ _02997_ _03008_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__a21o_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09218_ net1511 net319 net493 VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10490_ _05187_ _05188_ net816 VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__mux2_1
XFILLER_136_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ net1687 net330 net500 VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__mux2_1
XFILLER_136_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12160_ genblk2.pcpi_div.quotient_msk\[19\] net377 net365 net2794 VGND VGND VPWR
+ VPWR _01061_ sky130_fd_sc_hd__a22o_1
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout881_X net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout979_X net979 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11757__S net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11111_ net804 _05787_ _05789_ net840 VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__a211o_1
XFILLER_151_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12091_ net1005 net724 _06536_ net863 VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__a31o_1
Xhold780 cpuregs\[21\]\[23\] VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 genblk1.genblk1.pcpi_mul.next_rs1\[21\] VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09227__S net495 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12144__A2 net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13341__A1 net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11042_ net816 _05722_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__or2_1
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A mem_rdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ clknet_leaf_75_clk _01153_ VGND VGND VPWR VPWR decoded_imm\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12588__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12993_ net1510 net303 net450 VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__mux2_1
XFILLER_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1480 genblk2.pcpi_div.quotient_msk\[20\] VGND VGND VPWR VPWR net2794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13273__A net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1491 count_instr\[31\] VGND VGND VPWR VPWR net2805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11655__A1 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14732_ clknet_leaf_163_clk net2705 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11944_ _02443_ net726 net1046 VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11875_ _06343_ _06345_ _06299_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__a21o_1
X_14663_ clknet_leaf_151_clk _01048_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10826_ cpuregs\[24\]\[13\] net650 VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__or2_1
X_13614_ clknet_leaf_42_clk _00069_ VGND VGND VPWR VPWR cpuregs\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14594_ clknet_leaf_115_clk _00980_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11958__A2 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10757_ cpuregs\[14\]\[11\] cpuregs\[15\]\[11\] net666 VGND VGND VPWR VPWR _05446_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13545_ net306 net2072 net418 VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_133_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_133_clk sky130_fd_sc_hd__clkbuf_8
X_13476_ net1445 net317 net423 VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__mux2_1
XANTENNA__08306__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10688_ cpuregs\[22\]\[9\] cpuregs\[23\]\[9\] net671 VGND VGND VPWR VPWR _05379_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12336__B decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15215_ clknet_leaf_88_clk _00004_ VGND VGND VPWR VPWR cpu_state\[0\] sky130_fd_sc_hd__dfxtp_1
X_12427_ net917 _06665_ _06666_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__or3b_1
XFILLER_126_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12358_ net1873 net586 net362 VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__mux2_1
X_15146_ clknet_leaf_80_clk _06748_ VGND VGND VPWR VPWR reg_sh\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11309_ cpuregs\[28\]\[26\] cpuregs\[29\]\[26\] net703 VGND VGND VPWR VPWR _05983_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15077_ clknet_leaf_103_clk _01429_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12289_ mem_rdata_q\[29\] _06622_ _06623_ _06620_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_39_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14028_ clknet_leaf_53_clk _00482_ VGND VGND VPWR VPWR cpuregs\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09137__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08041__S net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06850_ mem_do_prefetch _02452_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__nand2_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08976__S net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10697__A2 _05386_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06781_ genblk2.pcpi_div.dividend\[30\] VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__inv_2
X_08520_ genblk1.genblk1.pcpi_mul.next_rs2\[7\] net1097 genblk1.genblk1.pcpi_mul.rd\[6\]
+ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__a21o_1
XANTENNA__10449__A2 net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11646__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08451_ net297 net2217 net531 VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__mux2_1
XFILLER_36_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10854__C1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14429__D alu_out\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15171__Q mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07402_ net1071 _02930_ _02931_ _02938_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__a31o_1
XFILLER_51_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08382_ reg_pc\[13\] reg_pc\[12\] _03789_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__and3_1
XANTENNA__09600__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08275__A0 net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07333_ genblk1.genblk1.pcpi_mul.pcpi_rd\[12\] genblk2.pcpi_div.pcpi_rd\[12\] net1110
+ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_124_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13122__S net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07264_ _02792_ _02795_ _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__a21o_1
X_09003_ net403 net1767 net517 VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__14515__Q decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13020__A0 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07195_ net1065 net1044 _02736_ _02744_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__a211o_1
XANTENNA__12961__S net454 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10909__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A _03844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1047_A net1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07627__Y _03148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13358__A net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10481__S net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout501 net503 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1214_A net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09047__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout512 net513 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_4
XFILLER_99_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09905_ net1128 _04444_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__and2_1
XFILLER_160_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout523 _03777_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkbuf_2
Xfanout534 _06240_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__buf_8
XANTENNA_fanout674_A net676 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout545 net546 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__clkbuf_4
Xfanout556 net557 VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__buf_2
Xfanout567 net570 VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkbuf_4
X_09836_ _04615_ _04620_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__nor2_1
Xfanout578 _03756_ VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1002_X net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout589 net590 VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout462_X net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06979_ genblk2.pcpi_div.quotient\[7\] genblk2.pcpi_div.quotient\[8\] _02544_ VGND
+ VGND VPWR VPWR _02556_ sky130_fd_sc_hd__or3_1
X_09767_ decoded_imm_j\[12\] _04433_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout841_A net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A _02693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11098__C1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08718_ genblk1.genblk1.pcpi_mul.next_rs2\[37\] net1099 _04072_ _04074_ VGND VGND
+ VPWR VPWR _04076_ sky130_fd_sc_hd__and4_1
XFILLER_92_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07803__B net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09698_ decoded_imm_j\[6\] _04427_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__and2_1
XFILLER_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ net902 _04015_ _04017_ net2781 net1212 VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_25_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_X net727 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11660_ decoded_imm_j\[18\] net10 net546 VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__mux2_1
XFILLER_42_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10611_ cpuregs\[19\]\[7\] net626 net593 VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__o21a_1
X_11591_ net2896 net740 _06190_ is_sb_sh_sw VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_115_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13032__S net446 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13330_ net567 _05637_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__nor2_1
XFILLER_128_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10542_ cpuregs\[17\]\[5\] net629 net609 _05236_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__o211a_1
XANTENNA__10612__A2 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13261_ _02180_ _02181_ _02185_ net395 net1035 VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__o32a_1
X_10473_ cpuregs\[4\]\[1\] net692 VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__or2_1
X_12212_ net748 net2813 VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__nor2_1
XFILLER_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15000_ clknet_leaf_147_clk _01352_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_13192_ net2303 net300 net429 VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__mux2_1
XFILLER_124_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07241__A1 net1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12143_ net2750 net382 net372 net2858 VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__a22o_1
XANTENNA__07241__B2 net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12074_ net1011 net1009 _06508_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__or3_1
XFILLER_104_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11025_ cpuregs\[19\]\[18\] net618 net589 VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__o21a_1
XFILLER_77_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input23_X net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output224_A net995 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11628__A1 instr_rdcycleh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12976_ net1712 net523 net447 VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__mux2_1
X_14715_ clknet_leaf_154_clk _01100_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11235__B net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11927_ _06389_ _06390_ _06391_ _06396_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__or4_2
X_14646_ clknet_leaf_161_clk _01031_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08384__X _03799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11858_ genblk2.pcpi_div.divisor\[6\] _02391_ _06328_ VGND VGND VPWR VPWR _06329_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__08257__A0 net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_106_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_8
X_10809_ cpuregs\[5\]\[13\] net620 net812 _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__o211a_1
X_14577_ clknet_leaf_96_clk _00963_ VGND VGND VPWR VPWR is_compare sky130_fd_sc_hd__dfxtp_1
X_11789_ genblk2.pcpi_div.divisor\[30\] genblk2.pcpi_div.dividend\[30\] VGND VGND
+ VPWR VPWR _06260_ sky130_fd_sc_hd__xor2_1
XANTENNA__11251__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13528_ net524 net1722 net416 VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__mux2_1
XANTENNA__10603__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11261__C1 net786 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_191_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13459_ net1413 net571 net426 VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09656__A decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput104 net104 VGND VGND VPWR VPWR mem_la_wdata[16] sky130_fd_sc_hd__buf_2
Xoutput115 net115 VGND VGND VPWR VPWR mem_la_wdata[26] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput126 net1170 VGND VGND VPWR VPWR mem_la_wdata[7] sky130_fd_sc_hd__buf_2
Xoutput137 net137 VGND VGND VPWR VPWR mem_wdata[11] sky130_fd_sc_hd__buf_2
X_15129_ clknet_leaf_0_clk _01481_ VGND VGND VPWR VPWR cpuregs\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xoutput148 net148 VGND VGND VPWR VPWR mem_wdata[21] sky130_fd_sc_hd__buf_2
Xoutput159 net159 VGND VGND VPWR VPWR mem_wdata[31] sky130_fd_sc_hd__buf_2
XFILLER_88_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13305__A1 net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07951_ net967 _03284_ _03285_ net928 _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__a221o_1
XANTENNA__15166__Q mem_rdata_q\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06902_ is_jalr_addi_slti_sltiu_xori_ori_andi is_lui_auipc_jal net1088 VGND VGND
+ VPWR VPWR _02497_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07882_ net244 net1015 VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__nand2b_1
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06833_ genblk1.genblk1.pcpi_mul.pcpi_ready net1113 VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__nor2_1
X_09621_ net3061 net877 _04437_ net847 VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__a22o_1
XANTENNA__13117__S net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09552_ _04396_ _04397_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__nor2_1
X_06764_ net2590 VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__inv_2
XANTENNA__10330__A net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08503_ _03887_ _03890_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__nand2_1
XFILLER_102_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09483_ _04352_ _04353_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__nor2_1
XFILLER_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12956__S net452 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_144_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08434_ _03837_ _03838_ net768 VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__mux2_1
XANTENNA__10842__A2 _05527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06954__S net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ reg_out\[10\] alu_out_q\[10\] net1153 VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__mux2_1
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07316_ net1063 net1028 _02857_ net1077 _02853_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__a221o_1
XANTENNA__11252__C1 net858 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08296_ reg_out\[25\] reg_next_pc\[25\] net925 VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_159_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07247_ reg_pc\[7\] decoded_imm\[7\] VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__nor2_1
XFILLER_164_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12347__A2 decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07178_ genblk1.genblk1.pcpi_mul.pcpi_rd\[2\] genblk2.pcpi_div.pcpi_rd\[2\] net1111
+ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout791_A net795 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout320 _03826_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10224__B net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout331 _03818_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_1
Xfanout342 _03807_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_1
Xfanout353 _03794_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout364 net370 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout375 net376 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_8
XFILLER_4_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout386 net388 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_2
XANTENNA__07814__A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout397 net398 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09819_ decoded_imm_j\[16\] _04437_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_161_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12830_ _03742_ _04283_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__or2_4
XFILLER_28_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10240__A decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12761_ net1836 net905 _02114_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__a21o_1
XANTENNA__11770__S net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14500_ clknet_leaf_94_clk _00889_ VGND VGND VPWR VPWR instr_and sky130_fd_sc_hd__dfxtp_1
X_11712_ net2040 net292 net376 VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__mux2_1
XANTENNA__11491__C1 net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15480_ clknet_leaf_9_clk _01816_ VGND VGND VPWR VPWR cpuregs\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12692_ net1211 net2900 net903 net2952 net713 VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__a221o_1
XANTENNA__09240__S net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10894__B net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08239__A0 net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14431_ clknet_leaf_87_clk alu_out\[31\] VGND VGND VPWR VPWR alu_out_q\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13232__A0 net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11643_ decoded_imm_j\[7\] net20 net545 VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__mux2_1
XFILLER_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09987__B1 net1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11574_ mem_rdata_q\[14\] mem_rdata_q\[12\] mem_rdata_q\[13\] VGND VGND VPWR VPWR
+ _06188_ sky130_fd_sc_hd__or3b_2
X_14362_ clknet_leaf_82_clk _00783_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_1
XFILLER_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 mem_rdata[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput28 mem_rdata[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XFILLER_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13313_ net567 _05563_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__nor2_1
X_10525_ cpuregs\[8\]\[5\] net675 VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__or2_1
X_14293_ clknet_leaf_123_clk _00747_ VGND VGND VPWR VPWR count_cycle\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13244_ net568 _05242_ _02165_ net960 _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__o221a_1
XFILLER_109_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10456_ cpuregs\[17\]\[0\] net635 net611 VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__o21a_1
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13175_ net1824 net407 net427 VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__mux2_1
XANTENNA__10415__A net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10387_ genblk2.pcpi_div.quotient_msk\[19\] genblk2.pcpi_div.quotient_msk\[18\] genblk2.pcpi_div.quotient_msk\[17\]
+ genblk2.pcpi_div.quotient_msk\[16\] VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__or4_1
XANTENNA__07708__B _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12126_ net997 net995 _06558_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__or3_1
XANTENNA__13299__B1 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12057_ net1013 _06501_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__or2_1
XFILLER_78_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11008_ cpuregs\[10\]\[18\] net647 VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__or2_1
XFILLER_65_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12959_ net306 net2209 net453 VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__mux2_1
XFILLER_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09150__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12026__A1 net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14629_ clknet_leaf_139_clk _01014_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10037__B1 net1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08150_ _03320_ _03325_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__nand2_1
XANTENNA__11785__B1 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07101_ genblk2.pcpi_div.quotient\[26\] _02660_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__or2_1
X_08081_ _03343_ _03437_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__or2_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07453__B2 net1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07032_ _02600_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__or2_1
XANTENNA__12329__A2 net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11537__A0 mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06803__A net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07205__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12016__S net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07205__B2 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ net1504 _04268_ net946 VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__mux2_1
XANTENNA__10760__A1 net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06964__B1 net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07934_ _03369_ _03394_ _03450_ _03393_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__a31o_1
XANTENNA__12540__A net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08289__X net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09325__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07193__X _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07865_ _03278_ _03311_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__nand2_1
XFILLER_84_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _03775_ reg_next_pc\[8\] net921 VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__mux2_2
X_06816_ net1134 instr_rdcycleh instr_rdinstr VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__or3_1
XANTENNA__07353__B decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07796_ _03312_ _03313_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__nand2_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09535_ _04386_ net1227 _04385_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__and3b_1
XFILLER_25_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout637_A net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09466_ count_instr\[20\] count_instr\[19\] _04338_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__and3_1
XFILLER_25_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11603__B mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12017__A1 net1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08417_ reg_pc\[20\] _03821_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__xor2_1
X_09397_ net267 net1234 net171 net182 VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_35_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout425_X net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_A net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1167_X net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08348_ net539 net2279 net528 VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__mux2_1
XFILLER_165_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08279_ net1018 _03723_ net981 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__mux2_2
XFILLER_164_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13517__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10310_ _04910_ _05015_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__or2_1
X_11290_ net1083 _05964_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__nand2_1
XANTENNA__11528__A0 mem_rdata_q\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08404__S net767 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_X net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10241_ decoded_imm\[4\] net1042 VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__nand2_2
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10235__A decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10172_ _04878_ _04877_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_163_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout961_X net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06955__B1 net1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1104 net1109 VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1115 net1116 VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__buf_2
Xfanout1126 genblk2.pcpi_div.outsign VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__buf_2
Xfanout1137 net1138 VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__buf_2
X_14980_ clknet_leaf_108_clk _01332_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1148 net1149 VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout1159 net245 VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__buf_4
XANTENNA__09235__S net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13931_ clknet_leaf_72_clk _00385_ VGND VGND VPWR VPWR cpuregs\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10503__A1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11066__A net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13862_ clknet_leaf_36_clk _00316_ VGND VGND VPWR VPWR cpuregs\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15601_ clknet_leaf_191_clk _01937_ VGND VGND VPWR VPWR cpuregs\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12813_ net341 net1972 net463 VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__mux2_1
XFILLER_62_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12596__S net468 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13793_ clknet_leaf_41_clk _00247_ VGND VGND VPWR VPWR cpuregs\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15532_ clknet_leaf_21_clk _01868_ VGND VGND VPWR VPWR cpuregs\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10806__A2 net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12744_ net1191 genblk1.genblk1.pcpi_mul.next_rs1\[21\] net916 net1008 VGND VGND
+ VPWR VPWR _02106_ sky130_fd_sc_hd__a22o_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12609__B net912 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12008__A1 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ clknet_leaf_38_clk _01799_ VGND VGND VPWR VPWR cpuregs\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12675_ net1195 net3006 net889 genblk1.genblk1.pcpi_mul.next_rs2\[39\] net712 VGND
+ VGND VPWR VPWR _01345_ sky130_fd_sc_hd__a221o_1
XFILLER_30_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__A2 net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14414_ clknet_leaf_177_clk alu_out\[14\] VGND VGND VPWR VPWR alu_out_q\[14\] sky130_fd_sc_hd__dfxtp_1
X_11626_ net3057 net737 _06206_ _06214_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_139_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ clknet_leaf_53_clk _01733_ VGND VGND VPWR VPWR cpuregs\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14345_ clknet_leaf_82_clk _06733_ VGND VGND VPWR VPWR reg_out\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11231__A2 net555 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11557_ mem_rdata_q\[13\] mem_rdata_q\[12\] VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__nand2b_1
XFILLER_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold609 cpuregs\[6\]\[28\] VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ net987 decoded_imm\[2\] net856 VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__a21o_1
XANTENNA__11519__A0 mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14276_ clknet_leaf_97_clk _00730_ VGND VGND VPWR VPWR count_cycle\[21\] sky130_fd_sc_hd__dfxtp_1
X_11488_ net1072 _02370_ _02487_ net1156 net1232 VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__o221a_1
XANTENNA_output99_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10990__A1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13227_ net1063 net1035 net754 net557 VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__a31o_1
X_10439_ cpuregs\[3\]\[0\] net634 net597 _05138_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__o211a_1
XFILLER_98_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13158_ net1412 net303 net434 VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__mux2_1
XANTENNA__10742__A1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12109_ _06373_ _06548_ _06372_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__a21oi_1
X_13089_ net308 net1814 net440 VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1309 genblk2.pcpi_div.divisor\[45\] VGND VGND VPWR VPWR net2623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09145__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09360__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07650_ net825 net799 net552 net776 VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__o31a_4
XANTENNA__08984__S net957 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07581_ net359 _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__nor2_1
X_09320_ net1400 net313 net481 VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09251_ net1591 net316 net490 VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__mux2_1
Xpicorv32_1249 VGND VGND VPWR VPWR picorv32_1249/HI eoi[7] sky130_fd_sc_hd__conb_1
X_08202_ _03372_ _03689_ _03465_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09182_ net330 net1729 net497 VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__mux2_1
X_08133_ _03611_ _03626_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13130__S net438 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06804__Y _02412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08064_ _02394_ net1023 _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__a21o_1
XANTENNA__07629__A net1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07015_ genblk2.pcpi_div.quotient\[12\] genblk2.pcpi_div.quotient\[13\] _02575_ VGND
+ VGND VPWR VPWR _02587_ sky130_fd_sc_hd__or3_1
XANTENNA__10981__B2 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1127_A net1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout587_A _03749_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07635__Y _03156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08966_ genblk1.genblk1.pcpi_mul.rd\[21\] genblk1.genblk1.pcpi_mul.rd\[53\] net956
+ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__mux2_1
XANTENNA__09055__S net514 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07917_ net1164 _02405_ _03288_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout375_X net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08897_ net1195 net2646 net888 _04225_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout754_A net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_57_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ net1188 net1157 VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__nand2_1
XFILLER_83_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout921_A net927 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07779_ _03295_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__and2_1
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07811__B net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09518_ count_instr\[38\] count_instr\[37\] _04372_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__and3_1
X_10790_ cpuregs\[2\]\[12\] cpuregs\[3\]\[12\] net659 VGND VGND VPWR VPWR _05478_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07114__B1 net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09449_ net2779 _04328_ net1228 VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout807_X net807 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12460_ net1172 net1175 _05098_ net717 VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__o31a_1
XFILLER_138_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11411_ net819 _06079_ _06081_ net836 VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__o211a_1
XANTENNA__09297__Y _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12391_ _04273_ _06663_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__or2_2
XANTENNA__10664__S net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12445__A net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13040__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11342_ cpuregs\[11\]\[27\] net639 net598 _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__o211a_1
XFILLER_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14130_ clknet_leaf_83_clk _00584_ VGND VGND VPWR VPWR count_instr\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14061_ clknet_leaf_50_clk _00515_ VGND VGND VPWR VPWR cpuregs\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_11273_ cpuregs\[20\]\[25\] cpuregs\[21\]\[25\] net702 VGND VGND VPWR VPWR _05948_
+ sky130_fd_sc_hd__mux2_1
X_13012_ net408 net2317 net443 VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__mux2_1
X_10224_ decoded_imm\[11\] net1028 VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__or2_1
XANTENNA__12713__A2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10155_ count_cycle\[54\] count_cycle\[55\] _04860_ _04867_ VGND VGND VPWR VPWR _04868_
+ sky130_fd_sc_hd__and4_1
XANTENNA__12180__A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11067__Y _05748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10086_ net3062 _04821_ _04823_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__o21a_1
X_14963_ clknet_leaf_147_clk _01315_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold6 cpuregs\[0\]\[16\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_8
X_13914_ clknet_leaf_6_clk _00368_ VGND VGND VPWR VPWR cpuregs\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14894_ clknet_leaf_140_clk _01246_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13845_ clknet_leaf_190_clk _00299_ VGND VGND VPWR VPWR cpuregs\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08309__S net983 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07105__B1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13776_ clknet_leaf_32_clk _00230_ VGND VGND VPWR VPWR cpuregs\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09645__A2 net880 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10988_ cpuregs\[26\]\[17\] net649 VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__or2_1
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11988__B1 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15515_ clknet_leaf_78_clk _01851_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dfxtp_1
X_12727_ net1190 net2133 net2421 net883 _02097_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15446_ clknet_leaf_9_clk _01785_ VGND VGND VPWR VPWR cpuregs\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12658_ net1212 net2730 net902 net3009 _02078_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_61_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07408__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11609_ instr_srl net561 _06183_ _06201_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__a22o_1
X_15377_ clknet_leaf_3_clk _01716_ VGND VGND VPWR VPWR cpuregs\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12589_ net338 net2141 net468 VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__mux2_1
XFILLER_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14328_ clknet_leaf_172_clk _06746_ VGND VGND VPWR VPWR reg_out\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_128_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12074__B net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold406 cpuregs\[13\]\[20\] VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 genblk1.genblk1.pcpi_mul.pcpi_rd\[22\] VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 cpuregs\[14\]\[24\] VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 cpuregs\[13\]\[5\] VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ clknet_leaf_128_clk _00713_ VGND VGND VPWR VPWR count_cycle\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_143_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09664__A decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout908 net910 VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__buf_2
Xfanout919 _03874_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__buf_2
X_08820_ genblk1.genblk1.pcpi_mul.rd\[52\] genblk1.genblk1.pcpi_mul.rdx\[52\] VGND
+ VGND VPWR VPWR _04162_ sky130_fd_sc_hd__or2_1
Xhold1106 reg_next_pc\[18\] VGND VGND VPWR VPWR net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 cpuregs\[17\]\[31\] VGND VGND VPWR VPWR net2431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1128 cpuregs\[27\]\[25\] VGND VGND VPWR VPWR net2442 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _04095_ _04098_ _04100_ _04102_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__o211a_1
XANTENNA__12468__A1 net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15174__Q mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10322__B net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_8
Xhold1139 cpuregs\[3\]\[29\] VGND VGND VPWR VPWR net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_07702_ cpuregs\[17\]\[3\] net630 _03148_ _03221_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__o211a_1
X_08682_ genblk1.genblk1.pcpi_mul.rd\[31\] genblk1.genblk1.pcpi_mul.next_rs2\[32\]
+ net1107 VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__nand3_1
XFILLER_26_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07633_ cpuregs\[2\]\[2\] net699 VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__or2_1
XANTENNA__13417__B1 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13125__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07564_ _03087_ _03088_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09303_ net1455 net542 net480 VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__mux2_1
XFILLER_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07495_ count_instr\[55\] net1133 net1141 count_cycle\[55\] VGND VGND VPWR VPWR _03025_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12964__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout335_A _03815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_A net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09234_ net1658 net574 net491 VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__mux2_1
XFILLER_22_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09165_ net585 net2320 net498 VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout502_A net503 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08116_ _03612_ _03613_ net1143 VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__mux2_1
X_09096_ net2047 net581 net507 VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08047_ _03299_ _03546_ _03298_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_79_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold940 cpuregs\[1\]\[4\] VGND VGND VPWR VPWR net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _01420_ VGND VGND VPWR VPWR net2265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 cpuregs\[11\]\[20\] VGND VGND VPWR VPWR net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold973 cpuregs\[19\]\[25\] VGND VGND VPWR VPWR net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold984 cpuregs\[1\]\[12\] VGND VGND VPWR VPWR net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 cpuregs\[18\]\[7\] VGND VGND VPWR VPWR net2309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout969_A _02432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09998_ net1206 net2605 VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__nor2_1
XANTENNA__07583__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08949_ net2549 _04251_ net943 VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__B net1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_X net757 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1640 count_instr\[51\] VGND VGND VPWR VPWR net2954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1651 _01107_ VGND VGND VPWR VPWR net2965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1662 count_instr\[27\] VGND VGND VPWR VPWR net2976 sky130_fd_sc_hd__dlygate4sd3_1
X_11960_ net866 _06326_ _06426_ _06425_ _06424_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__a32o_1
Xhold1673 count_cycle\[27\] VGND VGND VPWR VPWR net2987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11131__A1 net824 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1684 count_instr\[24\] VGND VGND VPWR VPWR net2998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1695 genblk1.genblk1.pcpi_mul.next_rs2\[27\] VGND VGND VPWR VPWR net3009 sky130_fd_sc_hd__dlygate4sd3_1
X_10911_ cpuregs\[18\]\[15\] net552 _05595_ net779 VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__o22a_1
XFILLER_45_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07886__A1 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11682__A2 net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout924_X net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11891_ _06358_ _06361_ _06360_ _06282_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_158_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13035__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13630_ clknet_leaf_120_clk _00084_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10842_ net1075 _05527_ net854 VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09627__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13561_ net524 net2396 net412 VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__mux2_1
X_10773_ _05459_ _05460_ net797 VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__mux2_1
XFILLER_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15300_ clknet_leaf_102_clk net1315 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_wait_q
+ sky130_fd_sc_hd__dfxtp_1
X_12512_ _05109_ net715 net1160 VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_136_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13492_ net1485 net572 net422 VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__mux2_1
XFILLER_157_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ clknet_leaf_180_clk _01572_ VGND VGND VPWR VPWR cpuregs\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12443_ _06677_ net2771 net383 VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__mux2_1
X_15162_ clknet_leaf_65_clk _01511_ VGND VGND VPWR VPWR mem_rdata_q\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12374_ net1452 _03810_ net361 VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__mux2_1
XFILLER_165_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10407__B net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14113_ clknet_leaf_41_clk _00567_ VGND VGND VPWR VPWR cpuregs\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_11325_ net775 _05990_ _05998_ _05982_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__a31oi_4
XFILLER_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15093_ clknet_leaf_194_clk _01445_ VGND VGND VPWR VPWR cpuregs\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12147__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14044_ clknet_leaf_195_clk _00498_ VGND VGND VPWR VPWR cpuregs\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11256_ _05929_ _05930_ net820 VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__mux2_1
XANTENNA_output254_A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10207_ decoded_imm\[20\] net1010 VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__nand2_1
XANTENNA__12114__S net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11187_ cpuregs\[27\]\[23\] net634 net600 _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__o211a_1
XFILLER_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11370__A1 net840 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10138_ count_cycle\[51\] _04854_ net1235 VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_59_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_10_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10069_ count_cycle\[26\] _04811_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__and2_1
X_14946_ clknet_leaf_17_clk _01298_ VGND VGND VPWR VPWR cpuregs\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12870__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10569__S net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14877_ clknet_leaf_36_clk _01229_ VGND VGND VPWR VPWR cpuregs\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13828_ clknet_leaf_43_clk _00282_ VGND VGND VPWR VPWR cpuregs\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13759_ clknet_leaf_9_clk _00213_ VGND VGND VPWR VPWR cpuregs\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07280_ _02821_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__nand2_1
XANTENNA__09659__A decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15429_ clknet_leaf_45_clk _01768_ VGND VGND VPWR VPWR cpuregs\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15169__Q mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold203 cpuregs\[23\]\[4\] VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 cpuregs\[22\]\[16\] VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 cpuregs\[29\]\[0\] VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 genblk1.genblk1.pcpi_mul.next_rs1\[25\] VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold247 cpuregs\[10\]\[18\] VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 cpuregs\[20\]\[0\] VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 cpuregs\[14\]\[6\] VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _04443_ _04444_ _04445_ _04673_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__and4_1
Xfanout705 net707 VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__clkbuf_2
Xfanout716 _06674_ VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__clkbuf_2
Xfanout727 net728 VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ net1146 _04634_ _04635_ _04633_ net1182 VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__o311ai_1
Xfanout738 net739 VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10333__A net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11361__A1 net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout749 net750 VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__buf_2
XANTENNA__07137__B1_N _02443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08803_ _04139_ _04142_ _04144_ _04146_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__o211a_1
XFILLER_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09783_ _04543_ _04557_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12959__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06995_ genblk2.pcpi_div.dividend\[11\] net1118 _02569_ VGND VGND VPWR VPWR _02570_
+ sky130_fd_sc_hd__and3_1
XANTENNA__09306__A1 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08734_ genblk1.genblk1.pcpi_mul.rd\[39\] genblk1.genblk1.pcpi_mul.next_rs2\[40\]
+ net1094 VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__nand3_1
XANTENNA__08297__X net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11113__B2 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12310__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09333__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08665_ genblk1.genblk1.pcpi_mul.next_rs2\[29\] net1106 _04028_ _04030_ VGND VGND
+ VPWR VPWR _04031_ sky130_fd_sc_hd__a22o_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout452_A net454 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10872__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07616_ net986 decoded_imm_j\[2\] _03135_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__o21a_2
XANTENNA__09609__A2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08596_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__inv_2
X_07547_ _03071_ _03072_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout717_A net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ _02976_ _02995_ _02993_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_153_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09217_ net1606 net322 net493 VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout505_X net505 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09148_ net1763 net333 net500 VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__mux2_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09079_ net1471 net328 net508 VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__mux2_1
XFILLER_107_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11110_ cpuregs\[5\]\[21\] net634 net818 _05788_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_9_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12090_ net724 _06536_ net1005 VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold770 cpuregs\[8\]\[31\] VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout874_X net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold781 cpuregs\[1\]\[24\] VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _01391_ VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ cpuregs\[14\]\[19\] cpuregs\[15\]\[19\] net680 VGND VGND VPWR VPWR _05722_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11352__A1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ clknet_leaf_75_clk _01152_ VGND VGND VPWR VPWR decoded_imm\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_129_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ net1381 net307 net449 VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__mux2_1
XANTENNA__09243__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1470 count_cycle\[12\] VGND VGND VPWR VPWR net2784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input13_A mem_rdata[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1481 _01061_ VGND VGND VPWR VPWR net2795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14731_ clknet_leaf_170_clk _01116_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold1492 genblk2.pcpi_div.quotient\[28\] VGND VGND VPWR VPWR net2806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11943_ genblk2.pcpi_div.dividend\[1\] _06412_ net276 VGND VGND VPWR VPWR _01010_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ clknet_leaf_138_clk _01047_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11874_ _06344_ _06332_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_28_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ clknet_leaf_1_clk _00068_ VGND VGND VPWR VPWR cpuregs\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_10825_ _05510_ _05511_ net796 VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__mux2_1
X_14593_ clknet_leaf_156_clk _00979_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dfxtp_1
XFILLER_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13544_ net310 net2111 net417 VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__mux2_1
X_10756_ net839 _05442_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__o21a_1
XFILLER_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13475_ net1693 net320 net423 VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__mux2_1
X_10687_ cpuregs\[20\]\[9\] cpuregs\[21\]\[9\] net671 VGND VGND VPWR VPWR _05378_
+ sky130_fd_sc_hd__mux2_1
X_15214_ clknet_leaf_99_clk _01563_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.instr_mulh
+ sky130_fd_sc_hd__dfxtp_1
X_12426_ net1218 genblk1.genblk1.pcpi_mul.mul_counter\[0\] genblk1.genblk1.pcpi_mul.mul_counter\[1\]
+ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__or3_1
XFILLER_127_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15145_ clknet_leaf_49_clk _01497_ VGND VGND VPWR VPWR cpuregs\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12357_ latched_rd\[0\] _04290_ latched_rd\[1\] VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__and3b_1
XFILLER_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output81_A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11591__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_947 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11308_ net785 _05972_ _05981_ net778 VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__o211a_1
X_15076_ clknet_leaf_103_clk net2368 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08322__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12288_ decoded_imm\[29\] net739 VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14027_ clknet_leaf_68_clk _00481_ VGND VGND VPWR VPWR cpuregs\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11239_ cpuregs\[1\]\[24\] net551 _05914_ net807 net836 VGND VGND VPWR VPWR _05915_
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06780_ mem_rdata_q\[14\] VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__inv_2
XFILLER_48_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09153__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14929_ clknet_leaf_179_clk _01281_ VGND VGND VPWR VPWR cpuregs\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_08450_ _03850_ _03851_ net768 VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__mux2_2
XFILLER_63_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07401_ net358 _02932_ _02937_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__o21bai_2
X_08381_ reg_pc\[12\] _03788_ reg_pc\[13\] VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__a21oi_1
X_07332_ count_cycle\[12\] net972 VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_98_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07263_ _02806_ _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__nand2_1
X_09002_ net408 net2081 net516 VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__mux2_1
X_07194_ net1062 _02739_ _02743_ net1082 _02742_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__a221o_1
XFILLER_118_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11582__B2 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09328__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13358__B net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11159__A net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout502 net503 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_8
X_09904_ net2564 net881 _04683_ net851 VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__a22o_1
XANTENNA__14531__Q decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout513 net515 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__buf_4
XANTENNA__12830__X _02118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout524 _03774_ VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__buf_2
XANTENNA__11334__A1 net840 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout535 _06240_ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1207_A _02378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout546 _03741_ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A mem_rdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout557 _02133_ VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__buf_2
X_09835_ _04617_ _04619_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__nor2_1
Xfanout568 net570 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout579 _03753_ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout667_A net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13374__A net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09766_ decoded_imm_j\[12\] _04433_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__or2_1
X_06978_ net1119 _02553_ genblk2.pcpi_div.dividend\[9\] VGND VGND VPWR VPWR _02555_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__09063__S net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08717_ genblk1.genblk1.pcpi_mul.next_rs2\[37\] net1099 _04072_ _04074_ VGND VGND
+ VPWR VPWR _04075_ sky130_fd_sc_hd__a22o_1
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09697_ decoded_imm_j\[6\] _04427_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout834_A _03137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout455_X net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout1197_X net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08648_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ genblk1.genblk1.pcpi_mul.next_rs2\[16\] net1094 genblk1.genblk1.pcpi_mul.rd\[15\]
+ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__a21o_1
XANTENNA__11622__A mem_rdata_q\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10610_ cpuregs\[17\]\[7\] net626 net608 _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__o211a_1
XFILLER_167_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11590_ net2922 net563 _06185_ _06192_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__a22o_1
XFILLER_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10541_ cpuregs\[16\]\[5\] net676 VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__or2_1
XANTENNA__10238__A decoded_imm\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13260_ reg_pc\[7\] net564 _02183_ _02184_ net391 VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout991_X net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10472_ cpuregs\[6\]\[1\] cpuregs\[7\]\[1\] net686 VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__mux2_1
XANTENNA__11768__S net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12211_ genblk2.pcpi_div.quotient_msk\[19\] net270 net2812 VGND VGND VPWR VPWR _06598_
+ sky130_fd_sc_hd__a21oi_1
X_13191_ net2154 net303 net430 VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__mux2_1
XFILLER_109_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09238__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12142_ genblk2.pcpi_div.quotient_msk\[1\] net382 net372 net2750 VGND VGND VPWR VPWR
+ _01043_ sky130_fd_sc_hd__a22o_1
XANTENNA__07241__A2 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08142__S _02364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07266__B _02799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12073_ _06273_ _06275_ _06520_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__or3_1
XANTENNA__11325__A1 net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11024_ cpuregs\[17\]\[18\] net618 net603 _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__o211a_1
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12599__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_144_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07282__A net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input16_X net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11628__A2 net738 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12975_ net1739 net525 net447 VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__mux2_1
XANTENNA_output217_A net1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14714_ clknet_leaf_153_clk _01099_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10836__B1 net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11926_ genblk2.pcpi_div.divisor\[35\] genblk2.pcpi_div.divisor\[34\] genblk2.pcpi_div.divisor\[33\]
+ genblk2.pcpi_div.divisor\[32\] VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__or4_1
XANTENNA__11617__A_N mem_rdata_q\[27\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14645_ clknet_leaf_161_clk _01030_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_11857_ _06310_ _06312_ _06326_ _06311_ _06308_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__a311o_1
XFILLER_82_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10808_ cpuregs\[4\]\[13\] net653 VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__or2_1
XFILLER_158_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14576_ clknet_leaf_88_clk _00962_ VGND VGND VPWR VPWR is_alu_reg_reg sky130_fd_sc_hd__dfxtp_1
XANTENNA__13250__A1 net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11788_ genblk2.pcpi_div.divisor\[31\] genblk2.pcpi_div.dividend\[31\] VGND VGND
+ VPWR VPWR _06259_ sky130_fd_sc_hd__and2b_1
X_13527_ net540 net1800 net415 VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__mux2_1
XFILLER_158_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10739_ cpuregs\[25\]\[11\] net625 net607 _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__o211a_1
XANTENNA__08009__A1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13458_ net1431 net575 net423 VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12409_ net335 net1977 net471 VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput105 net105 VGND VGND VPWR VPWR mem_la_wdata[17] sky130_fd_sc_hd__buf_2
X_13389_ net569 _05890_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__nor2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput116 net116 VGND VGND VPWR VPWR mem_la_wdata[27] sky130_fd_sc_hd__buf_2
XANTENNA__09148__S net500 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput127 net127 VGND VGND VPWR VPWR mem_la_wdata[8] sky130_fd_sc_hd__buf_2
X_15128_ clknet_leaf_192_clk _01480_ VGND VGND VPWR VPWR cpuregs\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xoutput138 net138 VGND VGND VPWR VPWR mem_wdata[12] sky130_fd_sc_hd__buf_2
Xoutput149 net149 VGND VGND VPWR VPWR mem_wdata[22] sky130_fd_sc_hd__buf_2
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15059_ clknet_leaf_104_clk _01411_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_07950_ net1047 net1178 net932 VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__and3_1
XANTENNA__08987__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11316__A1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06901_ is_sll_srl_sra is_sb_sh_sw _02436_ net1087 VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_71_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07881_ net1159 _02409_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__or2_1
XANTENNA__10524__C1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09620_ _03808_ reg_next_pc\[16\] net922 VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__mux2_1
X_06832_ _02379_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__or2_1
XANTENNA__07904__B net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07940__B1 net969 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09551_ net3051 _04395_ net1230 VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06763_ reg_pc\[2\] VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__inv_2
X_08502_ _03891_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__nand2_1
X_09482_ net2935 _04350_ net1239 VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08433_ reg_pc\[23\] _03834_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__xor2_1
XANTENNA__10757__S net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13133__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08248__A1 net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08364_ net409 net2182 net529 VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07315_ genblk1.genblk1.pcpi_mul.pcpi_rd\[11\] genblk2.pcpi_div.pcpi_rd\[11\] net1110
+ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__mux2_1
XANTENNA__14526__Q decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12972__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08295_ net1004 _03731_ net982 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__mux2_2
XANTENNA_fanout415_A _02357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_A net259 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07246_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__inv_2
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07208__C1 net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07177_ _02710_ _02726_ _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__o21a_1
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09058__S net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12752__B1 net918 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout784_A _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10505__B _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout310 net311 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1112_X net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout321 _03826_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_1
Xfanout332 net333 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout343 net344 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input8_X net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout354 net355 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout951_A net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout365 net370 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout376 _06234_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_4
XFILLER_74_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09818_ decoded_imm_j\[16\] _04437_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__nand2_1
Xfanout387 net388 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout398 _04887_ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__buf_2
XFILLER_59_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07814__B net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09749_ _04431_ _04529_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10240__B net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_X net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12760_ net1216 net1450 net918 net993 VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__a22o_1
XFILLER_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11711_ net1968 net295 net376 VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__mux2_1
X_12691_ net1211 net2952 net900 net2955 net713 VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__a221o_1
XANTENNA__13043__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14430_ clknet_leaf_67_clk alu_out\[30\] VGND VGND VPWR VPWR alu_out_q\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08239__A1 net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11642_ decoded_imm_j\[6\] net19 net545 VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__mux2_1
XANTENNA__13232__A1 net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09987__A1 net1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14361_ clknet_leaf_131_clk _00782_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_2
XFILLER_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11573_ instr_lh net741 _06181_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__a22o_1
XFILLER_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 mem_rdata[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13312_ _04922_ _04984_ _02229_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__o21a_1
Xinput29 mem_rdata[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10524_ net815 _05216_ _05218_ net829 VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__o211a_1
XFILLER_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14292_ clknet_leaf_128_clk _00746_ VGND VGND VPWR VPWR count_cycle\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09739__A1 net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13279__A net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13243_ reg_pc\[5\] net565 _02167_ _02169_ net391 VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__a2111oi_1
XFILLER_136_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10455_ cpuregs\[19\]\[0\] net635 net600 _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__o211a_1
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13174_ net1540 net520 net427 VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__mux2_1
X_10386_ genblk2.pcpi_div.quotient_msk\[23\] genblk2.pcpi_div.quotient_msk\[22\] genblk2.pcpi_div.quotient_msk\[21\]
+ genblk2.pcpi_div.quotient_msk\[20\] VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12125_ genblk2.pcpi_div.dividend\[29\] _06566_ net274 VGND VGND VPWR VPWR _01038_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12056_ genblk2.pcpi_div.dividend\[19\] net269 _06507_ VGND VGND VPWR VPWR _01028_
+ sky130_fd_sc_hd__o21ba_1
X_11007_ cpuregs\[9\]\[18\] net618 net603 _05688_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__o211a_1
XFILLER_65_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11961__S net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10809__B1 net812 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12958_ net309 net2164 net451 VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__mux2_1
XFILLER_46_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10285__A1 _04987_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11909_ _06267_ _06378_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__nor2_1
XFILLER_34_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10577__S net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12889_ mem_rdata_q\[26\] net19 net964 VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__mux2_1
XFILLER_61_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14628_ clknet_leaf_135_clk _01013_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12026__A2 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09978__B2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14559_ clknet_leaf_11_clk _00945_ VGND VGND VPWR VPWR cpuregs\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11785__A1 net1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07100_ genblk2.pcpi_div.quotient\[25\] _02651_ net1122 VGND VGND VPWR VPWR _02660_
+ sky130_fd_sc_hd__o21a_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08080_ _03341_ _03576_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__nor2_1
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07453__A2 net1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07031_ net1115 genblk2.pcpi_div.quotient\[16\] _02599_ net950 VGND VGND VPWR VPWR
+ _02601_ sky130_fd_sc_hd__a31o_1
XFILLER_161_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11537__A1 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07205__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15177__Q mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08982_ genblk1.genblk1.pcpi_mul.rd\[29\] genblk1.genblk1.pcpi_mul.rd\[61\] net956
+ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09606__S net927 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07933_ _03393_ _03395_ _03450_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__or3b_1
XANTENNA__13128__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09902__A1 net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07864_ _03271_ _03294_ _03380_ _03381_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__or4bb_1
XANTENNA__10512__A2 decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09603_ reg_pc\[7\] net882 _04428_ net846 VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__a22o_1
X_06815_ net1133 net1141 net1137 VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__nor3_1
X_07795_ net256 net994 VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__or2_1
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11724__X _06240_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09534_ count_instr\[44\] count_instr\[43\] _04382_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12265__A2 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09341__S net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09465_ _04340_ _04341_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12670__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08416_ reg_out\[20\] alu_out_q\[20\] net1155 VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09396_ net196 net193 net197 net198 VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_35_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08347_ _03767_ _03768_ net766 VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1062_X net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_X net418 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07649__X _03170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08278_ reg_out\[16\] reg_next_pc\[16\] net922 VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__mux2_1
XFILLER_165_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07229_ reg_pc\[6\] decoded_imm\[6\] VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__or2_1
XFILLER_164_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10240_ decoded_imm\[5\] net1040 VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__nor2_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout787_X net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10235__B net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10171_ count_cycle\[61\] count_cycle\[62\] count_cycle\[63\] _04873_ net1209 VGND
+ VGND VPWR VPWR _04878_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_163_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07384__X _06722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1105 net1108 VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__buf_2
Xfanout1116 net1117 VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__buf_1
XFILLER_121_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1127 net1128 VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__buf_2
XANTENNA__08420__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1138 instr_rdinstr VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout954_X net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1149 instr_jal VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13038__S net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13930_ clknet_leaf_46_clk _00384_ VGND VGND VPWR VPWR cpuregs\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10251__A decoded_imm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13861_ clknet_leaf_23_clk _00315_ VGND VGND VPWR VPWR cpuregs\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_190_clk_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15600_ clknet_leaf_190_clk _01936_ VGND VGND VPWR VPWR cpuregs\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12812_ net346 net2200 net463 VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__mux2_1
XFILLER_62_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13453__A1 net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12256__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13792_ clknet_leaf_8_clk _00246_ VGND VGND VPWR VPWR cpuregs\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09251__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15531_ clknet_leaf_22_clk _01867_ VGND VGND VPWR VPWR cpuregs\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12743_ net1191 genblk1.genblk1.pcpi_mul.next_rs1\[20\] net2105 net897 _02105_ VGND
+ VGND VPWR VPWR _01391_ sky130_fd_sc_hd__a221o_1
XFILLER_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12178__A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15462_ clknet_leaf_85_clk _00014_ VGND VGND VPWR VPWR mem_wordsize\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12674_ net1201 genblk1.genblk1.pcpi_mul.next_rs2\[39\] net892 net3035 net712 VGND
+ VGND VPWR VPWR _01344_ sky130_fd_sc_hd__a221o_1
X_14413_ clknet_leaf_177_clk alu_out\[13\] VGND VGND VPWR VPWR alu_out_q\[13\] sky130_fd_sc_hd__dfxtp_1
X_11625_ _06207_ _06213_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_139_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ clknet_leaf_71_clk _01732_ VGND VGND VPWR VPWR cpuregs\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13501__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14344_ clknet_leaf_82_clk _06732_ VGND VGND VPWR VPWR reg_out\[24\] sky130_fd_sc_hd__dfxtp_1
X_11556_ net1998 net563 _06175_ _06178_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__a22o_1
XFILLER_156_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10507_ net1179 net860 _05204_ _05205_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__o22a_1
X_14275_ clknet_leaf_97_clk _00729_ VGND VGND VPWR VPWR count_cycle\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11487_ _03739_ _06153_ _06154_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__o21a_1
XANTENNA__11021__S net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13226_ _02475_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__or2_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10438_ cpuregs\[2\]\[0\] net685 VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__or2_1
XFILLER_124_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10860__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13157_ net2324 net305 net433 VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__mux2_1
XFILLER_112_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10369_ net774 _05066_ _05074_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_143_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12108_ genblk2.pcpi_div.dividend\[26\] _06552_ net273 VGND VGND VPWR VPWR _01035_
+ sky130_fd_sc_hd__mux2_1
X_13088_ net313 net2062 net441 VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12039_ net721 _06492_ net1016 VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09896__B1 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_158_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11691__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07580_ net22 net938 net937 VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12247__A2 net379 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09161__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11455__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15729_ net119 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09250_ net1385 net320 net488 VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__mux2_1
XFILLER_167_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08201_ _03449_ _03688_ net990 VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09181_ net335 net2151 net497 VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__mux2_1
XANTENNA__09397__A net267 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08132_ _03331_ _03627_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__nand2_1
XANTENNA__08623__A1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12535__B net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08063_ _03379_ _03436_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__and2_1
XFILLER_107_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10981__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07014_ genblk2.pcpi_div.dividend\[14\] net1115 _02584_ net947 VGND VGND VPWR VPWR
+ _02586_ sky130_fd_sc_hd__a31o_1
XFILLER_162_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1022_A net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10733__A2 _05421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09336__S net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08965_ net2656 _04259_ net945 VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout482_A _04291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07916_ net1164 _02405_ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__o21a_1
X_08896_ _03914_ _03916_ _03913_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__a21bo_1
XFILLER_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07847_ _03360_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout747_A _06163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07778_ net253 net1000 VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__or2_1
XANTENNA__12238__A2 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09071__S net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09517_ count_instr\[37\] _04372_ count_instr\[38\] VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout914_A net919 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_X net535 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09448_ count_instr\[14\] count_instr\[13\] count_instr\[12\] _04325_ VGND VGND VPWR
+ VPWR _04330_ sky130_fd_sc_hd__and4_1
XANTENNA__13199__B1 net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09379_ net1813 net339 net399 VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout702_X net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11749__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11410_ net808 _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__or2_1
XANTENNA__07379__X _02917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12390_ latched_rd\[4\] latched_rd\[3\] latched_rd\[2\] VGND VGND VPWR VPWR _06663_
+ sky130_fd_sc_hd__or3b_1
XANTENNA__08415__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11341_ cpuregs\[10\]\[27\] net693 VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__or2_1
XFILLER_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10246__A net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14060_ clknet_leaf_54_clk _00514_ VGND VGND VPWR VPWR cpuregs\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11272_ cpuregs\[22\]\[25\] cpuregs\[23\]\[25\] net705 VGND VGND VPWR VPWR _05947_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13011_ net521 net2447 net443 VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__mux2_1
X_10223_ decoded_imm\[11\] net1028 VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__nand2_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12461__A net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09246__S net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10154_ count_cycle\[56\] count_cycle\[57\] VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__and2_1
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ clknet_leaf_147_clk _01314_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10085_ count_cycle\[32\] _04821_ net1207 VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__a21oi_1
Xhold7 cpuregs\[0\]\[17\] VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13913_ clknet_leaf_5_clk _00367_ VGND VGND VPWR VPWR cpuregs\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14893_ clknet_leaf_140_clk _01245_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13844_ clknet_leaf_178_clk _00298_ VGND VGND VPWR VPWR cpuregs\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12400__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12229__A2 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13775_ clknet_leaf_47_clk _00229_ VGND VGND VPWR VPWR cpuregs\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10987_ cpuregs\[25\]\[17\] net617 net603 _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__o211a_1
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12726_ _02406_ net911 VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__nor2_1
XFILLER_71_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15514_ clknet_leaf_78_clk _01850_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dfxtp_1
XANTENNA__07656__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15445_ clknet_leaf_9_clk _01784_ VGND VGND VPWR VPWR cpuregs\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12657_ _02397_ net913 VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_61_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ net3032 net561 net732 _06201_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__a22o_1
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15376_ clknet_leaf_2_clk _01715_ VGND VGND VPWR VPWR cpuregs\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07408__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12588_ net341 net2223 net467 VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__mux2_1
XANTENNA__08325__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14327_ clknet_leaf_174_clk _06745_ VGND VGND VPWR VPWR reg_out\[7\] sky130_fd_sc_hd__dfxtp_1
X_11539_ net1 net12 VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__nand2_1
Xhold407 cpuregs\[23\]\[25\] VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10963__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold418 genblk1.genblk1.pcpi_mul.next_rs1\[11\] VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 cpuregs\[24\]\[29\] VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ clknet_leaf_128_clk _00712_ VGND VGND VPWR VPWR count_cycle\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__06921__X _02509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11686__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13209_ net1065 net1040 net755 net557 VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__a31o_1
XANTENNA__10590__S net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14189_ clknet_leaf_101_clk _00643_ VGND VGND VPWR VPWR count_instr\[60\] sky130_fd_sc_hd__dfxtp_1
Xfanout909 net910 VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09156__S net503 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13114__A0 net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08750_ _04100_ _04102_ _04095_ _04098_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__a211o_1
Xhold1107 genblk1.genblk1.pcpi_mul.next_rs1\[13\] VGND VGND VPWR VPWR net2421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 genblk1.genblk1.pcpi_mul.next_rs1\[37\] VGND VGND VPWR VPWR net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08995__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1129 genblk1.genblk1.pcpi_mul.next_rs1\[54\] VGND VGND VPWR VPWR net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ cpuregs\[16\]\[3\] net676 VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__or2_1
X_08681_ net905 _04042_ _04044_ net2696 net1218 VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__a32o_1
XANTENNA__07344__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07344__B2 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07632_ net824 net810 VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__nor2_2
XANTENNA__13417__A1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07563_ reg_pc\[28\] decoded_imm\[28\] VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__nand2_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11979__A1 net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09302_ net1449 net573 net482 VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__mux2_1
X_07494_ net16 net938 net936 VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09233_ net1845 net577 net489 VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__mux2_1
XANTENNA__13141__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A _03818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09164_ net588 net1900 net498 VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__mux2_1
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08235__S net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14534__Q is_lui_auipc_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08115_ _03348_ _03437_ _03401_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__o21a_1
XANTENNA__12980__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09095_ net2538 net583 net506 VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1237_A net1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08046_ net967 _03286_ _03288_ net928 _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__a221o_1
Xhold930 cpuregs\[21\]\[30\] VGND VGND VPWR VPWR net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 cpuregs\[15\]\[0\] VGND VGND VPWR VPWR net2255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold952 cpuregs\[1\]\[10\] VGND VGND VPWR VPWR net2266 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold963 cpuregs\[10\]\[1\] VGND VGND VPWR VPWR net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12281__A _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold974 cpuregs\[17\]\[3\] VGND VGND VPWR VPWR net2288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1025_X net1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold985 cpuregs\[9\]\[7\] VGND VGND VPWR VPWR net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 cpuregs\[11\]\[5\] VGND VGND VPWR VPWR net2310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09066__S net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09997_ net849 _04766_ _04767_ net879 net2512 VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__a32o_1
XFILLER_135_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout864_A net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_X net485 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08948_ genblk1.genblk1.pcpi_mul.rd\[12\] genblk1.genblk1.pcpi_mul.rd\[44\] net954
+ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1630 genblk2.pcpi_div.quotient\[14\] VGND VGND VPWR VPWR net2944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1641 genblk1.genblk1.pcpi_mul.next_rs2\[55\] VGND VGND VPWR VPWR net2955 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_48_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08879_ _04210_ _04211_ _04205_ _04208_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__a211o_1
Xhold1652 genblk2.pcpi_div.quotient_msk\[4\] VGND VGND VPWR VPWR net2966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07335__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1663 genblk1.genblk1.pcpi_mul.next_rs2\[52\] VGND VGND VPWR VPWR net2977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1674 count_cycle\[16\] VGND VGND VPWR VPWR net2988 sky130_fd_sc_hd__dlygate4sd3_1
X_10910_ cpuregs\[19\]\[15\] net617 net589 VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__o21a_1
XFILLER_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1685 genblk2.pcpi_div.quotient\[1\] VGND VGND VPWR VPWR net2999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1696 genblk2.pcpi_div.dividend\[5\] VGND VGND VPWR VPWR net3010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11890_ _06286_ _06290_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__nand2_1
XFILLER_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07886__A2 _02410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10841_ net1075 decoded_imm\[13\] VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__or2_1
XFILLER_72_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_X net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07099__B1 net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13560_ net540 net2439 net411 VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__mux2_1
X_10772_ cpuregs\[30\]\[12\] cpuregs\[31\]\[12\] net650 VGND VGND VPWR VPWR _05460_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12511_ net2543 net387 _02003_ _02004_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__a22o_1
XFILLER_157_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10642__A1 net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13491_ net1771 net575 net419 VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13051__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15230_ clknet_leaf_22_clk _01571_ VGND VGND VPWR VPWR cpuregs\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ genblk2.pcpi_div.divisor\[33\] _06676_ net868 VGND VGND VPWR VPWR _06677_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_57_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15161_ clknet_leaf_65_clk _01510_ VGND VGND VPWR VPWR mem_rdata_q\[12\] sky130_fd_sc_hd__dfxtp_4
X_12373_ net1383 net340 net360 VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__mux2_1
XFILLER_126_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14112_ clknet_leaf_2_clk _00566_ VGND VGND VPWR VPWR cpuregs\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11324_ net836 _05993_ _05995_ _05997_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__a211o_1
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15092_ clknet_leaf_181_clk _01444_ VGND VGND VPWR VPWR cpuregs\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14043_ clknet_leaf_195_clk _00497_ VGND VGND VPWR VPWR cpuregs\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13287__A net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11255_ cpuregs\[4\]\[25\] cpuregs\[5\]\[25\] net702 VGND VGND VPWR VPWR _05930_
+ sky130_fd_sc_hd__mux2_1
X_10206_ decoded_imm\[21\] net216 VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__and2_1
X_11186_ cpuregs\[26\]\[23\] net685 VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__or2_1
XFILLER_122_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07574__A1 net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output247_A net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10137_ count_cycle\[51\] _04854_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_66_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11658__A0 decoded_imm_j\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10068_ count_cycle\[26\] _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14945_ clknet_leaf_36_clk _01297_ VGND VGND VPWR VPWR cpuregs\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11122__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14876_ clknet_leaf_38_clk _01228_ VGND VGND VPWR VPWR cpuregs\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13827_ clknet_leaf_13_clk _00281_ VGND VGND VPWR VPWR cpuregs\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13758_ clknet_leaf_11_clk _00212_ VGND VGND VPWR VPWR cpuregs\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12709_ net1339 net884 _02088_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__a21o_1
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_75_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13689_ clknet_leaf_107_clk _00143_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11270__A net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15428_ clknet_leaf_38_clk _01767_ VGND VGND VPWR VPWR cpuregs\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15359_ clknet_leaf_55_clk _01699_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
XFILLER_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 cpuregs\[30\]\[15\] VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold215 cpuregs\[22\]\[8\] VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 cpuregs\[13\]\[8\] VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold237 cpuregs\[14\]\[23\] VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 cpuregs\[28\]\[26\] VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13335__B1 net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09920_ _04445_ _04691_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__nor2_1
Xhold259 cpuregs\[23\]\[18\] VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07014__B1 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout706 net707 VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkbuf_4
Xfanout717 net718 VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__buf_2
X_09851_ _04438_ _04611_ _04439_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_111_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout728 _06244_ VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_84_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 net742 VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlymetal6s2s_1
X_08802_ _04144_ _04146_ _04139_ _04142_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__a211o_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09782_ _04526_ _04536_ _04568_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06994_ genblk2.pcpi_div.dividend\[10\] genblk2.pcpi_div.dividend\[9\] _02553_ VGND
+ VGND VPWR VPWR _02569_ sky130_fd_sc_hd__or3_1
XANTENNA__09614__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08733_ net892 _04086_ _04088_ net2691 net1201 VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__a32o_1
XFILLER_67_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11113__A2 net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _03873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13136__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12310__B2 mem_rdata_q\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08664_ genblk1.genblk1.pcpi_mul.rd\[28\] genblk1.genblk1.pcpi_mul.rdx\[28\] VGND
+ VGND VPWR VPWR _04030_ sky130_fd_sc_hd__or2_1
X_07615_ net986 decoded_imm_j\[2\] _03135_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__o21ai_2
XANTENNA__14529__Q decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12975__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08595_ _03963_ _03966_ _03968_ _03970_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout445_A net446 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07546_ reg_pc\[27\] decoded_imm\[27\] VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__nand2_1
XFILLER_35_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ _03006_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout612_A net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09216_ net2190 net326 net494 VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__mux2_1
XFILLER_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09147_ net1764 net338 net501 VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout400_X net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_X net1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07253__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09078_ net1514 net332 net508 VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__mux2_1
XFILLER_136_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout981_A net983 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13326__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08029_ _03360_ _03530_ _03411_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__a21o_1
Xhold760 cpuregs\[6\]\[1\] VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 cpuregs\[25\]\[22\] VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 cpuregs\[27\]\[30\] VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ cpuregs\[12\]\[19\] cpuregs\[13\]\[19\] net680 VGND VGND VPWR VPWR _05721_
+ sky130_fd_sc_hd__mux2_1
Xhold793 genblk1.genblk1.pcpi_mul.next_rs1\[44\] VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout867_X net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10243__B net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ net1442 net310 net449 VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__mux2_1
Xhold1460 count_instr\[18\] VGND VGND VPWR VPWR net2774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13046__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12301__A1 mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1471 genblk2.pcpi_div.quotient_msk\[15\] VGND VGND VPWR VPWR net2785 sky130_fd_sc_hd__dlygate4sd3_1
X_14730_ clknet_leaf_170_clk _01115_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11942_ _06411_ _06410_ _06408_ net866 VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__a2bb2o_1
Xhold1482 count_instr\[39\] VGND VGND VPWR VPWR net2796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 _06607_ VGND VGND VPWR VPWR net2807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14661_ clknet_leaf_152_clk net2530 VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _06305_ _06342_ _06306_ _06333_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__or4b_1
XFILLER_33_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13612_ clknet_leaf_0_clk _00067_ VGND VGND VPWR VPWR cpuregs\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_10824_ cpuregs\[30\]\[13\] cpuregs\[31\]\[13\] net651 VGND VGND VPWR VPWR _05511_
+ sky130_fd_sc_hd__mux2_1
X_14592_ clknet_leaf_159_clk _00978_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11361__Y _06034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13543_ net312 net1878 net417 VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__mux2_1
X_10755_ cpuregs\[1\]\[11\] net549 _05443_ net796 net823 VGND VGND VPWR VPWR _05444_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12186__A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13474_ net1779 net324 net425 VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__mux2_1
X_10686_ net830 _05372_ _05374_ _05376_ net789 VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__a2111o_1
X_15213_ clknet_leaf_98_clk _01562_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.instr_mulhsu
+ sky130_fd_sc_hd__dfxtp_1
X_12425_ net1218 genblk1.genblk1.pcpi_mul.mul_counter\[0\] net3012 VGND VGND VPWR
+ VPWR _06665_ sky130_fd_sc_hd__o21a_1
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08036__A2 net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15144_ clknet_leaf_53_clk _01496_ VGND VGND VPWR VPWR cpuregs\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12356_ net910 _06659_ _06660_ _06661_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__a31o_1
XFILLER_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11591__A2 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11307_ net794 _05976_ _05978_ _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__or4_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15075_ clknet_leaf_103_clk _01427_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12287_ decoded_imm\[30\] net739 net559 mem_rdata_q\[30\] net532 VGND VGND VPWR VPWR
+ _01144_ sky130_fd_sc_hd__a221o_1
XANTENNA__12125__S net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output74_A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14026_ clknet_leaf_45_clk _00480_ VGND VGND VPWR VPWR cpuregs\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11238_ cpuregs\[2\]\[24\] cpuregs\[3\]\[24\] net699 VGND VGND VPWR VPWR _05914_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11169_ cpuregs\[20\]\[22\] cpuregs\[21\]\[22\] net682 VGND VGND VPWR VPWR _05847_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08398__X _03810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14928_ clknet_leaf_23_clk _01280_ VGND VGND VPWR VPWR cpuregs\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10854__A1 net812 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14859_ clknet_leaf_23_clk _01211_ VGND VGND VPWR VPWR cpuregs\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07400_ net1065 net1018 _02936_ net1079 _02935_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__a221o_1
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ reg_out\[13\] alu_out_q\[13\] net1153 VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__mux2_1
X_07331_ net1140 count_cycle\[44\] net977 _02871_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__a211o_1
XANTENNA__12096__A net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_X clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07483__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07262_ reg_pc\[8\] decoded_imm\[8\] VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__nand2_1
XFILLER_149_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09001_ net521 net1685 net516 VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__mux2_1
X_07193_ genblk1.genblk1.pcpi_mul.pcpi_rd\[3\] genblk2.pcpi_div.pcpi_rd\[3\] net1111
+ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__mux2_1
XANTENNA__10047__C _04791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11031__A1 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14812__Q decoded_imm\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12035__S net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09903_ _04443_ _04682_ net1184 VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__mux2_1
Xfanout503 _04284_ VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_4_9_0_clk_X clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout514 net515 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_4
XANTENNA__07538__A1 genblk2.pcpi_div.pcpi_rd\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout525 _03774_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__buf_1
Xfanout536 _06240_ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__buf_4
XANTENNA_fanout395_A net398 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout547 net548 VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11727__X _06242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09834_ _04522_ _04569_ _04570_ _04618_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__and4_1
XANTENNA__10542__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout558 _02133_ VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__buf_2
Xfanout569 net570 VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09344__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09765_ net845 _04554_ _04555_ net875 net2446 VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__a32o_1
XANTENNA__13374__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06977_ genblk2.pcpi_div.dividend\[9\] net1119 _02553_ VGND VGND VPWR VPWR _02554_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11098__A1 net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08716_ genblk1.genblk1.pcpi_mul.rd\[36\] genblk1.genblk1.pcpi_mul.rdx\[36\] VGND
+ VGND VPWR VPWR _04074_ sky130_fd_sc_hd__or2_1
XFILLER_55_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09696_ _04491_ _04492_ net2821 net878 VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__a2bb2o_1
X_08647_ _04007_ _04010_ _04012_ _04014_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_124_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout827_A net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13390__A net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08578_ genblk1.genblk1.pcpi_mul.rd\[15\] genblk1.genblk1.pcpi_mul.next_rs2\[16\]
+ net1094 VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__nand3_1
XANTENNA__12718__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11622__B mem_rdata_q\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07529_ net359 _03051_ _03056_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout615_X net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10540_ _05233_ _05234_ net802 VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__mux2_1
XFILLER_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10238__B net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10471_ net1181 net860 _05169_ _05170_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12734__A _02408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ net748 _06597_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__nor2_1
XANTENNA__07828__A net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13190_ net2369 net305 net429 VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__mux2_1
XFILLER_108_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout984_X net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12141_ net2602 net385 net372 genblk2.pcpi_div.quotient_msk\[1\] VGND VGND VPWR VPWR
+ _01042_ sky130_fd_sc_hd__a22o_1
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12072_ _06275_ _06520_ _06273_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__o21ai_1
Xhold590 cpuregs\[16\]\[19\] VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ cpuregs\[16\]\[18\] net647 VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__or2_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09254__S net491 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ net1497 net539 net447 VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__mux2_1
XFILLER_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07850__X _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1290 genblk1.genblk1.pcpi_mul.rd\[4\] VGND VGND VPWR VPWR net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_14713_ clknet_leaf_154_clk _01098_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_11925_ genblk2.pcpi_div.divisor\[55\] genblk2.pcpi_div.divisor\[54\] genblk2.pcpi_div.divisor\[53\]
+ genblk2.pcpi_div.divisor\[52\] VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__or4_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13504__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14644_ clknet_leaf_161_clk _01029_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_11856_ _06312_ _06326_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__and2_1
XFILLER_72_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10807_ cpuregs\[6\]\[13\] cpuregs\[7\]\[13\] net653 VGND VGND VPWR VPWR _05494_
+ sky130_fd_sc_hd__mux2_1
X_14575_ clknet_leaf_89_clk _00961_ VGND VGND VPWR VPWR is_alu_reg_imm sky130_fd_sc_hd__dfxtp_2
X_11787_ net867 _05095_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__nor2_1
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11261__A1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10738_ cpuregs\[24\]\[11\] net664 VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__or2_1
X_13526_ net541 net2075 net415 VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__mux2_1
XFILLER_158_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13457_ net1399 net579 net426 VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__mux2_1
X_10669_ cpuregs\[14\]\[9\] cpuregs\[15\]\[9\] net667 VGND VGND VPWR VPWR _05360_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07217__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12408_ net338 net1756 net472 VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__mux2_1
XANTENNA__07297__X _02840_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08333__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13388_ net961 _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__nor2_1
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput106 net106 VGND VGND VPWR VPWR mem_la_wdata[18] sky130_fd_sc_hd__buf_2
Xoutput117 net117 VGND VGND VPWR VPWR mem_la_wdata[28] sky130_fd_sc_hd__buf_2
X_15127_ clknet_leaf_195_clk _01479_ VGND VGND VPWR VPWR cpuregs\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xoutput128 net128 VGND VGND VPWR VPWR mem_la_wdata[9] sky130_fd_sc_hd__buf_2
X_12339_ decoded_imm\[5\] net735 _06643_ mem_rdata_q\[25\] _06649_ VGND VGND VPWR
+ VPWR _01169_ sky130_fd_sc_hd__a221o_1
Xoutput139 net139 VGND VGND VPWR VPWR mem_wdata[13] sky130_fd_sc_hd__buf_2
XFILLER_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15058_ clknet_leaf_105_clk net2290 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11694__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06900_ net1232 _02439_ _02440_ _02445_ _02495_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__a41o_1
X_14009_ clknet_leaf_191_clk _00463_ VGND VGND VPWR VPWR cpuregs\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07744__Y _03263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07880_ net1161 _02407_ _03347_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__o31a_1
XFILLER_96_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09164__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06831_ _00003_ net975 _02422_ _02435_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__or4_2
X_09550_ count_instr\[50\] _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__and2_1
X_06762_ net1089 VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__inv_2
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08501_ genblk1.genblk1.pcpi_mul.next_rs2\[4\] net1098 genblk1.genblk1.pcpi_mul.rd\[3\]
+ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__a21o_1
X_09481_ count_instr\[25\] count_instr\[24\] _04344_ _04348_ VGND VGND VPWR VPWR _04352_
+ sky130_fd_sc_hd__and4_1
XFILLER_36_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11723__A net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08432_ reg_out\[23\] alu_out_q\[23\] net1155 VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__mux2_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08363_ _03778_ _03781_ net766 VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__mux2_1
XANTENNA__14807__Q decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08248__A2 net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07314_ count_cycle\[11\] net971 net841 _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__o211a_1
XANTENNA__11252__A1 net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08294_ reg_out\[24\] reg_next_pc\[24\] net925 VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__mux2_1
XFILLER_165_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07245_ reg_pc\[7\] decoded_imm\[7\] VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__and2_1
XANTENNA__10773__S net797 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_A net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09339__S net475 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07208__B1 _02756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07176_ _02710_ _02726_ net991 VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__a21oi_1
XFILLER_106_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14542__Q is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12752__A1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12752__B2 net1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07367__B decoded_imm\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout300 _03852_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_1
Xfanout311 _03839_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout398_X net398 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout322 _03826_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_2
Xfanout333 _03815_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout344 net345 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__buf_1
Xfanout355 net357 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08479__A genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09074__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout366 net370 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout377 net384 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_4
X_09817_ net2617 net876 _04599_ _04603_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__a22o_1
Xfanout388 net390 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_161_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout399 _04293_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__buf_4
XANTENNA_fanout565_X net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A _00015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09748_ _04529_ _04431_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__and2b_1
XFILLER_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09679_ _04473_ _04474_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__and3_1
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08485__Y _03879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11710_ net2011 net300 net375 VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__mux2_1
X_12690_ net1210 net2955 net900 genblk1.genblk1.pcpi_mul.next_rs2\[54\] net713 VGND
+ VGND VPWR VPWR _01360_ sky130_fd_sc_hd__a221o_1
XFILLER_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08418__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11641_ net3064 net18 net545 VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__mux2_1
XFILLER_70_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14360_ clknet_leaf_80_clk _00781_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_2
X_11572_ net3036 net740 _06176_ is_lb_lh_lw_lbu_lhu VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__a22o_1
XFILLER_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13311_ _04922_ _04984_ net960 VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__a21oi_1
Xinput19 mem_rdata[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
X_10523_ net801 _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__or2_1
XFILLER_167_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14291_ clknet_leaf_128_clk _00745_ VGND VGND VPWR VPWR count_cycle\[36\] sky130_fd_sc_hd__dfxtp_1
X_13242_ net1038 net758 _02168_ _02474_ net1063 VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09249__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10454_ cpuregs\[18\]\[0\] net686 VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__or2_1
XFILLER_164_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12743__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12743__B2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07277__B decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13173_ net2116 net526 net427 VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__mux2_1
X_10385_ genblk2.pcpi_div.quotient_msk\[31\] genblk2.pcpi_div.quotient_msk\[30\] genblk2.pcpi_div.quotient_msk\[29\]
+ genblk2.pcpi_div.quotient_msk\[28\] VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__or4_1
XFILLER_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12124_ _06563_ _06565_ net869 VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13295__A net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12055_ _06505_ _06506_ net269 _06504_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__o211a_1
XFILLER_96_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12403__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10506__B1 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11006_ cpuregs\[8\]\[18\] net648 VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__or2_1
XFILLER_120_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10431__B _02702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12259__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12957_ net315 net2414 net453 VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__mux2_1
XFILLER_34_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11908_ _06377_ _06378_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__or2_1
XANTENNA__07686__B1 net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08328__S net531 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12888_ mem_rdata_q\[25\] net18 net964 VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__mux2_1
XFILLER_33_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627_ clknet_leaf_135_clk _01012_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11839_ _06309_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__inv_2
XFILLER_159_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09948__A net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14558_ clknet_leaf_199_clk _00944_ VGND VGND VPWR VPWR cpuregs\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11689__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13509_ net1690 net317 net419 VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__mux2_1
X_14489_ clknet_leaf_92_clk _00878_ VGND VGND VPWR VPWR instr_slli sky130_fd_sc_hd__dfxtp_1
XANTENNA__08650__A2 net1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09159__S net502 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07030_ net1115 _02599_ genblk2.pcpi_div.quotient\[16\] VGND VGND VPWR VPWR _02600_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07468__A net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08998__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08981_ net1626 _04267_ net946 VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__mux2_1
X_07932_ _03373_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__nand2_1
XANTENNA__12498__B1 net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10622__A net773 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07863_ _03268_ _03314_ _03373_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__and3_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06814_ net2572 net2550 net1649 VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__or3_1
X_09602_ _03770_ reg_next_pc\[7\] net921 VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__mux2_2
X_07794_ net256 net994 VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__nand2_1
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09622__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ count_instr\[43\] _04382_ count_instr\[44\] VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_104_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13144__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09464_ net3040 _04338_ net1229 VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_121_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08238__S net940 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ net324 net2450 net530 VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__mux2_1
X_09395_ net2361 net280 net401 VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__mux2_1
XANTENNA__12983__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout525_A _03774_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08346_ reg_pc\[6\] _03764_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__xor2_1
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08277_ net1020 _03722_ net980 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__mux2_2
XFILLER_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09069__S net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07228_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__inv_2
XFILLER_165_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12725__B2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07159_ genblk1.genblk1.pcpi_mul.pcpi_rd\[1\] genblk2.pcpi_div.pcpi_rd\[1\] net1112
+ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1222_X net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10170_ count_cycle\[61\] count_cycle\[62\] _04873_ count_cycle\[63\] VGND VGND VPWR
+ VPWR _04877_ sky130_fd_sc_hd__a31o_1
XANTENNA__10803__Y _05491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1106 net1107 VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__clkbuf_2
Xfanout1117 net1124 VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__buf_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1128 decoded_imm_j\[20\] VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13150__A1 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1139 net1140 VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__buf_2
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10251__B net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_X net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13860_ clknet_leaf_43_clk _00314_ VGND VGND VPWR VPWR cpuregs\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07841__A net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12811_ net349 net1996 net463 VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__mux2_1
XANTENNA__07117__C1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13791_ clknet_leaf_7_clk _00245_ VGND VGND VPWR VPWR cpuregs\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13054__S net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15530_ clknet_leaf_29_clk _01866_ VGND VGND VPWR VPWR cpuregs\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12742_ _02410_ net912 VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__nor2_1
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10672__C1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12893__S net965 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15461_ clknet_leaf_85_clk _00013_ VGND VGND VPWR VPWR mem_wordsize\[1\] sky130_fd_sc_hd__dfxtp_1
X_12673_ net1201 genblk1.genblk1.pcpi_mul.next_rs2\[38\] net892 net2894 net712 VGND
+ VGND VPWR VPWR _01343_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_190_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_190_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11624_ _06188_ _06212_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__or2_1
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14412_ clknet_leaf_178_clk alu_out\[12\] VGND VGND VPWR VPWR alu_out_q\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11216__A1 net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06891__A1 net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ clknet_leaf_52_clk _01731_ VGND VGND VPWR VPWR cpuregs\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11555_ is_beq_bne_blt_bge_bltu_bgeu net1233 net747 VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__and3_2
XFILLER_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14343_ clknet_leaf_75_clk _06731_ VGND VGND VPWR VPWR reg_out\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12194__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10707__A net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10506_ net986 decoded_imm\[1\] net856 VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a21o_1
X_14274_ clknet_leaf_97_clk _00728_ VGND VGND VPWR VPWR count_cycle\[19\] sky130_fd_sc_hd__dfxtp_1
X_11486_ _02368_ _06152_ net1208 VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13225_ net1045 net1042 net757 VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__mux2_1
XFILLER_109_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10437_ _05135_ _05136_ net818 VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__mux2_1
XANTENNA__10727__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13156_ net1506 net308 net432 VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__mux2_1
X_10368_ net833 _05069_ _05071_ _05073_ net793 VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__a2111o_1
X_12107_ net863 _06547_ _06548_ _06550_ _06551_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__a32o_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13087_ net318 net1698 net440 VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__mux2_1
X_10299_ _04997_ _05004_ _04999_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__a21o_1
X_12038_ net1019 _06484_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__or2_1
XANTENNA__11257__B net702 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09896__A1 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06919__X _02507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07751__A net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13444__A2 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13989_ clknet_leaf_22_clk _00443_ VGND VGND VPWR VPWR cpuregs\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15728_ net1179 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12652__B1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_181_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_181_clk sky130_fd_sc_hd__clkbuf_8
X_08200_ _03312_ _03682_ _03313_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_32_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09180_ _03810_ net1808 net497 VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__mux2_1
X_08131_ _03328_ _03332_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09397__B net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08062_ net967 _03375_ net932 _03374_ _03564_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__a221o_1
X_07013_ net1115 _02584_ net3043 VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12707__A1 net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12707__B2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12391__X _06664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12183__A2 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12551__B net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10623__Y _05316_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13139__S net431 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11448__A net817 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08964_ genblk1.genblk1.pcpi_mul.rd\[20\] genblk1.genblk1.pcpi_mul.rd\[52\] net955
+ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__mux2_1
XANTENNA__08139__A1 net966 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08139__B2 net929 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07915_ _03302_ _03432_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__nand2_1
XANTENNA__12978__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08895_ net1200 net2674 net893 _04224_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__a22o_1
XANTENNA__11143__B1 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12891__A0 mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07846_ _03361_ _03363_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__nand2_2
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09352__S net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07777_ net253 net1000 VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__nand2_1
XANTENNA__10498__S net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09639__B2 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09516_ net3060 _04372_ _04374_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__o21a_1
XANTENNA__12643__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11997__A2 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09447_ _04328_ _04329_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout430_X net430 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_172_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_172_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1172_X net1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout528_X net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13199__A1 net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09378_ net1843 net344 net399 VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__mux2_1
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07600__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12726__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08329_ reg_out\[3\] alu_out_q\[3\] net1154 VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__mux2_1
XFILLER_138_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10184__A_N net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11340_ cpuregs\[9\]\[27\] net638 net613 _06012_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__o211a_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout897_X net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11271_ _05933_ _05936_ _03171_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__o21a_1
XANTENNA__12742__A _02410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13010_ net526 net2299 net443 VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__mux2_1
XFILLER_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10222_ decoded_imm\[12\] net1026 VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08431__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13049__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10153_ count_cycle\[56\] _04864_ count_cycle\[57\] VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a21o_1
X_10084_ _04821_ _04822_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__nor2_1
X_14961_ clknet_leaf_145_clk _01313_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 cpuregs\[0\]\[31\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13912_ clknet_leaf_181_clk _00366_ VGND VGND VPWR VPWR cpuregs\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12882__A0 mem_rdata_q\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14892_ clknet_leaf_151_clk _01244_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13843_ clknet_leaf_24_clk _00297_ VGND VGND VPWR VPWR cpuregs\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11437__A1 net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10986_ cpuregs\[24\]\[17\] net648 VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13774_ clknet_leaf_37_clk _00228_ VGND VGND VPWR VPWR cpuregs\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11988__A2 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15513_ clknet_leaf_175_clk _01849_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dfxtp_1
X_12725_ net1190 net1732 net2133 net883 _02096_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_163_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_163_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13512__S net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15444_ clknet_leaf_10_clk _01783_ VGND VGND VPWR VPWR cpuregs\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12656_ net3014 net902 _02077_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_61_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ net2572 net561 _06193_ _06201_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__a22o_1
XANTENNA__11540__B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15375_ clknet_leaf_194_clk _01714_ VGND VGND VPWR VPWR cpuregs\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12587_ net346 net2401 net467 VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__mux2_1
XANTENNA__10948__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14326_ clknet_leaf_174_clk _06744_ VGND VGND VPWR VPWR reg_out\[6\] sky130_fd_sc_hd__dfxtp_1
X_11538_ mem_rdata_q\[31\] net2588 net736 VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__mux2_1
XFILLER_117_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold408 cpuregs\[16\]\[7\] VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11967__S net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold419 cpuregs\[10\]\[13\] VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ cpuregs\[26\]\[30\] net690 VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__or2_1
X_14257_ clknet_leaf_127_clk _00711_ VGND VGND VPWR VPWR count_cycle\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12165__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13208_ _02137_ _02138_ _02475_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__a21o_1
X_14188_ clknet_leaf_100_clk _00642_ VGND VGND VPWR VPWR count_instr\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13139_ net1670 net537 net431 VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__mux2_1
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1108 cpuregs\[1\]\[23\] VGND VGND VPWR VPWR net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 _01407_ VGND VGND VPWR VPWR net2433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12798__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07700_ _03218_ _03219_ net801 VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__mux2_1
XANTENNA__12873__A0 mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08680_ _04043_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__inv_2
XANTENNA__09172__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07631_ net986 decoded_imm_j\[3\] _03150_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__o21a_2
XANTENNA__10884__C1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06809__B net983 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07562_ reg_pc\[28\] decoded_imm\[28\] VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__or2_1
XANTENNA__12625__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09301_ net1503 net578 net480 VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__mux2_1
XANTENNA__10636__C1 net827 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_154_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_154_clk sky130_fd_sc_hd__clkbuf_8
X_07493_ _03007_ _03010_ _03021_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__a21o_1
XFILLER_22_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09232_ net1360 net581 net491 VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__mux2_1
XFILLER_167_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09163_ _03744_ _03745_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__or2_1
XANTENNA__14815__Q decoded_imm\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08114_ _03611_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__inv_2
X_09094_ net2250 net587 net506 VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__mux2_1
XFILLER_162_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08045_ _03287_ net934 VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__nor2_1
XANTENNA__10781__S net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold920 _01417_ VGND VGND VPWR VPWR net2234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 cpuregs\[19\]\[13\] VGND VGND VPWR VPWR net2245 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A instr_rdinstrh VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold942 reg_next_pc\[8\] VGND VGND VPWR VPWR net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09347__S net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold953 cpuregs\[1\]\[17\] VGND VGND VPWR VPWR net2267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold964 cpuregs\[7\]\[19\] VGND VGND VPWR VPWR net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 genblk1.genblk1.pcpi_mul.next_rs1\[40\] VGND VGND VPWR VPWR net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold986 genblk1.genblk1.pcpi_mul.pcpi_rd\[21\] VGND VGND VPWR VPWR net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11178__A net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold997 cpuregs\[6\]\[3\] VGND VGND VPWR VPWR net2311 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ net1185 _04452_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1018_X net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09871__A net1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout380_X net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08947_ net2739 _04250_ net943 VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout478_X net478 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A net858 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1620 _06587_ VGND VGND VPWR VPWR net2934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12864__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1631 genblk1.genblk1.pcpi_mul.next_rs2\[61\] VGND VGND VPWR VPWR net2945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1642 genblk1.genblk1.pcpi_mul.next_rs2\[62\] VGND VGND VPWR VPWR net2956 sky130_fd_sc_hd__dlygate4sd3_1
X_08878_ genblk1.genblk1.pcpi_mul.rd\[61\] genblk1.genblk1.pcpi_mul.next_rs2\[62\]
+ net1107 VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__nand3_1
Xhold1653 genblk1.genblk1.pcpi_mul.rd\[43\] VGND VGND VPWR VPWR net2967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1664 genblk1.genblk1.pcpi_mul.next_rs2\[46\] VGND VGND VPWR VPWR net2978 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09082__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1675 genblk2.pcpi_div.dividend\[31\] VGND VGND VPWR VPWR net2989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1686 _06580_ VGND VGND VPWR VPWR net3000 sky130_fd_sc_hd__dlygate4sd3_1
X_07829_ _03344_ _03346_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__and2_1
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1697 genblk2.pcpi_div.quotient\[4\] VGND VGND VPWR VPWR net3011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout645_X net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ _05500_ _05509_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__a21oi_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10771_ cpuregs\[28\]\[12\] cpuregs\[29\]\[12\] net650 VGND VGND VPWR VPWR _05459_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout812_X net812 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_145_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_145_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_158_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_142_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12510_ _02001_ _02002_ net385 VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__o21ba_1
X_13490_ net1775 net579 net422 VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__mux2_1
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08426__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12441_ net1178 _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_23_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15160_ clknet_leaf_89_clk _01509_ VGND VGND VPWR VPWR mem_rdata_q\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12372_ net1441 net345 net361 VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__mux2_1
XFILLER_165_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_157_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11323_ cpuregs\[18\]\[26\] net555 _05996_ net786 VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__o22a_1
X_14111_ clknet_leaf_2_clk _00565_ VGND VGND VPWR VPWR cpuregs\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15091_ clknet_leaf_182_clk _01443_ VGND VGND VPWR VPWR cpuregs\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12472__A net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12147__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09257__S net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14042_ clknet_leaf_196_clk _00496_ VGND VGND VPWR VPWR cpuregs\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11254_ cpuregs\[6\]\[25\] cpuregs\[7\]\[25\] net706 VGND VGND VPWR VPWR _05929_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10205_ decoded_imm\[21\] net1009 VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__nor2_1
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08220__B1 net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11185_ cpuregs\[25\]\[23\] net634 net610 _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__o211a_1
X_10136_ _04854_ _04855_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__nor2_1
XANTENNA__13507__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10067_ _04811_ net1236 _04810_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__and3b_1
XANTENNA__12411__S net474 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14944_ clknet_leaf_38_clk _01296_ VGND VGND VPWR VPWR cpuregs\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11658__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14875_ clknet_leaf_18_clk _01227_ VGND VGND VPWR VPWR cpuregs\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkload1_A clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13826_ clknet_leaf_12_clk _00280_ VGND VGND VPWR VPWR cpuregs\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12607__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08287__A0 net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13757_ clknet_leaf_1_clk _00211_ VGND VGND VPWR VPWR cpuregs\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_136_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_136_clk sky130_fd_sc_hd__clkbuf_8
X_10969_ cpuregs\[8\]\[17\] net655 VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__or2_1
XANTENNA__11551__A net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12708_ net1198 genblk1.genblk1.pcpi_mul.next_rs1\[3\] net914 net1043 VGND VGND VPWR
+ VPWR _02088_ sky130_fd_sc_hd__a22o_1
X_13688_ clknet_leaf_113_clk _00142_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_130_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13032__A0 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15427_ clknet_leaf_57_clk _01766_ VGND VGND VPWR VPWR cpuregs\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12639_ net1200 genblk1.genblk1.pcpi_mul.next_rs2\[19\] net919 net244 VGND VGND VPWR
+ VPWR _02069_ sky130_fd_sc_hd__a22o_1
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11043__C1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15358_ clknet_leaf_55_clk _01698_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_1
XANTENNA__11697__S net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14309_ clknet_leaf_101_clk _00763_ VGND VGND VPWR VPWR count_cycle\[54\] sky130_fd_sc_hd__dfxtp_1
Xhold205 cpuregs\[15\]\[13\] VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 cpuregs\[24\]\[8\] VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15289_ clknet_leaf_30_clk _01630_ VGND VGND VPWR VPWR cpuregs\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold227 cpuregs\[30\]\[21\] VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__B1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold238 cpuregs\[20\]\[12\] VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold249 cpuregs\[30\]\[11\] VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13335__B2 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14370__Q net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _04438_ _04439_ _04611_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__and3_1
Xfanout707 _03139_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__buf_2
Xfanout718 net720 VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_111_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 net730 VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__clkbuf_4
XFILLER_98_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ genblk1.genblk1.pcpi_mul.rd\[49\] genblk1.genblk1.pcpi_mul.next_rs2\[50\]
+ net1096 VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__nand3_1
X_06993_ net951 _02566_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__or3_1
X_09781_ _04525_ _04534_ _04535_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__and3_1
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08732_ _04087_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__inv_2
XANTENNA__11649__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08663_ _04028_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__inv_2
XFILLER_82_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07614_ net1080 decoded_imm_j\[17\] VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__or2_1
X_08594_ _03968_ _03970_ _03963_ _03966_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__a211o_1
XANTENNA__09630__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07545_ reg_pc\[27\] decoded_imm\[27\] VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_127_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_127_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout340_A _03807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_clk_X clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13152__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10085__B1 net1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07476_ reg_pc\[22\] decoded_imm\[22\] VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_153_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09215_ net1713 net330 net492 VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__mux2_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12991__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout605_A net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09146_ net1656 net340 net500 VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__mux2_1
XANTENNA__13388__A net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07253__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09077_ net1852 net336 net508 VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__mux2_1
XANTENNA__07253__B2 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13326__A1 net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08028_ net968 _03362_ net934 _03361_ _03534_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__o221a_1
XANTENNA__09077__S net508 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 cpuregs\[6\]\[5\] VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net975 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout595_X net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold761 cpuregs\[16\]\[5\] VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 cpuregs\[6\]\[25\] VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08202__B1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold783 cpuregs\[11\]\[11\] VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold794 _01414_ VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09979_ _04741_ _04744_ _04742_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__a21o_1
XANTENNA__11636__A mem_rdata_q\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ net1826 net314 net449 VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1450 net218 VGND VGND VPWR VPWR net2764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1461 genblk2.pcpi_div.divisor\[25\] VGND VGND VPWR VPWR net2775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1472 _01056_ VGND VGND VPWR VPWR net2786 sky130_fd_sc_hd__dlygate4sd3_1
X_11941_ net1049 net1052 net726 net866 VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__a31o_1
Xhold1483 count_cycle\[60\] VGND VGND VPWR VPWR net2797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1494 genblk2.pcpi_div.quotient\[22\] VGND VGND VPWR VPWR net2808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14660_ clknet_leaf_139_clk _01045_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient_msk\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11872_ _06302_ _06303_ _06337_ _06342_ _06301_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_28_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08269__A0 net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13611_ clknet_leaf_10_clk _00066_ VGND VGND VPWR VPWR cpuregs\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_10823_ cpuregs\[28\]\[13\] cpuregs\[29\]\[13\] net651 VGND VGND VPWR VPWR _05510_
+ sky130_fd_sc_hd__mux2_1
X_14591_ clknet_leaf_104_clk _00977_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_118_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13062__S net534 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13542_ net316 net1757 net417 VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__mux2_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10754_ cpuregs\[2\]\[11\] cpuregs\[3\]\[11\] net653 VGND VGND VPWR VPWR _05443_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10685_ cpuregs\[27\]\[9\] net627 net594 _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__o211a_1
X_13473_ net1576 net329 net423 VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__mux2_1
X_15212_ clknet_leaf_49_clk _01561_ VGND VGND VPWR VPWR cpuregs\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12424_ net910 net1217 net2990 VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__mux2_1
XFILLER_127_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09776__A decoded_imm_j\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15143_ clknet_leaf_73_clk _01495_ VGND VGND VPWR VPWR cpuregs\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12355_ net1218 genblk1.genblk1.pcpi_mul.mul_counter\[5\] net956 net917 VGND VGND
+ VPWR VPWR _06661_ sky130_fd_sc_hd__a22o_1
XANTENNA__12406__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11306_ cpuregs\[11\]\[26\] net643 net601 _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__o211a_1
X_15074_ clknet_leaf_103_clk _01426_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12286_ mem_rdata_q\[31\] net559 _06621_ net532 VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__a211o_1
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11237_ net808 _05910_ _05912_ net839 VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__a211o_1
X_14025_ clknet_leaf_49_clk _00479_ VGND VGND VPWR VPWR cpuregs\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__S net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output67_A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11168_ net831 _05841_ _05843_ _05845_ net792 VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__a2111o_1
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10119_ count_cycle\[44\] _04841_ count_cycle\[45\] VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a21o_1
X_11099_ cpuregs\[8\]\[20\] net657 VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__or2_1
XFILLER_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14927_ clknet_leaf_23_clk _01279_ VGND VGND VPWR VPWR cpuregs\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11980__S net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14858_ clknet_leaf_17_clk _01210_ VGND VGND VPWR VPWR cpuregs\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13809_ clknet_leaf_21_clk _00263_ VGND VGND VPWR VPWR cpuregs\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_109_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_8
X_14789_ clknet_leaf_109_clk _01142_ VGND VGND VPWR VPWR genblk2.pcpi_div.instr_rem
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07330_ count_instr\[44\] net1131 net1136 count_instr\[12\] VGND VGND VPWR VPWR _02871_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08066__S net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07261_ reg_pc\[8\] decoded_imm\[8\] VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__or2_1
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09000_ net526 net1957 net516 VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA__09686__A decoded_imm_j\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07192_ count_cycle\[3\] net971 net842 _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_113_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07235__A1 _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11031__A2 net855 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09902_ net1150 _04679_ _04680_ _04681_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__a22o_1
Xfanout504 _04279_ VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_8
XFILLER_116_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout515 _04276_ VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkbuf_4
Xfanout526 net527 VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkbuf_2
Xfanout537 net538 VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkbuf_2
X_09833_ _04567_ _04582_ _04593_ _04606_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__and4_1
Xfanout548 _03741_ VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout290_A _03860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout559 _06622_ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__buf_2
XFILLER_59_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13147__S net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net390 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09764_ net1183 _04432_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__or2_1
X_06976_ genblk2.pcpi_div.dividend\[8\] genblk2.pcpi_div.dividend\[7\] _02541_ VGND
+ VGND VPWR VPWR _02553_ sky130_fd_sc_hd__or3_1
X_08715_ _04072_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__inv_2
XANTENNA__12295__A1 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12986__S net447 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09695_ net1182 _04426_ net848 VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout555_A _03156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09160__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08646_ _04012_ _04014_ _04007_ _04010_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__a211o_1
XANTENNA__07171__B1 net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09360__S net478 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13390__B _04884_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout722_A net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08577_ net891 _03954_ _03956_ net2626 net1192 VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout1085_X net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09999__B1 net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07528_ net1069 net1003 _03055_ net1085 _03054_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__a221o_1
XFILLER_167_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout510_X net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07459_ net1073 _02984_ _02991_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout608_X net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07668__X _03189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10470_ net987 decoded_imm\[0\] net856 VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__a21o_1
XFILLER_136_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12734__B net911 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07226__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09129_ _03743_ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__or2_2
XFILLER_68_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07828__B net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12140_ net1223 _06258_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__and2_1
XFILLER_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12071_ _06276_ _06514_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__and2b_1
Xhold580 cpuregs\[24\]\[0\] VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 cpuregs\[8\]\[1\] VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _05702_ _05703_ net809 VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__mux2_1
XANTENNA__07844__A net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11730__B1 _06243_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13057__S net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12286__A1 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ net1871 net542 net448 VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__mux2_1
XANTENNA__12896__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1280 genblk1.genblk1.pcpi_mul.next_rs1\[38\] VGND VGND VPWR VPWR net2594 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ clknet_leaf_162_clk _01097_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1291 count_cycle\[0\] VGND VGND VPWR VPWR net2605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10836__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11924_ genblk2.pcpi_div.divisor\[43\] genblk2.pcpi_div.divisor\[42\] genblk2.pcpi_div.divisor\[41\]
+ genblk2.pcpi_div.divisor\[40\] VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__or4_1
XANTENNA__07162__B1 net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09270__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14643_ clknet_leaf_161_clk _01028_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11855_ _06314_ _06325_ _06312_ _06313_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__o211ai_2
XANTENNA_output105_A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10806_ net1164 net854 _05492_ _05493_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__a22o_1
XFILLER_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14574_ clknet_leaf_50_clk _00960_ VGND VGND VPWR VPWR cpuregs\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_11786_ genblk2.pcpi_div.outsign _05120_ _06256_ _06257_ VGND VGND VPWR VPWR _01008_
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13525_ net574 net1795 net418 VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__mux2_1
XFILLER_158_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10737_ _05424_ _05425_ net800 VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__mux2_1
XFILLER_158_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13456_ net1677 net583 net425 VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__mux2_1
XANTENNA__06923__A net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10668_ net839 _05356_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_11_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12407_ net342 net1954 net471 VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__mux2_1
XANTENNA__07217__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10599_ net801 _05289_ _05291_ net829 VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__o211a_1
X_13387_ _05013_ _05015_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_93_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput107 net107 VGND VGND VPWR VPWR mem_la_wdata[19] sky130_fd_sc_hd__buf_2
Xoutput118 net118 VGND VGND VPWR VPWR mem_la_wdata[29] sky130_fd_sc_hd__buf_2
XFILLER_154_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15126_ clknet_leaf_3_clk _01478_ VGND VGND VPWR VPWR cpuregs\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xoutput129 net129 VGND VGND VPWR VPWR mem_la_write sky130_fd_sc_hd__buf_2
XFILLER_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12338_ net1148 decoded_imm_j\[5\] net743 VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__and3_1
XFILLER_114_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15057_ clknet_leaf_105_clk net2481 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_12269_ net176 _04298_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__nor2_1
X_14008_ clknet_leaf_190_clk _00462_ VGND VGND VPWR VPWR cpuregs\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10524__A1 net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06830_ _02427_ _02430_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__or3_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07940__A2 _02384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06761_ mem_do_rinst VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__inv_2
XFILLER_83_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08500_ genblk1.genblk1.pcpi_mul.rd\[3\] genblk1.genblk1.pcpi_mul.next_rs2\[4\] net1098
+ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__nand3_1
X_09480_ _04350_ _04351_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__nor2_1
XANTENNA__10827__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09180__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08431_ net313 net2222 net530 VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__mux2_1
XFILLER_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08362_ _03779_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__nor2_1
XANTENNA__11237__C1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07313_ net1139 count_cycle\[43\] net976 _02854_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__a211o_1
XANTENNA__07456__A1 genblk2.pcpi_div.pcpi_rd\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08293_ net1006 _03730_ net982 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__mux2_2
XANTENNA__11252__A2 _05926_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07244_ _02761_ _02776_ _02777_ _02775_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a31oi_1
XFILLER_165_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07208__A1 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07175_ _02723_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__nand2_1
XFILLER_118_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1045_A net225 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1212_A net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout301 _03849_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09355__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout312 net315 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout323 _03826_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__buf_1
Xfanout334 _03815_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout672_A net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout345 _03802_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_2
Xfanout356 net357 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08479__B net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout367 net370 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_2
X_09816_ net1183 _04436_ _04602_ _02489_ net846 VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1000_X net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout378 net379 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_2
XFILLER_47_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout389 net390 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07931__A2 net995 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09747_ _04536_ _04537_ _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout460_X net460 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06959_ net1126 _02538_ genblk2.pcpi_div.dividend\[6\] VGND VGND VPWR VPWR _02539_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout558_X net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09678_ _04475_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__inv_2
XANTENNA__09090__S net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13217__A0 _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08629_ net903 _03998_ _04000_ net2660 net1210 VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__a32o_1
X_11640_ decoded_imm_j\[4\] net17 net546 VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__mux2_1
XFILLER_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10249__B net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11571_ _02382_ net547 _06187_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09841__C1 net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07398__X _02935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13310_ _02226_ _02227_ _02228_ net395 net1024 VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__o32a_1
XANTENNA__07839__A net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10522_ cpuregs\[12\]\[5\] cpuregs\[13\]\[5\] net675 VGND VGND VPWR VPWR _05217_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14290_ clknet_leaf_127_clk _00744_ VGND VGND VPWR VPWR count_cycle\[35\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08434__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13241_ net1042 net753 VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__or2_1
X_10453_ _05151_ _05152_ net816 VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__mux2_1
XANTENNA__10265__A decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10384_ genblk2.pcpi_div.quotient_msk\[27\] genblk2.pcpi_div.quotient_msk\[26\] genblk2.pcpi_div.quotient_msk\[25\]
+ genblk2.pcpi_div.quotient_msk\[24\] VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__or4_1
X_13172_ net1549 net537 net427 VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__mux2_1
XFILLER_109_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12123_ net995 _06564_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09265__S net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12054_ _06280_ _06283_ _06498_ net867 VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__a31o_1
XANTENNA__10506__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09372__A1 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11005_ net796 _05684_ _05686_ net823 VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__o211a_1
XANTENNA__07383__B1 _02909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input21_X net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout890 net891 VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__buf_2
XANTENNA_output222_A net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13_0_clk_X clknet_4_13_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13515__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10809__A2 net620 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12956_ net317 net2065 net452 VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__mux2_1
XANTENNA__06918__A net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11907_ genblk2.pcpi_div.divisor\[25\] genblk2.pcpi_div.dividend\[25\] VGND VGND
+ VPWR VPWR _06378_ sky130_fd_sc_hd__and2b_1
X_12887_ mem_rdata_q\[24\] net17 net964 VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__mux2_1
X_14626_ clknet_leaf_135_clk _01011_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ genblk2.pcpi_div.divisor\[5\] genblk2.pcpi_div.dividend\[5\] VGND VGND VPWR
+ VPWR _06309_ sky130_fd_sc_hd__and2b_1
XFILLER_159_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07438__A1 genblk2.pcpi_div.pcpi_rd\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14557_ clknet_leaf_195_clk _00943_ VGND VGND VPWR VPWR cpuregs\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11769_ _06245_ _06246_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_40_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_119_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07749__A net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13508_ net1794 net320 net419 VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__mux2_1
XANTENNA__08344__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14488_ clknet_leaf_95_clk _00877_ VGND VGND VPWR VPWR instr_sw sky130_fd_sc_hd__dfxtp_1
XFILLER_158_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13439_ _05031_ _05033_ net961 VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15109_ clknet_leaf_34_clk _01461_ VGND VGND VPWR VPWR cpuregs\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07610__A1 genblk2.pcpi_div.pcpi_rd\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08980_ genblk1.genblk1.pcpi_mul.rd\[28\] genblk1.genblk1.pcpi_mul.rd\[60\] net957
+ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__mux2_1
XFILLER_170_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09175__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07931_ _02398_ net995 _03447_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__o22a_1
XANTENNA__11718__B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07862_ _03291_ _03297_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09601_ reg_pc\[6\] net876 _04427_ net846 VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__a22o_1
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09903__S net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06813_ mem_do_wdata net1234 _02418_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__and3_1
XFILLER_113_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07793_ _03308_ _03310_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__nand2_1
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09532_ count_instr\[43\] _04382_ _04384_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__o21a_1
XANTENNA__07126__B1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14818__Q decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09463_ count_instr\[19\] _04338_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_121_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08414_ _03819_ _03822_ net767 VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__mux2_1
X_09394_ net2263 net282 net401 VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07429__A1 net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08345_ reg_out\[6\] alu_out_q\[6\] net1153 VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout420_A net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1162_A net241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13160__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net519 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10433__B1 net1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08276_ reg_out\[15\] reg_next_pc\[15\] net921 VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__mux2_1
XANTENNA__12284__B net739 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08107__X alu_out\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07227_ reg_pc\[6\] decoded_imm\[6\] VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__nand2_1
XFILLER_138_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1048_X net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07158_ reg_pc\[1\] decoded_imm\[1\] VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__nand2_1
XFILLER_133_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07601__A1 net1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_168_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07601__B2 net1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07089_ net1121 _02650_ genblk2.pcpi_div.quotient\[24\] VGND VGND VPWR VPWR _02651_
+ sky130_fd_sc_hd__a21o_1
XFILLER_161_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09085__S net511 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1107 net1108 VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1120 VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__buf_2
XFILLER_114_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1129 decoded_imm_j\[20\] VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_98_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13438__A0 net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10959__S net811 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_X net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12810_ net352 net1781 net463 VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__mux2_1
XFILLER_90_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11449__C1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13790_ clknet_leaf_11_clk _00244_ VGND VGND VPWR VPWR cpuregs\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12110__B1 net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12741_ net2511 net897 _02104_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__a21o_1
XANTENNA__07668__A1 net775 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15460_ clknet_leaf_85_clk _00012_ VGND VGND VPWR VPWR mem_wordsize\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12672_ net1200 net2894 net892 net2953 net712 VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_13_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ clknet_leaf_177_clk alu_out\[11\] VGND VGND VPWR VPWR alu_out_q\[11\] sky130_fd_sc_hd__dfxtp_1
X_11623_ mem_rdata_q\[3\] _02401_ _06208_ _06211_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__or4_1
X_15391_ clknet_leaf_50_clk _01730_ VGND VGND VPWR VPWR cpuregs\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__A2 net859 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13070__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14342_ clknet_leaf_76_clk _06730_ VGND VGND VPWR VPWR reg_out\[22\] sky130_fd_sc_hd__dfxtp_1
X_11554_ _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__inv_2
XFILLER_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14463__Q net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10505_ net987 _05203_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__nor2_1
X_14273_ clknet_leaf_97_clk _00727_ VGND VGND VPWR VPWR count_cycle\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11485_ net1061 _02487_ _05125_ _06152_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__or4_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13224_ net960 _04958_ _02152_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__nor3_1
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10436_ cpuregs\[4\]\[0\] cpuregs\[5\]\[0\] net697 VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__mux2_1
X_13155_ net1680 net312 net433 VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__mux2_1
X_10367_ cpuregs\[27\]\[31\] net638 net599 _05072_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__o211a_1
XFILLER_88_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12414__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12106_ net1001 net725 _06549_ net863 VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__a31oi_1
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13086_ net321 net2003 net440 VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__mux2_1
X_10298_ decoded_imm\[18\] net1014 VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_89_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_8
X_12037_ _06290_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__xor2_1
XANTENNA__10869__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07751__B net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08339__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13988_ clknet_leaf_43_clk _00442_ VGND VGND VPWR VPWR cpuregs\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15727_ net1181 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07659__A1 net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12939_ net571 net2036 net451 VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__mux2_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ clknet_leaf_104_clk _00995_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dfxtp_1
X_15589_ clknet_leaf_57_clk _01925_ VGND VGND VPWR VPWR cpuregs\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_13_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_08130_ _03330_ _03333_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__nand2_1
XFILLER_159_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__14373__Q net241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08061_ _03376_ net930 VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__nor2_1
XANTENNA__07198__B decoded_imm\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07012_ genblk2.pcpi_div.dividend\[13\] _02578_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__or2_1
XFILLER_161_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08963_ net1676 _04258_ net944 VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__mux2_1
XFILLER_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07914_ _03356_ _03365_ _03431_ _03417_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__o31ai_1
XFILLER_97_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08894_ _03892_ _03894_ _03891_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11143__A1 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07845_ net1165 net1028 VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__or2_1
XANTENNA__12891__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10779__S net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout468_A _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13155__S net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07776_ _03292_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__nor2_1
XFILLER_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09639__A2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09515_ count_instr\[37\] _04372_ net1206 VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12994__S net450 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12643__B2 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09869__A net1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09446_ net2974 _04326_ net1228 VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__o21ai_1
XFILLER_40_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13199__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06873__A2 net975 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09377_ net1762 net348 net399 VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout423_X net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_A net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1165_X net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08328_ net581 net2206 net531 VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__mux2_1
XFILLER_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08259_ net1038 _03713_ net980 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_134_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11270_ net794 _05940_ _05942_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__or4_1
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout792_X net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12742__B net912 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10221_ _04924_ _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__nand2_1
XANTENNA__07586__B1 _03109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10152_ net2758 _04864_ _04865_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__a21oi_1
XFILLER_161_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10083_ net2788 _04820_ net1235 VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__o21ai_1
X_14960_ clknet_leaf_144_clk _01312_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 cpuregs\[0\]\[7\] VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07852__A net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13911_ clknet_leaf_181_clk _00365_ VGND VGND VPWR VPWR cpuregs\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_input29_A mem_rdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12882__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14891_ clknet_leaf_105_clk _01243_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10689__S net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10342__C1 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10893__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_28_clk _00296_ VGND VGND VPWR VPWR cpuregs\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13773_ clknet_leaf_57_clk _00227_ VGND VGND VPWR VPWR cpuregs\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ _05666_ _05667_ net796 VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__mux2_1
XFILLER_71_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15512_ clknet_leaf_175_clk _01848_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dfxtp_1
X_12724_ _02405_ net911 VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__nor2_1
X_15443_ clknet_leaf_1_clk _01782_ VGND VGND VPWR VPWR cpuregs\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12655_ net1212 genblk1.genblk1.pcpi_mul.next_rs2\[27\] net917 net253 VGND VGND VPWR
+ VPWR _02077_ sky130_fd_sc_hd__a22o_1
XANTENNA__12409__S net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11606_ net2654 net562 _06189_ _06201_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__a22o_1
XFILLER_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15374_ clknet_leaf_193_clk _01713_ VGND VGND VPWR VPWR cpuregs\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12586_ net349 net2159 net467 VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14193__Q reg_pc\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07274__C1 _02817_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14325_ clknet_leaf_134_clk _06743_ VGND VGND VPWR VPWR reg_out\[5\] sky130_fd_sc_hd__dfxtp_1
X_11537_ mem_rdata_q\[30\] net194 net736 VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__mux2_1
Xhold409 net45 VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output97_A net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14256_ clknet_leaf_127_clk net2907 VGND VGND VPWR VPWR count_cycle\[1\] sky130_fd_sc_hd__dfxtp_1
X_11468_ cpuregs\[25\]\[30\] net637 net612 _06137_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__o211a_1
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13207_ net1045 net759 VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__or2_1
X_10419_ mem_do_prefetch _02490_ _05121_ _05122_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__o211a_1
X_14187_ clknet_leaf_100_clk _00641_ VGND VGND VPWR VPWR count_instr\[58\] sky130_fd_sc_hd__dfxtp_1
X_11399_ net1083 _06069_ net857 VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13138_ net1524 net541 net432 VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__mux2_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07893__A_N net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13069_ net575 net2008 net440 VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__mux2_1
Xhold1109 net185 VGND VGND VPWR VPWR net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07329__B1 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12322__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07762__A net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12873__A1 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11676__A2 net747 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10900__B net649 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07630_ net986 decoded_imm_j\[3\] _03150_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__o21ai_1
XFILLER_54_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14368__Q net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07561_ _03037_ _03048_ _03083_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__o31a_1
XANTENNA__12667__X _02083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12625__B2 net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09300_ net1380 net581 net482 VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07492_ _03007_ _03010_ _03021_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__nand3_1
X_09231_ net1490 net583 net490 VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__mux2_1
XFILLER_22_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09162_ net2061 net280 net503 VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__mux2_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13050__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08113_ _03593_ _03608_ _03610_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__o21a_1
XFILLER_148_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09093_ _04275_ _04277_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__nor2_4
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09628__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08044_ net770 _03548_ _03549_ _03542_ VGND VGND VPWR VPWR alu_out\[12\] sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_116_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold910 cpuregs\[2\]\[5\] VGND VGND VPWR VPWR net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 cpuregs\[9\]\[17\] VGND VGND VPWR VPWR net2235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 cpuregs\[13\]\[28\] VGND VGND VPWR VPWR net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 cpuregs\[6\]\[23\] VGND VGND VPWR VPWR net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 cpuregs\[5\]\[4\] VGND VGND VPWR VPWR net2268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11364__A1 _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold965 cpuregs\[18\]\[6\] VGND VGND VPWR VPWR net2279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold976 _01410_ VGND VGND VPWR VPWR net2290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_1_0_clk_X clknet_4_1_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold987 cpuregs\[17\]\[11\] VGND VGND VPWR VPWR net2301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 cpuregs\[1\]\[11\] VGND VGND VPWR VPWR net2312 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ net1152 _04765_ _04764_ _02380_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__a211o_1
XANTENNA__12989__S net448 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_A _03751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08946_ genblk1.genblk1.pcpi_mul.rd\[11\] genblk1.genblk1.pcpi_mul.rd\[43\] net954
+ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1610 genblk1.genblk1.pcpi_mul.rd\[39\] VGND VGND VPWR VPWR net2924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1621 count_instr\[25\] VGND VGND VPWR VPWR net2935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1632 _01367_ VGND VGND VPWR VPWR net2946 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08877_ genblk1.genblk1.pcpi_mul.next_rs2\[62\] net1106 genblk1.genblk1.pcpi_mul.rd\[61\]
+ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__a21o_1
XFILLER_57_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1643 _01368_ VGND VGND VPWR VPWR net2957 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout373_X net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1654 count_cycle\[59\] VGND VGND VPWR VPWR net2968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1665 genblk1.genblk1.pcpi_mul.next_rs2\[35\] VGND VGND VPWR VPWR net2979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1676 genblk1.genblk1.pcpi_mul.mul_counter\[0\] VGND VGND VPWR VPWR net2990 sky130_fd_sc_hd__dlygate4sd3_1
X_07828_ net1160 net1016 VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__nand2_1
Xhold1687 count_cycle\[52\] VGND VGND VPWR VPWR net3001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1698 genblk1.genblk1.pcpi_mul.mul_counter\[1\] VGND VGND VPWR VPWR net3012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07740__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout540_X net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07759_ net1177 net1045 VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__or2_1
XFILLER_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10770_ net1165 net853 _05457_ _05458_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__a22o_1
XANTENNA__09493__B1 net1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09429_ _04316_ _04317_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout805_X net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12440_ net1180 net717 VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13041__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12371_ net1446 net348 net360 VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__mux2_1
XFILLER_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14110_ clknet_leaf_11_clk _00564_ VGND VGND VPWR VPWR cpuregs\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13201__X _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11322_ cpuregs\[19\]\[26\] net642 net602 VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__o21a_1
XFILLER_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08442__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15090_ clknet_leaf_179_clk _01442_ VGND VGND VPWR VPWR cpuregs\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14041_ clknet_leaf_191_clk _00495_ VGND VGND VPWR VPWR cpuregs\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11253_ _02396_ _05133_ _05928_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10204_ _04908_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__nand2_1
XANTENNA__06901__D net1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08220__A1 net1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08220__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12899__S net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11184_ cpuregs\[24\]\[23\] net685 VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__or2_1
X_10135_ net2783 _04853_ net1229 VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11107__A1 net247 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09273__S net485 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10066_ count_cycle\[23\] count_cycle\[24\] count_cycle\[25\] _04804_ VGND VGND VPWR
+ VPWR _04811_ sky130_fd_sc_hd__and4_1
X_14943_ clknet_leaf_15_clk _01295_ VGND VGND VPWR VPWR cpuregs\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10866__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14874_ clknet_leaf_39_clk _01226_ VGND VGND VPWR VPWR cpuregs\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_13825_ clknet_leaf_42_clk _00279_ VGND VGND VPWR VPWR cpuregs\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_91_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12607__B2 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13523__S net418 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10618__B1 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13756_ clknet_leaf_4_clk _00210_ VGND VGND VPWR VPWR cpuregs\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_10968_ net798 _05648_ _05650_ net824 VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__o211a_1
XANTENNA__11551__B net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12707_ net1191 net1491 net2544 net897 _02087_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__a221o_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11291__B1 _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13687_ clknet_leaf_113_clk _00141_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_10899_ _05582_ _05583_ net796 VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__mux2_1
X_15426_ clknet_leaf_53_clk _01765_ VGND VGND VPWR VPWR cpuregs\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12638_ net2633 net890 _02068_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__a21o_1
XFILLER_129_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15357_ clknet_leaf_55_clk _01697_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12569_ net258 _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14308_ clknet_leaf_98_clk _00762_ VGND VGND VPWR VPWR count_cycle\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15288_ clknet_leaf_40_clk _01629_ VGND VGND VPWR VPWR cpuregs\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold206 net150 VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 cpuregs\[8\]\[18\] VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold228 genblk1.genblk1.pcpi_mul.next_rs1\[9\] VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 cpuregs\[24\]\[28\] VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ clknet_leaf_175_clk _00693_ VGND VGND VPWR VPWR reg_next_pc\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12543__B1 _02396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout708 net709 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_111_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__C1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 net720 VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__buf_2
X_08800_ genblk1.genblk1.pcpi_mul.rd\[49\] genblk1.genblk1.pcpi_mul.next_rs2\[50\]
+ net1096 VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_74_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09780_ _04568_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__inv_2
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12602__S net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06992_ net1118 _02565_ genblk2.pcpi_div.quotient\[11\] VGND VGND VPWR VPWR _02567_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_112_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09183__S net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08731_ _04079_ _04082_ _04084_ _04085_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__o211a_1
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08662_ genblk1.genblk1.pcpi_mul.rd\[28\] genblk1.genblk1.pcpi_mul.rdx\[28\] VGND
+ VGND VPWR VPWR _04028_ sky130_fd_sc_hd__nand2_1
XFILLER_66_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07613_ net991 _03127_ _03134_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08593_ genblk1.genblk1.pcpi_mul.rd\[17\] genblk1.genblk1.pcpi_mul.next_rs2\[18\]
+ net1100 VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__nand3_1
X_07544_ _03064_ _03068_ _03070_ _02703_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__o22a_1
XANTENNA__12557__B net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07475_ reg_pc\[22\] decoded_imm\[22\] VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__or2_1
XFILLER_139_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout333_A _03815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1075_A cpu_state\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09214_ net1714 net333 net492 VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09145_ net1758 net343 net500 VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout500_A net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09358__S net477 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09076_ net1599 net339 net508 VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__mux2_1
XANTENNA__08262__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07253__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13326__A2 _05599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08027_ _03364_ net930 VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__or2_1
XFILLER_162_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold740 cpuregs\[2\]\[30\] VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1030_X net1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold751 cpuregs\[3\]\[21\] VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 cpuregs\[8\]\[30\] VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1128_X net1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold773 cpuregs\[23\]\[5\] VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 cpuregs\[31\]\[27\] VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold795 net179 VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09978_ _04749_ _04750_ net2586 net879 VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11636__B mem_rdata_q\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08929_ net1436 _04241_ net944 VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__mux2_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout755_X net755 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1440 _06609_ VGND VGND VPWR VPWR net2754 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1451 genblk1.genblk1.pcpi_mul.rd\[13\] VGND VGND VPWR VPWR net2765 sky130_fd_sc_hd__dlygate4sd3_1
X_11940_ net1052 net726 net1049 VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_146_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1462 genblk2.pcpi_div.quotient_msk\[16\] VGND VGND VPWR VPWR net2776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 count_cycle\[17\] VGND VGND VPWR VPWR net2787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08010__B net934 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1484 genblk2.pcpi_div.quotient_msk\[10\] VGND VGND VPWR VPWR net2798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1495 _06601_ VGND VGND VPWR VPWR net2809 sky130_fd_sc_hd__dlygate4sd3_1
X_11871_ _06304_ _06341_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout922_X net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ clknet_leaf_199_clk _00065_ VGND VGND VPWR VPWR cpuregs\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_10822_ net788 _05504_ _05506_ _05508_ net776 VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__o41a_1
XFILLER_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14590_ clknet_leaf_114_clk _00976_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_9_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13541_ net320 net2044 net415 VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__mux2_1
X_10753_ _05440_ _05441_ net813 VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13472_ net1595 net334 net423 VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__mux2_1
X_10684_ cpuregs\[26\]\[9\] net670 VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__or2_1
X_15211_ clknet_leaf_50_clk _01560_ VGND VGND VPWR VPWR cpuregs\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11025__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12423_ net279 net2010 net473 VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__mux2_1
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15142_ clknet_leaf_46_clk _01494_ VGND VGND VPWR VPWR cpuregs\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09268__S net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12354_ genblk1.genblk1.pcpi_mul.mul_counter\[4\] _06658_ _02415_ VGND VGND VPWR
+ VPWR _06660_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08172__S net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ cpuregs\[10\]\[26\] net694 VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__or2_1
XFILLER_114_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15073_ clknet_leaf_103_clk net2237 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12285_ _02428_ net745 VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__and2_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11328__A1 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14024_ clknet_leaf_71_clk _00478_ VGND VGND VPWR VPWR cpuregs\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07864__X _03382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11236_ cpuregs\[5\]\[24\] net642 net819 _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_56_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output252_A net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13518__S net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12422__S net473 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11167_ cpuregs\[27\]\[22\] net633 net597 _05844_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__o211a_1
X_10118_ count_cycle\[44\] _04841_ _04843_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__o21a_1
X_11098_ net798 _05775_ _05777_ net824 VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__o211a_1
XFILLER_64_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10049_ _04798_ _04799_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__nor2_1
XFILLER_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14926_ clknet_leaf_17_clk _01278_ VGND VGND VPWR VPWR cpuregs\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14857_ clknet_leaf_32_clk _01209_ VGND VGND VPWR VPWR cpuregs\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07180__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13808_ clknet_leaf_29_clk _00262_ VGND VGND VPWR VPWR cpuregs\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14788_ clknet_leaf_109_clk _01141_ VGND VGND VPWR VPWR genblk2.pcpi_div.instr_divu
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12056__A2 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13253__A1 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08347__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13739_ clknet_leaf_105_clk _00193_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07260_ _02795_ _02796_ _02805_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__a21o_1
XFILLER_32_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11016__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15409_ clknet_leaf_4_clk _01748_ VGND VGND VPWR VPWR cpuregs\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_07191_ count_instr\[3\] net1135 net976 _02740_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09178__S net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07235__A2 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14381__Q net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13308__A2 net564 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09901_ _04443_ _04673_ net1150 VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout505 _04279_ VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__buf_2
Xfanout516 net517 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__buf_4
Xfanout527 _03774_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__buf_1
X_09832_ _04593_ _04596_ _04606_ _04616_ _04605_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__a32o_1
XFILLER_101_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout538 net540 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__buf_1
XFILLER_99_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10641__A net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_141_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout549 net551 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__buf_4
XANTENNA__10542__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09763_ net1149 _04550_ _04553_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__a21o_1
X_06975_ _02551_ _02552_ net951 _02549_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout283_A _03870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08714_ genblk1.genblk1.pcpi_mul.rd\[36\] genblk1.genblk1.pcpi_mul.rdx\[36\] VGND
+ VGND VPWR VPWR _04072_ sky130_fd_sc_hd__nand2_1
X_09694_ _04486_ _04487_ _04490_ net1182 VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__o211a_1
XANTENNA__07950__A net1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08645_ genblk1.genblk1.pcpi_mul.rd\[25\] genblk1.genblk1.pcpi_mul.next_rs2\[26\]
+ net1105 VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_156_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout548_A _03741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13163__S net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1192_A net1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11472__A net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__inv_2
XANTENNA__13244__A1 net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08257__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13244__B2 net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07527_ genblk1.genblk1.pcpi_mul.pcpi_rd\[25\] genblk2.pcpi_div.pcpi_rd\[25\] net1113
+ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_22_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A net716 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1078_X net1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07458_ net358 _02985_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__o21bai_1
XFILLER_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11007__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13399__A _02412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_X net503 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10816__A net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07389_ _02880_ _02892_ _02907_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand3_1
XFILLER_136_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09088__S net510 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09128_ latched_rd\[1\] latched_rd\[0\] VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__nand2_1
XFILLER_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10766__C1 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09059_ latched_rd\[3\] latched_rd\[4\] latched_rd\[2\] VGND VGND VPWR VPWR _04277_
+ sky130_fd_sc_hd__nand3b_4
XFILLER_151_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12070_ genblk2.pcpi_div.dividend\[21\] _06519_ net270 VGND VGND VPWR VPWR _01030_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold570 cpuregs\[6\]\[2\] VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 cpuregs\[10\]\[8\] VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold592 cpuregs\[27\]\[21\] VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ cpuregs\[20\]\[18\] cpuregs\[21\]\[18\] net647 VGND VGND VPWR VPWR _05703_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07844__B net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ net1821 net573 net448 VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__mux2_1
XFILLER_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1270 count_instr\[49\] VGND VGND VPWR VPWR net2584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input11_A mem_rdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07860__A net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1281 genblk2.pcpi_div.quotient\[26\] VGND VGND VPWR VPWR net2595 sky130_fd_sc_hd__dlygate4sd3_1
X_14711_ clknet_leaf_153_clk _01096_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_11923_ genblk2.pcpi_div.divisor\[39\] genblk2.pcpi_div.divisor\[38\] genblk2.pcpi_div.divisor\[37\]
+ genblk2.pcpi_div.divisor\[36\] VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__or4_1
Xhold1292 pcpi_timeout_counter\[2\] VGND VGND VPWR VPWR net2606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12691__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13073__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14642_ clknet_leaf_165_clk _01027_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13235__A1 net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11854_ _06316_ _06323_ _06324_ _06315_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__o211a_1
X_10805_ net1075 _05491_ net854 VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11246__B1 net611 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14573_ clknet_leaf_54_clk _00959_ VGND VGND VPWR VPWR cpuregs\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11785_ net1189 genblk2.pcpi_div.instr_rem net866 net1216 VGND VGND VPWR VPWR _06257_
+ sky130_fd_sc_hd__a211o_1
X_13524_ net576 net1661 net415 VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__mux2_1
XANTENNA__09787__A _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10736_ cpuregs\[30\]\[11\] cpuregs\[31\]\[11\] net665 VGND VGND VPWR VPWR _05425_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13455_ net1581 net587 net426 VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__mux2_1
X_10667_ cpuregs\[1\]\[9\] net550 _05357_ net800 net828 VGND VGND VPWR VPWR _05358_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__12417__S net474 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12406_ _03802_ net2000 net471 VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ net1007 net393 _02293_ _02295_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__a22o_1
X_10598_ net815 _05290_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15125_ clknet_leaf_192_clk _01477_ VGND VGND VPWR VPWR cpuregs\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xoutput108 net1179 VGND VGND VPWR VPWR mem_la_wdata[1] sky130_fd_sc_hd__buf_2
X_12337_ decoded_imm\[6\] net735 _06643_ mem_rdata_q\[26\] _06648_ VGND VGND VPWR
+ VPWR _01168_ sky130_fd_sc_hd__a221o_1
XFILLER_142_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 net1177 VGND VGND VPWR VPWR mem_la_wdata[2] sky130_fd_sc_hd__buf_2
XFILLER_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15056_ clknet_leaf_102_clk _01408_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12268_ net1192 _05096_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__nor2_1
X_14007_ clknet_leaf_183_clk _00461_ VGND VGND VPWR VPWR cpuregs\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09914__A1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11219_ _05893_ _05894_ net819 VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__mux2_1
XFILLER_68_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12199_ genblk2.pcpi_div.quotient_msk\[13\] net271 net2834 VGND VGND VPWR VPWR _06592_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_96_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11721__A1 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput90 net90 VGND VGND VPWR VPWR mem_la_addr[4] sky130_fd_sc_hd__buf_2
XFILLER_68_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10180__B net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06760_ latched_store VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__inv_2
X_14909_ clknet_leaf_121_clk _01261_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12682__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07153__A1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ _03832_ _03835_ net768 VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__mux2_1
XANTENNA__06900__A1 net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14376__Q net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08361_ reg_pc\[9\] reg_pc\[8\] _03772_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__and3_1
XFILLER_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07312_ count_instr\[43\] net1131 net1135 count_instr\[11\] VGND VGND VPWR VPWR _02854_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09697__A decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08292_ reg_out\[23\] reg_next_pc\[23\] net926 VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__mux2_1
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07243_ net1071 _02779_ _02780_ _02789_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__a31o_1
XANTENNA__06833__B net1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07174_ reg_pc\[2\] decoded_imm\[2\] VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__or2_1
XFILLER_117_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12201__A2 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08106__A _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1038_A net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11960__A1 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09636__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13158__S net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout302 _03849_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_1
XANTENNA_fanout498_A net499 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout313 net315 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10371__A net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout324 net325 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout335 _03815_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1205_A _02378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout346 _03802_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input3_A mem_rdata[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout357 _03791_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_2
X_09815_ _04600_ _04601_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__nor2_1
XANTENNA__12997__S net449 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout368 net369 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_2
Xfanout379 net384 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_2
XANTENNA_fanout665_A net672 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09746_ _04536_ _04537_ _02480_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13465__A1 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06958_ genblk2.pcpi_div.dividend\[5\] genblk2.pcpi_div.dividend\[4\] _02528_ VGND
+ VGND VPWR VPWR _02538_ sky130_fd_sc_hd__or3_1
XFILLER_86_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09371__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11473__Y _06143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09677_ decoded_imm_j\[4\] _04425_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__and2_1
XANTENNA__12673__C1 net712 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06889_ net991 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout832_A net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_X net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08628_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__inv_2
XFILLER_82_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout620_X net620 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08559_ _03940_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout718_X net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11570_ _02369_ net6 _02452_ _06186_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__or4_1
XFILLER_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10521_ cpuregs\[14\]\[5\] cpuregs\[15\]\[5\] net675 VGND VGND VPWR VPWR _05216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10546__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12728__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13240_ net1047 net754 _02166_ net709 VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__o211a_1
XFILLER_155_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10452_ cpuregs\[20\]\[0\] cpuregs\[21\]\[0\] net687 VGND VGND VPWR VPWR _05152_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10265__B net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13171_ net1753 net541 net428 VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__mux2_1
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10383_ _05084_ _05085_ _05087_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__or3_1
XFILLER_163_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12122_ net997 _06558_ net725 VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_36_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08303__X net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08450__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13068__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12053_ _06280_ _06498_ _06283_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_53_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11004_ net809 _05685_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__or2_1
XANTENNA__07383__A1 net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout880 net881 VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07383__B2 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout891 net898 VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12259__A2 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09281__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input14_X net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12955_ net323 net2028 net452 VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__mux2_1
XFILLER_34_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output215_A net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11906_ genblk2.pcpi_div.dividend\[25\] genblk2.pcpi_div.divisor\[25\] VGND VGND
+ VPWR VPWR _06377_ sky130_fd_sc_hd__and2b_1
XFILLER_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12886_ mem_rdata_q\[23\] net16 net964 VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__mux2_1
XANTENNA__07686__A2 net623 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11837_ genblk2.pcpi_div.divisor\[6\] genblk2.pcpi_div.dividend\[6\] VGND VGND VPWR
+ VPWR _06308_ sky130_fd_sc_hd__xor2_1
X_14625_ clknet_leaf_129_clk _01010_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13531__S net416 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14556_ clknet_leaf_195_clk _00942_ VGND VGND VPWR VPWR cpuregs\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11768_ net167 net130 net536 VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux2_1
XFILLER_158_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10442__A1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10719_ cpuregs\[25\]\[10\] net627 net608 _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__o211a_1
X_13507_ net1952 net324 net421 VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__mux2_1
X_14487_ clknet_leaf_94_clk _00876_ VGND VGND VPWR VPWR instr_andi sky130_fd_sc_hd__dfxtp_1
XFILLER_158_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07749__B net996 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11699_ net1769 net340 net373 VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__mux2_1
X_13438_ net996 _02341_ net398 VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__mux2_1
XFILLER_127_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13369_ _02275_ _02276_ _02280_ net397 net1010 VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__o32a_1
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11942__B2 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15108_ clknet_leaf_33_clk _01460_ VGND VGND VPWR VPWR cpuregs\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_170_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08213__X alu_out\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07930_ _02399_ net996 net994 _02398_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__a22o_1
XFILLER_130_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15039_ clknet_leaf_129_clk net2106 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11718__C net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12498__A2 net716 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09980__A net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07861_ _03377_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__or2_2
XFILLER_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07374__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09600_ _03767_ reg_next_pc\[6\] net921 VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_108_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06812_ net1234 _02417_ _02418_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__and3_1
XFILLER_96_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07792_ _03309_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ count_instr\[43\] _04382_ net1214 VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a21oi_1
XFILLER_25_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09462_ _04338_ _04339_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__nor2_1
XFILLER_92_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08413_ _03820_ _03821_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__nor2_1
X_09393_ net2145 net288 net402 VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08344_ net542 net2537 net528 VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__mux2_1
XFILLER_149_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08275_ net1022 _03721_ net980 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__mux2_1
XANTENNA_fanout413_A _02358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1155_A net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07226_ net1071 _02763_ _02764_ _02773_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__a31o_1
XFILLER_165_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07157_ reg_pc\[1\] decoded_imm\[1\] VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__or2_1
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09366__S net402 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08270__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07601__A2 net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07088_ genblk2.pcpi_div.quotient\[23\] _02644_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout782_A _03152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1108 net1109 VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1208_X net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1119 net1120 VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input6_X net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_X net570 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09729_ _04502_ _04505_ _04511_ _04512_ _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout835_X net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ net1190 net2089 net914 net1011 VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__a22o_1
XANTENNA__10672__A1 net813 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12671_ net1202 net2953 net894 net2979 net712 VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__a221o_1
XFILLER_169_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12756__A _02412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ clknet_leaf_171_clk alu_out\[10\] VGND VGND VPWR VPWR alu_out_q\[10\] sky130_fd_sc_hd__dfxtp_1
X_11622_ mem_rdata_q\[19\] mem_rdata_q\[18\] _06209_ _06210_ VGND VGND VPWR VPWR _06211_
+ sky130_fd_sc_hd__or4_1
XFILLER_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15390_ clknet_leaf_57_clk _01729_ VGND VGND VPWR VPWR cpuregs\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_168_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10547__Y _05242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14341_ clknet_leaf_76_clk _06729_ VGND VGND VPWR VPWR reg_out\[21\] sky130_fd_sc_hd__dfxtp_1
X_11553_ net746 _06175_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__and2_1
XFILLER_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10504_ net774 _05194_ _05202_ _05186_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__a31oi_4
X_14272_ clknet_leaf_97_clk _00726_ VGND VGND VPWR VPWR count_cycle\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11484_ cpu_state\[2\] _02471_ _06148_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__a211o_1
XFILLER_109_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13223_ _04948_ _04957_ _04956_ _04949_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__o211a_1
X_10435_ cpuregs\[6\]\[0\] cpuregs\[7\]\[0\] net684 VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__mux2_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09276__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13154_ net1759 net318 net432 VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__mux2_1
X_10366_ cpuregs\[26\]\[31\] net693 VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__or2_1
XFILLER_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12105_ net724 _06549_ net1001 VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__a21o_1
XFILLER_152_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13085_ net325 net2025 net441 VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__mux2_1
X_10297_ _04993_ _05002_ _04995_ _04915_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__and4b_1
X_12036_ _02360_ genblk2.pcpi_div.dividend\[16\] _06358_ VGND VGND VPWR VPWR _06490_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13526__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09750__C1 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13429__A1 net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06929__A _02509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08305__A0 net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13987_ clknet_leaf_13_clk _00441_ VGND VGND VPWR VPWR cpuregs\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12938_ net576 net2114 net451 VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12869_ net29 net2947 _02450_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__mux2_1
XFILLER_34_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ clknet_leaf_104_clk _00994_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dfxtp_1
XFILLER_21_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08355__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15588_ clknet_leaf_54_clk _01924_ VGND VGND VPWR VPWR cpuregs\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14539_ clknet_leaf_91_clk _00927_ VGND VGND VPWR VPWR is_sll_srl_sra sky130_fd_sc_hd__dfxtp_1
X_08060_ net770 _03562_ _03563_ _03557_ VGND VGND VPWR VPWR alu_out\[14\] sky130_fd_sc_hd__a31o_1
XFILLER_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07011_ net950 _02583_ _02581_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__o21ai_1
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09186__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07595__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08962_ genblk1.genblk1.pcpi_mul.rd\[19\] genblk1.genblk1.pcpi_mul.rd\[51\] net955
+ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__mux2_1
XANTENNA__11679__A0 is_sb_sh_sw VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07913_ _03384_ _03427_ _03429_ _03318_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__o221a_1
XFILLER_102_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08893_ net1217 net2941 net904 _04223_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__a22o_1
XANTENNA__11143__A2 _05820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07844_ net1165 net1028 VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__nor2_1
XANTENNA__06839__A net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07775_ net251 net1004 VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__nor2_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09514_ _04372_ _04373_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__nor2_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09445_ count_instr\[13\] count_instr\[12\] _04325_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout530_A _03746_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout628_A net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13171__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09376_ net1684 net351 net399 VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__mux2_1
XANTENNA__08265__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08327_ _03752_ _02371_ net767 VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__mux2_2
XFILLER_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_X net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09272__A1 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_X net416 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1158_X net1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08258_ reg_out\[6\] reg_next_pc\[6\] net921 VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__mux2_1
XFILLER_20_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07209_ count_instr\[36\] net1130 net1135 count_instr\[4\] VGND VGND VPWR VPWR _02758_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08189_ _03266_ net935 net771 _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09096__S net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10220_ decoded_imm\[13\] net1024 VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__or2_1
XFILLER_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout785_X net785 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07586__A1 net1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10151_ count_cycle\[56\] _04864_ net1238 VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_18_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10082_ count_cycle\[29\] count_cycle\[30\] count_cycle\[31\] _04816_ VGND VGND VPWR
+ VPWR _04821_ sky130_fd_sc_hd__and4_2
XFILLER_0_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout952_X net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12331__A1 decoded_imm\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12331__B2 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13910_ clknet_leaf_180_clk _00364_ VGND VGND VPWR VPWR cpuregs\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07852__B net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14890_ clknet_leaf_105_clk _01242_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.mul_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13841_ clknet_leaf_21_clk _00295_ VGND VGND VPWR VPWR cpuregs\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_114_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13772_ clknet_leaf_52_clk _00226_ VGND VGND VPWR VPWR cpuregs\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10984_ cpuregs\[30\]\[17\] cpuregs\[31\]\[17\] net647 VGND VGND VPWR VPWR _05667_
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15511_ clknet_leaf_175_clk _01847_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_27_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12723_ net1190 net1335 net1732 net883 _02095_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__a221o_1
XANTENNA__07510__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13081__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15442_ clknet_leaf_195_clk _01781_ VGND VGND VPWR VPWR cpuregs\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12654_ net2724 net902 _02076_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__a21o_1
X_11605_ net2800 net561 _06180_ _06201_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__a22o_1
XFILLER_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15373_ clknet_leaf_181_clk _01712_ VGND VGND VPWR VPWR cpuregs\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12585_ net352 net2030 net467 VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11536_ mem_rdata_q\[29\] net2643 net736 VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__mux2_1
X_14324_ clknet_leaf_130_clk _06742_ VGND VGND VPWR VPWR reg_out\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11070__A1 net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14255_ clknet_leaf_127_clk _00709_ VGND VGND VPWR VPWR count_cycle\[0\] sky130_fd_sc_hd__dfxtp_1
X_11467_ cpuregs\[24\]\[30\] net690 VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__or2_1
X_13206_ _02384_ net759 VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nand2_1
X_10418_ net2852 _02490_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__nand2_1
X_14186_ clknet_leaf_100_clk _00640_ VGND VGND VPWR VPWR count_instr\[57\] sky130_fd_sc_hd__dfxtp_1
X_11398_ net1081 decoded_imm\[28\] VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__or2_1
XFILLER_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13137_ net1601 net571 net433 VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__mux2_1
X_10349_ cpuregs\[10\]\[31\] net694 VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__or2_1
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13068_ net579 net1953 net441 VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__mux2_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12019_ net1023 _06474_ _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12322__B2 mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10884__A1 net799 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07560_ _03058_ _03071_ _03083_ _03084_ _03072_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10636__A1 net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07491_ _03019_ _03020_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07501__A1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09230_ net1555 net587 net490 VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__mux2_1
XFILLER_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06825__C net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14384__Q net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09161_ net1934 net284 net502 VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09254__A1 _03844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08112_ net1159 net1013 _03609_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__a21oi_1
X_09092_ net1995 net278 net510 VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08043_ _03302_ _03547_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_116_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold900 cpuregs\[17\]\[16\] VGND VGND VPWR VPWR net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 cpuregs\[31\]\[1\] VGND VGND VPWR VPWR net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 genblk1.genblk1.pcpi_mul.next_rs1\[55\] VGND VGND VPWR VPWR net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold933 cpuregs\[18\]\[25\] VGND VGND VPWR VPWR net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 net57 VGND VGND VPWR VPWR net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold955 cpuregs\[9\]\[12\] VGND VGND VPWR VPWR net2269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11364__A2 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold966 cpuregs\[9\]\[1\] VGND VGND VPWR VPWR net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 cpuregs\[21\]\[19\] VGND VGND VPWR VPWR net2291 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _04761_ _04762_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1020_A net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold988 cpuregs\[11\]\[24\] VGND VGND VPWR VPWR net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 cpuregs\[9\]\[29\] VGND VGND VPWR VPWR net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09644__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08945_ net2435 _04249_ net943 VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout480_A net483 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1600 genblk1.genblk1.pcpi_mul.next_rs2\[5\] VGND VGND VPWR VPWR net2914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12313__A1 decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A _03756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13166__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1611 genblk2.pcpi_div.quotient\[5\] VGND VGND VPWR VPWR net2925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 mem_rdata_q\[4\] VGND VGND VPWR VPWR net2936 sky130_fd_sc_hd__dlygate4sd3_1
X_08876_ _04209_ _04208_ net2815 net1217 VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_4_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1633 mem_rdata_q\[6\] VGND VGND VPWR VPWR net2947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1644 genblk1.genblk1.pcpi_mul.next_rs2\[59\] VGND VGND VPWR VPWR net2958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1655 genblk1.genblk1.pcpi_mul.next_rs2\[58\] VGND VGND VPWR VPWR net2969 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10875__A1 net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07827_ net1160 net1016 VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__and2_1
Xhold1666 net198 VGND VGND VPWR VPWR net2980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1677 count_cycle\[62\] VGND VGND VPWR VPWR net2991 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_A _06163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_X net366 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1688 genblk1.genblk1.pcpi_mul.next_rs2\[23\] VGND VGND VPWR VPWR net3002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1699 count_instr\[55\] VGND VGND VPWR VPWR net3013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07758_ net1177 net1045 VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__and2_1
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout533_X net533 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07689_ net788 _03204_ _03206_ _03208_ net776 VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__o41a_1
XANTENNA_fanout912_A net913 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09428_ net2973 _04314_ net1225 VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__o21ai_1
XFILLER_158_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09359_ net1417 net292 net477 VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12370_ net1340 net351 net360 VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__mux2_1
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11321_ cpuregs\[17\]\[26\] net642 net615 _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__o211a_1
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14040_ clknet_leaf_186_clk _00494_ VGND VGND VPWR VPWR cpuregs\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12001__B1 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11252_ net1081 _05926_ _05927_ net858 VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__a211o_1
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10203_ decoded_imm\[22\] net1007 VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__or2_1
X_11183_ _05858_ _05859_ net819 VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__mux2_1
XANTENNA__08220__A2 net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10563__B1 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10134_ count_cycle\[47\] count_cycle\[50\] _04846_ _04852_ VGND VGND VPWR VPWR _04854_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11107__A2 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13076__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09705__C1 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10065_ count_cycle\[25\] _04808_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__or2_1
X_14942_ clknet_leaf_38_clk _01294_ VGND VGND VPWR VPWR cpuregs\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14873_ clknet_leaf_6_clk _01225_ VGND VGND VPWR VPWR cpuregs\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13824_ clknet_leaf_1_clk _00278_ VGND VGND VPWR VPWR cpuregs\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12068__B1 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13755_ clknet_leaf_4_clk _00209_ VGND VGND VPWR VPWR cpuregs\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10967_ net810 _05649_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12706_ _02402_ net911 VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__nor2_1
XFILLER_93_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10898_ cpuregs\[30\]\[15\] cpuregs\[31\]\[15\] net649 VGND VGND VPWR VPWR _05583_
+ sky130_fd_sc_hd__mux2_1
X_13686_ clknet_leaf_114_clk _00140_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_15425_ clknet_leaf_71_clk _01764_ VGND VGND VPWR VPWR cpuregs\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12637_ net1196 genblk1.genblk1.pcpi_mul.next_rs2\[18\] net915 net1160 VGND VGND
+ VPWR VPWR _02068_ sky130_fd_sc_hd__a22o_1
XFILLER_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11043__A1 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15356_ clknet_leaf_93_clk _01696_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfxtp_1
X_12568_ _05118_ net719 VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__nand2_1
XANTENNA__12240__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11519_ mem_rdata_q\[12\] net174 net740 VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__mux2_1
X_14307_ clknet_leaf_98_clk _00761_ VGND VGND VPWR VPWR count_cycle\[52\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_44_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15287_ clknet_leaf_14_clk _01628_ VGND VGND VPWR VPWR cpuregs\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12499_ genblk2.pcpi_div.divisor\[46\] net870 VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__nor2_1
Xhold207 cpuregs\[14\]\[15\] VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 cpuregs\[30\]\[3\] VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _01379_ VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14238_ clknet_leaf_176_clk _00692_ VGND VGND VPWR VPWR reg_next_pc\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14169_ clknet_leaf_125_clk _00623_ VGND VGND VPWR VPWR count_instr\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout709 _02501_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_111_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ net1118 genblk2.pcpi_div.quotient\[11\] _02565_ VGND VGND VPWR VPWR _02566_
+ sky130_fd_sc_hd__and3_1
XFILLER_140_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08730_ _04084_ _04085_ _04079_ _04082_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__a211o_1
XANTENNA__14379__Q net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08661_ net1212 net2921 net901 _04027_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_53_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07612_ net359 _03128_ _03133_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12059__B1 net1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08592_ genblk1.genblk1.pcpi_mul.rd\[17\] genblk1.genblk1.pcpi_mul.next_rs2\[18\]
+ net1096 VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_157_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07543_ net1142 count_cycle\[58\] count_cycle\[26\] net978 _03069_ VGND VGND VPWR
+ VPWR _03070_ sky130_fd_sc_hd__a221o_1
XFILLER_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11234__S net699 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07474_ _02998_ _03000_ _03005_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__or3_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09213_ net1734 net338 net493 VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11019__D1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1068_A net1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09144_ net1422 net347 net500 VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07300__X _02843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09075_ net1850 net343 net509 VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__mux2_1
XFILLER_162_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1235_A net1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11990__C1 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08026_ _03532_ _03533_ _03527_ VGND VGND VPWR VPWR alu_out\[10\] sky130_fd_sc_hd__o21ai_1
XANTENNA__07159__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold730 cpuregs\[16\]\[20\] VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 net200 VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout695_A net696 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold752 cpuregs\[27\]\[23\] VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 cpuregs\[23\]\[31\] VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold774 cpuregs\[16\]\[27\] VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold785 cpuregs\[7\]\[2\] VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold796 cpuregs\[19\]\[8\] VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09374__S net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07683__A net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09977_ net1185 _04450_ net849 VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout862_A net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11409__S net704 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08928_ genblk1.genblk1.pcpi_mul.rd\[2\] genblk1.genblk1.pcpi_mul.rd\[34\] net955
+ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__mux2_1
XANTENNA__11636__C mem_rdata_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1430 _01132_ VGND VGND VPWR VPWR net2744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 genblk1.genblk1.pcpi_mul.rd\[54\] VGND VGND VPWR VPWR net2755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 genblk2.pcpi_div.quotient\[23\] VGND VGND VPWR VPWR net2766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout650_X net650 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ genblk1.genblk1.pcpi_mul.rd\[58\] genblk1.genblk1.pcpi_mul.next_rs2\[59\]
+ net1108 VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__nand3_1
Xhold1463 _01057_ VGND VGND VPWR VPWR net2777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1474 count_cycle\[31\] VGND VGND VPWR VPWR net2788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1485 count_instr\[36\] VGND VGND VPWR VPWR net2799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1496 genblk2.pcpi_div.quotient_msk\[21\] VGND VGND VPWR VPWR net2810 sky130_fd_sc_hd__dlygate4sd3_1
X_11870_ _06300_ _06302_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__nor2_1
XFILLER_73_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09403__A net267 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10821_ cpuregs\[11\]\[13\] net619 net590 _05507_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_28_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout915_X net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10752_ cpuregs\[4\]\[11\] cpuregs\[5\]\[11\] net666 VGND VGND VPWR VPWR _05441_
+ sky130_fd_sc_hd__mux2_1
X_13540_ net324 net1904 net417 VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13471_ net1694 net336 net423 VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__mux2_1
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10683_ cpuregs\[25\]\[9\] net627 net608 _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__o211a_1
XANTENNA__09218__A1 net319 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12422_ net284 net1999 net473 VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__mux2_1
X_15210_ clknet_leaf_72_clk _01559_ VGND VGND VPWR VPWR cpuregs\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__06762__A net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14752__Q genblk2.pcpi_div.pcpi_ready VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12353_ genblk1.genblk1.pcpi_mul.mul_counter\[4\] _02415_ _06658_ VGND VGND VPWR
+ VPWR _06659_ sky130_fd_sc_hd__or3_1
X_15141_ clknet_leaf_49_clk _01493_ VGND VGND VPWR VPWR cpuregs\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10784__B1 net589 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ cpuregs\[9\]\[26\] net643 net615 _05977_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__o211a_1
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15072_ clknet_leaf_103_clk _01424_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12284_ decoded_imm\[31\] net739 VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__and2_1
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14023_ clknet_leaf_71_clk _00477_ VGND VGND VPWR VPWR cpuregs\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11235_ cpuregs\[4\]\[24\] net699 VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__or2_1
XANTENNA__10536__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09284__S net486 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11166_ cpuregs\[26\]\[22\] net683 VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__or2_1
XANTENNA_output245_A net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11319__S net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10117_ count_cycle\[44\] _04841_ net1206 VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11097_ net810 _05776_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__or2_1
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10048_ net2885 _04797_ net1229 VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__o21ai_1
X_14925_ clknet_leaf_31_clk _01277_ VGND VGND VPWR VPWR cpuregs\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold90 cpuregs\[20\]\[2\] VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13534__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07704__B2 net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14856_ clknet_leaf_48_clk _01208_ VGND VGND VPWR VPWR cpuregs\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07180__A2 net1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13807_ clknet_leaf_45_clk _00261_ VGND VGND VPWR VPWR cpuregs\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14787_ clknet_leaf_91_clk _01140_ VGND VGND VPWR VPWR mem_state\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13253__A2 net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11999_ net1032 net1030 _06448_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_119_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13738_ clknet_leaf_108_clk _00192_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13669_ clknet_leaf_145_clk _00123_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15408_ clknet_leaf_3_clk _01747_ VGND VGND VPWR VPWR cpuregs\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07768__A net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08363__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07190_ count_instr\[35\] net1130 net1139 count_cycle\[35\] VGND VGND VPWR VPWR _02740_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08216__X net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15339_ clknet_leaf_166_clk _01679_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12516__B2 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09900_ _04443_ _04672_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__or2_1
Xfanout506 _04279_ VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09194__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout517 net519 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__buf_4
X_09831_ _04590_ _04604_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__nand2_1
Xfanout528 _03746_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkload13_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout539 net540 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__clkbuf_2
XFILLER_101_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07943__A1 net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06974_ net1120 genblk2.pcpi_div.quotient\[8\] _02550_ net951 VGND VGND VPWR VPWR
+ _02552_ sky130_fd_sc_hd__a31o_1
X_09762_ net984 _04551_ _04552_ _02380_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__a31o_1
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07008__A net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08713_ net1200 net2931 net894 _04071_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__a22o_1
XFILLER_55_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09693_ net1149 _04488_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__or3b_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout276_A net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07950__B net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08644_ genblk1.genblk1.pcpi_mul.rd\[25\] genblk1.genblk1.pcpi_mul.next_rs2\[26\]
+ net1105 VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__and3_1
XFILLER_55_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12568__B net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _03947_ _03950_ _03952_ _03953_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__o211a_1
XANTENNA__13741__Q genblk1.genblk1.pcpi_mul.mul_waiting VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10369__A net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout443_A net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13244__A2 _05242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07526_ count_cycle\[25\] net973 net843 _03053_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__o211a_1
XANTENNA__12452__B1 net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07457_ net1067 net1010 _02989_ net1086 _02988_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout610_A net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07136__A_N net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09369__S net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08273__S net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07388_ reg_pc\[14\] decoded_imm\[14\] _02905_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__nand3_1
XANTENNA__13399__B net756 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09127_ latched_rd\[2\] latched_rd\[4\] latched_rd\[3\] VGND VGND VPWR VPWR _04281_
+ sky130_fd_sc_hd__nand3_2
XFILLER_108_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09058_ net278 net2419 net515 VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__mux2_1
X_08009_ net770 _03517_ _03518_ _03514_ VGND VGND VPWR VPWR alu_out\[8\] sky130_fd_sc_hd__a31o_1
XFILLER_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold560 cpuregs\[30\]\[2\] VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08187__A1 net1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold571 cpuregs\[15\]\[16\] VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 net184 VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ cpuregs\[22\]\[18\] cpuregs\[23\]\[18\] net647 VGND VGND VPWR VPWR _05702_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold593 cpuregs\[7\]\[3\] VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout865_X net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11730__A2 _06242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ net1532 net578 net448 VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1260 genblk1.genblk1.pcpi_mul.rd\[12\] VGND VGND VPWR VPWR net2574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _00632_ VGND VGND VPWR VPWR net2585 sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ clknet_leaf_162_clk _01095_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1282 _06605_ VGND VGND VPWR VPWR net2596 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ genblk2.pcpi_div.dividend\[31\] genblk2.pcpi_div.divisor\[31\] VGND VGND
+ VPWR VPWR _06393_ sky130_fd_sc_hd__and2b_1
XANTENNA__07860__B net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1293 reg_next_pc\[30\] VGND VGND VPWR VPWR net2607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08448__S net1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12691__B1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14641_ clknet_leaf_165_clk _01026_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11853_ genblk2.pcpi_div.dividend\[3\] genblk2.pcpi_div.divisor\[3\] VGND VGND VPWR
+ VPWR _06324_ sky130_fd_sc_hd__nand2b_1
XFILLER_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10804_ net1075 decoded_imm\[12\] VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__or2_1
X_14572_ clknet_leaf_69_clk _00958_ VGND VGND VPWR VPWR cpuregs\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_11784_ net1157 net258 _05118_ _03368_ genblk2.pcpi_div.instr_div VGND VGND VPWR
+ VPWR _06256_ sky130_fd_sc_hd__o311a_1
XANTENNA__08111__A1 net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13523_ net579 net1558 net418 VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__mux2_1
X_10735_ cpuregs\[28\]\[11\] cpuregs\[29\]\[11\] net665 VGND VGND VPWR VPWR _05424_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09279__S net484 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13454_ _03745_ _02127_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__nor2_1
X_10666_ cpuregs\[2\]\[9\] cpuregs\[3\]\[9\] net667 VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__mux2_1
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12405_ _03799_ net1727 net471 VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13385_ _04879_ _02294_ net393 VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__a21oi_1
X_10597_ cpuregs\[14\]\[7\] cpuregs\[15\]\[7\] net673 VGND VGND VPWR VPWR _05290_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15124_ clknet_leaf_187_clk _01476_ VGND VGND VPWR VPWR cpuregs\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR mem_la_wdata[20] sky130_fd_sc_hd__buf_2
X_12336_ net1148 decoded_imm_j\[6\] net744 VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__and3_1
XFILLER_108_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13529__S net416 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15055_ clknet_leaf_102_clk net2433 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_12267_ genblk2.pcpi_div.divisor\[30\] net380 net368 net2173 VGND VGND VPWR VPWR
+ _01136_ sky130_fd_sc_hd__a22o_1
XFILLER_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14006_ clknet_leaf_190_clk _00460_ VGND VGND VPWR VPWR cpuregs\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output72_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11218_ cpuregs\[28\]\[24\] cpuregs\[29\]\[24\] net697 VGND VGND VPWR VPWR _05894_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__S net1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11557__B mem_rdata_q\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12198_ net748 net2962 VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__nor2_1
Xoutput80 net80 VGND VGND VPWR VPWR mem_la_addr[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput91 net91 VGND VGND VPWR VPWR mem_la_addr[5] sky130_fd_sc_hd__buf_2
X_11149_ cpuregs\[1\]\[22\] net551 _05826_ net804 net831 VGND VGND VPWR VPWR _05827_
+ sky130_fd_sc_hd__a221o_1
XFILLER_110_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10888__S net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07138__C1 net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12131__C1 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07689__B1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14908_ clknet_leaf_142_clk _01260_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08358__S net529 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07153__A2 decoded_imm\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14839_ clknet_leaf_11_clk _01191_ VGND VGND VPWR VPWR cpuregs\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08360_ reg_pc\[8\] _03772_ reg_pc\[9\] VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11237__A1 net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12434__B1 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07311_ _02811_ _02852_ net1060 VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__o21a_1
X_08291_ net1007 _03729_ net982 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__mux2_2
XANTENNA__11512__S net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07242_ net1062 _02783_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__a21o_1
XANTENNA__09189__S net498 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07173_ reg_pc\[2\] decoded_imm\[2\] VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__nor2_1
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10748__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13162__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout303 net304 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout314 net315 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10371__B _05076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout325 net327 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11173__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A _04888_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07916__A1 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout336 net337 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_2
Xfanout347 net348 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_2
X_09814_ _04436_ _04586_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__and2b_1
XFILLER_59_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout358 _02914_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_2
Xfanout369 net370 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1100_A net1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09745_ _04524_ _04526_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__nand2_1
XFILLER_86_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06957_ genblk2.pcpi_div.quotient\[6\] _02535_ net953 VGND VGND VPWR VPWR _02537_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__13174__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11476__A1 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06888_ net1072 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__nand2_1
XANTENNA__08268__S net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09676_ decoded_imm_j\[4\] _04425_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__or2_1
XFILLER_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08627_ _03991_ _03994_ _03996_ _03997_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__o211a_1
XFILLER_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout446_X net446 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net826 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_X net1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12510__B1_N net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08558_ genblk1.genblk1.pcpi_mul.rd\[12\] genblk1.genblk1.pcpi_mul.rdx\[12\] VGND
+ VGND VPWR VPWR _03940_ sky130_fd_sc_hd__nand2_1
XANTENNA__12976__A1 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07509_ _03033_ _03036_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__nand2_1
XFILLER_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08489_ genblk1.genblk1.pcpi_mul.rd\[1\] genblk1.genblk1.pcpi_mul.next_rs2\[2\] net1101
+ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__and3_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10987__B1 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09099__S net507 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10520_ _05212_ _05214_ net785 VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__a21o_1
XFILLER_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12728__B2 net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10451_ cpuregs\[22\]\[0\] cpuregs\[23\]\[0\] net687 VGND VGND VPWR VPWR _05151_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10739__B1 net607 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11400__A1 net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13170_ net1640 net571 net429 VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__mux2_1
XFILLER_136_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10382_ genblk2.pcpi_div.quotient_msk\[3\] genblk2.pcpi_div.quotient_msk\[2\] genblk2.pcpi_div.quotient_msk\[1\]
+ genblk2.pcpi_div.quotient_msk\[0\] VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__or4_1
XFILLER_163_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout982_X net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12121_ _06384_ _06385_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_36_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12052_ net861 _06502_ _06503_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_53_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold390 cpuregs\[20\]\[21\] VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07907__A1 _02392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11003_ cpuregs\[14\]\[18\] cpuregs\[15\]\[18\] net655 VGND VGND VPWR VPWR _05685_
+ sky130_fd_sc_hd__mux2_1
Xfanout870 net871 VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__buf_2
XANTENNA__07383__A2 _02917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07871__A _03382_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout881 net882 VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net893 VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__buf_2
XFILLER_19_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13084__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12954_ net326 net2427 net452 VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__mux2_1
Xhold1090 cpuregs\[7\]\[31\] VGND VGND VPWR VPWR net2404 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ _06372_ _06375_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__or2_1
X_12885_ mem_rdata_q\[22\] net15 net962 VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_193_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_193_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_output208_A net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14624_ clknet_leaf_122_clk _01009_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11836_ genblk2.pcpi_div.divisor\[7\] genblk2.pcpi_div.dividend\[7\] VGND VGND VPWR
+ VPWR _06307_ sky130_fd_sc_hd__and2b_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14555_ clknet_leaf_3_clk _00941_ VGND VGND VPWR VPWR cpuregs\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08096__B1 _03465_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11767_ net268 net96 VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_101_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11332__S net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13506_ net1980 net329 net419 VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_140_clk_A clknet_4_7_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10718_ cpuregs\[24\]\[10\] net668 VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__or2_1
X_14486_ clknet_leaf_95_clk _00875_ VGND VGND VPWR VPWR instr_ori sky130_fd_sc_hd__dfxtp_1
XFILLER_158_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11698_ net1663 net345 net374 VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__mux2_1
XANTENNA__13427__A2_N _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12719__B2 net883 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13437_ _04879_ _02335_ _02337_ _02338_ _02340_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__o41a_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_3_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10649_ cpuregs\[27\]\[8\] net626 net594 _05340_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__o211a_1
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13368_ reg_pc\[20\] net566 _02278_ _02279_ net393 VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_155_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15107_ clknet_leaf_73_clk _01459_ VGND VGND VPWR VPWR cpuregs\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12319_ decoded_imm\[14\] net743 _06632_ _06638_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__o22a_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13299_ net708 _02196_ _02218_ net564 reg_pc\[12\] VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__a32o_1
XANTENNA__13144__A1 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15038_ clknet_leaf_135_clk _01390_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10191__B net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07860_ net240 net1022 VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__nor2_1
XFILLER_95_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07781__A net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06811_ mem_state\[0\] mem_state\[1\] VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__or2_1
X_07791_ net1172 net1041 VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__nor2_1
XFILLER_113_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11507__S net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09530_ _04382_ _04383_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__nor2_1
XANTENNA__12655__B1 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14387__Q net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09461_ net2774 _04337_ net1229 VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_184_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_184_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_121_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08412_ reg_pc\[19\] reg_pc\[18\] _03813_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__and3_1
X_09392_ net1989 net292 net401 VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__mux2_1
XFILLER_52_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08343_ _03762_ _03765_ net767 VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__mux2_1
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08274_ reg_out\[14\] reg_next_pc\[14\] net920 VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__mux2_1
XANTENNA__11091__C1 net838 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07225_ net1062 _02767_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__a21o_1
XANTENNA__13368__D1 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_A net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13383__A1 net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07156_ net12 net130 _02695_ net9 _02707_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__a221o_1
XANTENNA__06860__A net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08404__X _03815_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11394__B1 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13169__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07087_ genblk2.pcpi_div.dividend\[24\] net1121 _02647_ net948 VGND VGND VPWR VPWR
+ _02649_ sky130_fd_sc_hd__a31o_1
XFILLER_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout396_X net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1109 genblk1.genblk1.pcpi_mul.rs1\[0\] VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__buf_2
XANTENNA_fanout775_A _03170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12894__A0 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12801__S net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09382__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_A _02690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07989_ _03303_ _03308_ _03494_ _03309_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a31o_1
XANTENNA__11417__S net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11449__A1 net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09728_ _04503_ _04511_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__or2_1
XFILLER_170_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout730_X net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_175_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_175_clk sky130_fd_sc_hd__clkbuf_8
X_09659_ decoded_imm_j\[1\] _04422_ _04457_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__nand3_1
XFILLER_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout828_X net828 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12670_ net1202 net2979 net894 net3007 net713 VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__a221o_1
XFILLER_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12756__B net913 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11621_ mem_rdata_q\[0\] mem_rdata_q\[1\] VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14340_ clknet_leaf_76_clk _06728_ VGND VGND VPWR VPWR reg_out\[20\] sky130_fd_sc_hd__dfxtp_1
X_11552_ mem_rdata_q\[14\] mem_rdata_q\[13\] mem_rdata_q\[12\] VGND VGND VPWR VPWR
+ _06175_ sky130_fd_sc_hd__nor3_2
XFILLER_168_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10503_ net832 _05197_ _05199_ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__a211o_1
XFILLER_155_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11483_ _05125_ _06149_ _02387_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__and3b_1
X_14271_ clknet_leaf_84_clk _00725_ VGND VGND VPWR VPWR count_cycle\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12177__A2 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10434_ net1083 net1088 net1231 VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__o21ai_2
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13222_ _03227_ net568 VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__nor2_1
XANTENNA__08461__S net530 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06770__A net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11385__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13079__S net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10365_ cpuregs\[25\]\[31\] net638 net613 _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__o211a_1
X_13153_ net1647 net320 net432 VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__mux2_1
XFILLER_88_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12104_ net1003 _06542_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__or2_1
X_13084_ net329 net1561 net439 VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__mux2_1
XFILLER_151_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10296_ _04999_ _05001_ _04997_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__o21a_1
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11137__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12035_ genblk2.pcpi_div.dividend\[16\] _06489_ net269 VGND VGND VPWR VPWR _01025_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12885__A0 mem_rdata_q\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09292__S net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10360__A1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13429__A2 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12012__A net1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12637__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13986_ clknet_leaf_12_clk _00440_ VGND VGND VPWR VPWR cpuregs\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12937_ net580 net2184 net453 VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_166_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_166_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_103_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13542__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ net28 net3015 _02450_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11570__B net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14607_ clknet_leaf_114_clk _00993_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dfxtp_1
X_11819_ _06287_ _06288_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__nor2_1
X_15587_ clknet_leaf_59_clk _01923_ VGND VGND VPWR VPWR cpuregs\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12799_ net585 net2074 net465 VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14538_ clknet_leaf_88_clk _00926_ VGND VGND VPWR VPWR is_sb_sh_sw sky130_fd_sc_hd__dfxtp_2
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10186__B net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14469_ clknet_leaf_95_clk _00858_ VGND VGND VPWR VPWR instr_bne sky130_fd_sc_hd__dfxtp_1
X_07010_ genblk2.pcpi_div.quotient\[13\] _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12168__A2 net380 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08224__X net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11376__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09991__A net1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07595__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08961_ net2483 _04257_ net944 VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__mux2_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11128__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07912_ net1169 net1036 VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12876__A0 mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08892_ _04220_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07843_ net1165 net1028 VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__nand2_1
XFILLER_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06839__B net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07774_ net251 net1004 VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__and2_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09513_ net2799 _04370_ net1226 VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_157_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_157_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_37_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout356_A net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09444_ _04326_ _04327_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__nor2_1
XFILLER_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09375_ net1899 net355 net400 VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__mux2_1
XFILLER_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08326_ reg_out\[2\] alu_out_q\[2\] net1154 VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08257_ net1040 _03712_ net980 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__mux2_2
XFILLER_165_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_X net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11700__S net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12159__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09377__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07208_ net1062 _02754_ _02756_ net842 VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__a211o_1
X_08188_ _03268_ _03677_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08281__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07139_ _02383_ net17 _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__o21a_1
XANTENNA__08232__B1 net1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07586__A2 net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10150_ _04864_ net1238 _04863_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout778_X net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12867__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10081_ _04820_ net1235 _04819_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_7_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07625__S net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12331__A2 net735 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09406__A net1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08310__A net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10342__A1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_X net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11147__S net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_28_clk _00294_ VGND VGND VPWR VPWR cpuregs\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12619__B1 net915 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08299__A0 net1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13771_ clknet_leaf_70_clk _00225_ VGND VGND VPWR VPWR cpuregs\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_148_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_148_clk sky130_fd_sc_hd__clkbuf_8
X_10983_ cpuregs\[28\]\[17\] cpuregs\[29\]\[17\] net646 VGND VGND VPWR VPWR _05666_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11671__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15510_ clknet_leaf_173_clk _01846_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12722_ _02404_ net911 VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__nor2_1
XANTENNA__08456__S net768 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08309__X net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15441_ clknet_leaf_195_clk _01780_ VGND VGND VPWR VPWR cpuregs\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12653_ net1212 genblk1.genblk1.pcpi_mul.next_rs2\[26\] net918 net252 VGND VGND VPWR
+ VPWR _02076_ sky130_fd_sc_hd__a22o_1
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11604_ net1145 net563 _06175_ _06202_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__a22o_1
X_15372_ clknet_leaf_182_clk _01711_ VGND VGND VPWR VPWR cpuregs\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12584_ net357 net2181 net467 VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__mux2_1
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10802__C1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07274__A1 net1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14323_ clknet_leaf_133_clk _06741_ VGND VGND VPWR VPWR reg_out\[3\] sky130_fd_sc_hd__dfxtp_1
X_11535_ mem_rdata_q\[28\] net2729 net736 VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__mux2_1
XFILLER_129_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07274__B2 net1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11070__A2 net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06771__Y _02379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09287__S net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14254_ clknet_leaf_87_clk _00708_ VGND VGND VPWR VPWR reg_next_pc\[31\] sky130_fd_sc_hd__dfxtp_1
X_11466_ _06134_ _06135_ net805 VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__mux2_1
XANTENNA__08044__X alu_out\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13205_ net569 _05203_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__nor2_1
X_10417_ net1208 _02451_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__nor2_1
XFILLER_136_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08223__B1 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14185_ clknet_leaf_100_clk _00639_ VGND VGND VPWR VPWR count_instr\[56\] sky130_fd_sc_hd__dfxtp_1
X_11397_ net774 _06060_ _06068_ _06052_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__a31oi_4
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13136_ net1489 net575 net432 VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__mux2_1
XFILLER_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10348_ cpuregs\[9\]\[31\] net638 net612 _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__o211a_1
XANTENNA__10581__B2 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_930 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13537__S net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10279_ _04923_ _04924_ _04926_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__and3_1
XFILLER_97_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13067_ net584 net2277 net442 VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__mux2_1
XANTENNA__12322__A2 decoded_imm_j\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11565__B mem_rdata_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12018_ net1023 _06474_ net867 VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11530__A0 mem_rdata_q\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13969_ clknet_leaf_21_clk _00423_ VGND VGND VPWR VPWR cpuregs\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_139_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_139_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_100_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07490_ reg_pc\[23\] decoded_imm\[23\] VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__nand2_1
XANTENNA__10468__Y _05168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08593__C net1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15639_ clknet_leaf_0_clk _01975_ VGND VGND VPWR VPWR cpuregs\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09160_ net2124 net287 net502 VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11597__B1 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08111_ net1159 net1013 _03337_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__o21a_1
X_09091_ net1498 net283 net510 VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__mux2_1
XFILLER_148_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11520__S net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08042_ _03302_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__nand2_1
XANTENNA__09197__S net494 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold901 cpuregs\[5\]\[20\] VGND VGND VPWR VPWR net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 cpuregs\[25\]\[19\] VGND VGND VPWR VPWR net2226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _01425_ VGND VGND VPWR VPWR net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 cpuregs\[11\]\[7\] VGND VGND VPWR VPWR net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 cpuregs\[11\]\[21\] VGND VGND VPWR VPWR net2259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A2 net1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold956 cpuregs\[11\]\[15\] VGND VGND VPWR VPWR net2270 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__B1 net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold967 instr_addi VGND VGND VPWR VPWR net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 cpuregs\[19\]\[4\] VGND VGND VPWR VPWR net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 cpuregs\[13\]\[26\] VGND VGND VPWR VPWR net2303 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net1152 _04763_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__nor2_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08944_ genblk1.genblk1.pcpi_mul.rd\[10\] genblk1.genblk1.pcpi_mul.rd\[42\] net954
+ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__mux2_1
Xhold1601 genblk1.genblk1.pcpi_mul.next_rs2\[47\] VGND VGND VPWR VPWR net2915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09714__B1 net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1612 genblk2.pcpi_div.quotient\[18\] VGND VGND VPWR VPWR net2926 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11521__A0 mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08875_ net904 _04207_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1623 genblk2.pcpi_div.quotient\[7\] VGND VGND VPWR VPWR net2937 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout473_A net474 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1634 genblk1.genblk1.pcpi_mul.next_rs2\[48\] VGND VGND VPWR VPWR net2948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1645 _01365_ VGND VGND VPWR VPWR net2959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1656 genblk1.genblk1.pcpi_mul.next_rs2\[18\] VGND VGND VPWR VPWR net2970 sky130_fd_sc_hd__dlygate4sd3_1
X_07826_ net1160 net1016 VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__or2_1
XFILLER_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1667 _00827_ VGND VGND VPWR VPWR net2981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1678 count_instr\[35\] VGND VGND VPWR VPWR net2992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1689 genblk1.genblk1.pcpi_mul.next_rs2\[29\] VGND VGND VPWR VPWR net3003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07740__A2 net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07757_ _03273_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout640_A net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout738_A net739 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13182__S net428 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08276__S net921 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07688_ cpuregs\[11\]\[3\] net623 net592 _03207_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__o211a_1
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09427_ count_instr\[7\] count_instr\[6\] _04313_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout905_A _03879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1170_X net1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09358_ net1584 net296 net477 VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08309_ net1188 _03738_ net983 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_23_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09289_ net2082 net298 net487 VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__mux2_1
XANTENNA__13211__A net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11320_ cpuregs\[16\]\[26\] net702 VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__or2_1
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12001__A1 net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11251_ net1080 decoded_imm\[24\] VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__nor2_1
XFILLER_134_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10202_ decoded_imm\[22\] net1007 VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__nand2_1
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11182_ cpuregs\[28\]\[23\] cpuregs\[29\]\[23\] net697 VGND VGND VPWR VPWR _05859_
+ sky130_fd_sc_hd__mux2_1
X_10133_ _04853_ net1229 _04851_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__and3b_1
XANTENNA__11666__A mem_rdata_q\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10064_ _04808_ _04809_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input34_A resetn VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14941_ clknet_leaf_8_clk _01293_ VGND VGND VPWR VPWR cpuregs\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_94_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14872_ clknet_leaf_6_clk _01224_ VGND VGND VPWR VPWR cpuregs\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07192__B1 net842 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_0_clk _00277_ VGND VGND VPWR VPWR cpuregs\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12068__A1 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12497__A net240 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13092__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13754_ clknet_leaf_3_clk _00208_ VGND VGND VPWR VPWR cpuregs\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_10966_ cpuregs\[14\]\[17\] cpuregs\[15\]\[17\] net655 VGND VGND VPWR VPWR _05649_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12705_ net1491 net897 _02086_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__a21o_1
X_13685_ clknet_leaf_115_clk _00139_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_10897_ cpuregs\[28\]\[15\] cpuregs\[29\]\[15\] net646 VGND VGND VPWR VPWR _05582_
+ sky130_fd_sc_hd__mux2_1
X_15424_ clknet_leaf_52_clk _01763_ VGND VGND VPWR VPWR cpuregs\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12636_ net2890 net890 _02067_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__a21o_1
XFILLER_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15355_ clknet_leaf_93_clk _01695_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfxtp_1
X_12567_ _02047_ net2634 net389 VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__mux2_1
XFILLER_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12436__S net865 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14306_ clknet_leaf_98_clk _00760_ VGND VGND VPWR VPWR count_cycle\[51\] sky130_fd_sc_hd__dfxtp_1
X_11518_ mem_rdata_q\[11\] net1782 net738 VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__mux2_1
X_15286_ clknet_leaf_15_clk _01627_ VGND VGND VPWR VPWR cpuregs\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_12498_ _05106_ net716 net240 VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__o21ai_1
Xhold208 cpuregs\[26\]\[7\] VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 cpuregs\[15\]\[10\] VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ clknet_leaf_177_clk _00691_ VGND VGND VPWR VPWR reg_next_pc\[14\] sky130_fd_sc_hd__dfxtp_1
X_11449_ net805 _06116_ _06118_ net833 VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_78_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12543__A2 net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14168_ clknet_leaf_126_clk _00622_ VGND VGND VPWR VPWR count_instr\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_140_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10554__A1 net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13119_ net321 net2276 net436 VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ genblk2.pcpi_div.quotient\[9\] genblk2.pcpi_div.quotient\[10\] _02556_ VGND
+ VGND VPWR VPWR _02565_ sky130_fd_sc_hd__or3_1
X_14099_ clknet_leaf_25_clk _00553_ VGND VGND VPWR VPWR cpuregs\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_39_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07970__A2 net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08660_ _04025_ _04026_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07611_ net1188 net1069 _03132_ net1085 _03131_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__a221o_1
XFILLER_94_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12059__A1 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08591_ genblk1.genblk1.pcpi_mul.next_rs2\[18\] net1100 genblk1.genblk1.pcpi_mul.rd\[17\]
+ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__a21o_1
X_07542_ count_instr\[58\] net1133 net1137 count_instr\[26\] VGND VGND VPWR VPWR _03069_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_157_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10639__B net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06836__C net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07473_ net1066 net1009 _03004_ net1086 _03003_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__a221o_1
XANTENNA__07486__A1 net1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07486__B2 net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09212_ net1697 net340 net492 VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__mux2_1
XFILLER_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ net1683 net351 net500 VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06852__B net1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10778__D1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A _03831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09074_ net1745 net347 net508 VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__mux2_1
XFILLER_135_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10374__B _05079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08025_ _03360_ _03531_ _03465_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__a21o_1
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold720 cpuregs\[7\]\[20\] VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 cpuregs\[16\]\[30\] VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold742 cpuregs\[8\]\[15\] VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold753 cpuregs\[8\]\[5\] VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold764 cpuregs\[8\]\[26\] VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap483 _04291_ VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout590_A net592 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10545__A1 net829 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold775 genblk1.genblk1.pcpi_mul.next_rs1\[19\] VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold786 cpuregs\[15\]\[27\] VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13177__S net427 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold797 cpuregs\[16\]\[23\] VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ net1152 _04747_ _04748_ _04746_ net1185 VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__o311a_1
XFILLER_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1016_X net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08927_ net1467 _04240_ net945 VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__mux2_1
XFILLER_57_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11636__D mem_rdata_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_A _05134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1420 genblk2.pcpi_div.divisor\[5\] VGND VGND VPWR VPWR net2734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_X net476 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1431 count_cycle\[37\] VGND VGND VPWR VPWR net2745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 genblk2.pcpi_div.quotient_msk\[9\] VGND VGND VPWR VPWR net2756 sky130_fd_sc_hd__dlygate4sd3_1
X_08858_ genblk1.genblk1.pcpi_mul.next_rs2\[59\] net1108 genblk1.genblk1.pcpi_mul.rd\[58\]
+ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__a21o_1
Xhold1453 _06602_ VGND VGND VPWR VPWR net2767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1464 instr_bge VGND VGND VPWR VPWR net2778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09390__S net402 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1475 genblk1.genblk1.pcpi_mul.rd\[29\] VGND VGND VPWR VPWR net2789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1486 instr_sll VGND VGND VPWR VPWR net2800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_936 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07809_ _03325_ _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__and2_1
Xhold1497 genblk1.genblk1.pcpi_mul.mul_counter\[4\] VGND VGND VPWR VPWR net2811 sky130_fd_sc_hd__dlygate4sd3_1
X_08789_ _04129_ _04132_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__nand2_1
XANTENNA__11425__S net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10820_ cpuregs\[10\]\[13\] net652 VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_28_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13206__A _02384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09403__B net1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07204__A net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10751_ cpuregs\[6\]\[11\] cpuregs\[7\]\[11\] net666 VGND VGND VPWR VPWR _05440_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout810_X net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13470_ net1521 net341 net423 VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__mux2_1
X_10682_ cpuregs\[24\]\[9\] net671 VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__or2_1
X_12421_ net285 net1590 net473 VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__mux2_1
X_15140_ clknet_leaf_71_clk _01492_ VGND VGND VPWR VPWR cpuregs\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12352_ genblk1.genblk1.pcpi_mul.mul_counter\[0\] genblk1.genblk1.pcpi_mul.mul_counter\[3\]
+ genblk1.genblk1.pcpi_mul.mul_counter\[2\] genblk1.genblk1.pcpi_mul.mul_counter\[1\]
+ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__or4_1
XANTENNA__10284__B net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11981__B1 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11303_ cpuregs\[8\]\[26\] net703 VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__or2_1
XFILLER_126_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15071_ clknet_leaf_103_clk net2376 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12283_ net745 _06619_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__and2_1
XANTENNA__07874__A _03389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14022_ clknet_leaf_36_clk _00476_ VGND VGND VPWR VPWR cpuregs\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11234_ cpuregs\[6\]\[24\] cpuregs\[7\]\[24\] net699 VGND VGND VPWR VPWR _05910_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11733__B1 _06243_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13087__S net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12930__C1 net710 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07401__A1 net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11165_ cpuregs\[25\]\[22\] net633 net610 _05842_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__o211a_1
XFILLER_96_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ _04841_ _04842_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__nor2_1
XANTENNA__12289__A1 mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11096_ cpuregs\[14\]\[20\] cpuregs\[15\]\[20\] net657 VGND VGND VPWR VPWR _05776_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output238_A net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10047_ count_cycle\[18\] count_cycle\[19\] _04791_ _04795_ VGND VGND VPWR VPWR _04798_
+ sky130_fd_sc_hd__and4_1
X_14924_ clknet_leaf_48_clk _01276_ VGND VGND VPWR VPWR cpuregs\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold80 cpuregs\[28\]\[5\] VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 decoded_rd\[4\] VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07704__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14855_ clknet_leaf_30_clk _01207_ VGND VGND VPWR VPWR cpuregs\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13806_ clknet_leaf_36_clk _00260_ VGND VGND VPWR VPWR cpuregs\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14786_ clknet_leaf_91_clk _01139_ VGND VGND VPWR VPWR mem_state\[0\] sky130_fd_sc_hd__dfxtp_1
X_11998_ _06340_ _06341_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13737_ clknet_leaf_108_clk _00191_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10949_ cpuregs\[26\]\[16\] net656 VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__or2_1
XANTENNA__10178__C _04883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13550__S net418 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13668_ clknet_leaf_144_clk _00122_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_15407_ clknet_leaf_194_clk _01746_ VGND VGND VPWR VPWR cpuregs\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_12619_ net1195 genblk1.genblk1.pcpi_mul.next_rs2\[9\] net915 net1168 VGND VGND VPWR
+ VPWR _02059_ sky130_fd_sc_hd__a22o_1
XANTENNA__07768__B net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13599_ clknet_leaf_27_clk _00054_ VGND VGND VPWR VPWR cpuregs\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15338_ clknet_leaf_166_clk _01678_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15269_ clknet_leaf_176_clk _01610_ VGND VGND VPWR VPWR cpuregs\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout507 _04279_ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__buf_4
X_09830_ decoded_imm_j\[17\] _04438_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__xnor2_1
Xfanout518 net519 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkbuf_8
Xfanout529 _03746_ VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__buf_2
XFILLER_59_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07943__A2 net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09761_ _04432_ _04540_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__or2_1
X_06973_ net1120 _02550_ genblk2.pcpi_div.quotient\[8\] VGND VGND VPWR VPWR _02551_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_79_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08712_ _04069_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11488__C1 net1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09692_ _04423_ _04424_ _04425_ _04426_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__a31o_1
XANTENNA__07156__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08643_ genblk1.genblk1.pcpi_mul.next_rs2\[26\] net1105 genblk1.genblk1.pcpi_mul.rd\[25\]
+ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__a21o_1
XANTENNA__13229__B1 net396 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07950__C net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08574_ _03952_ _03953_ _03947_ _03950_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_124_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07525_ count_instr\[25\] net1137 net979 _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__a211o_1
XFILLER_23_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07459__A1 net1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout1080_A net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13460__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_A net438 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1178_A net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10463__B1 net611 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07456_ genblk1.genblk1.pcpi_mul.pcpi_rd\[20\] genblk2.pcpi_div.pcpi_rd\[20\] net1112
+ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__mux2_1
XFILLER_168_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07311__X _02853_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07678__B net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_A net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07387_ _02922_ _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__nand2_1
XANTENNA__13401__B1 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09126_ latched_rd\[4\] latched_rd\[3\] VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2_1
XANTENNA__10766__A1 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09057_ net284 net2514 net515 VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__mux2_1
XANTENNA__07631__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12804__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09385__S net399 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08008_ _03354_ _03516_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__or2_1
XANTENNA__12507__A2 net718 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold550 cpuregs\[24\]\[18\] VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout593_X net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold561 cpuregs\[31\]\[20\] VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout972_A net975 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold572 cpuregs\[25\]\[16\] VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 cpuregs\[29\]\[7\] VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 cpuregs\[31\]\[28\] VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09959_ net1129 _04448_ _04726_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout760_X net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12970_ net1874 net582 net449 VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1250 reg_next_pc\[22\] VGND VGND VPWR VPWR net2564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 genblk1.genblk1.pcpi_mul.next_rs1\[28\] VGND VGND VPWR VPWR net2575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11921_ genblk2.pcpi_div.divisor\[47\] genblk2.pcpi_div.divisor\[46\] genblk2.pcpi_div.divisor\[45\]
+ genblk2.pcpi_div.divisor\[44\] VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__or4_1
Xhold1272 reg_next_pc\[29\] VGND VGND VPWR VPWR net2586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1283 reg_next_pc\[27\] VGND VGND VPWR VPWR net2597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 instr_sra VGND VGND VPWR VPWR net2608 sky130_fd_sc_hd__dlygate4sd3_1
X_14640_ clknet_leaf_164_clk _01025_ VGND VGND VPWR VPWR genblk2.pcpi_div.dividend\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_11852_ _06319_ _06322_ _06317_ _06318_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__o211a_1
XFILLER_61_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10803_ net772 _05466_ _05474_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__a31oi_4
X_14571_ clknet_leaf_51_clk _00957_ VGND VGND VPWR VPWR cpuregs\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11246__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11783_ _04299_ _06255_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_52_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08111__A2 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13522_ net583 net1844 net417 VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__mux2_1
X_10734_ net1166 net853 _05422_ _05423_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__a22o_1
XANTENNA__06773__A net1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13453_ net992 net394 _02352_ _02354_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10665_ _05354_ _05355_ net813 VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__mux2_1
XFILLER_139_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12404_ net352 net1879 net471 VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13384_ reg_pc\[22\] _05079_ _05855_ is_lui_auipc_jal VGND VGND VPWR VPWR _02294_
+ sky130_fd_sc_hd__o2bb2a_1
X_10596_ cpuregs\[12\]\[7\] cpuregs\[13\]\[7\] net673 VGND VGND VPWR VPWR _05289_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15123_ clknet_leaf_184_clk _01475_ VGND VGND VPWR VPWR cpuregs\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ decoded_imm\[7\] net735 _06643_ mem_rdata_q\[27\] _06647_ VGND VGND VPWR
+ VPWR _01167_ sky130_fd_sc_hd__a221o_1
XANTENNA__07622__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15054_ clknet_leaf_102_clk net2473 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11397__Y _06069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12266_ net2873 net380 net368 net2891 VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__a22o_1
XFILLER_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10509__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14005_ clknet_leaf_190_clk _00459_ VGND VGND VPWR VPWR cpuregs\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11217_ cpuregs\[30\]\[24\] cpuregs\[31\]\[24\] net697 VGND VGND VPWR VPWR _05893_
+ sky130_fd_sc_hd__mux2_1
X_12197_ genblk2.pcpi_div.quotient_msk\[12\] net271 net2961 VGND VGND VPWR VPWR _06591_
+ sky130_fd_sc_hd__a21oi_1
Xoutput70 net70 VGND VGND VPWR VPWR mem_la_addr[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput81 net81 VGND VGND VPWR VPWR mem_la_addr[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput92 net92 VGND VGND VPWR VPWR mem_la_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11148_ cpuregs\[2\]\[22\] cpuregs\[3\]\[22\] net683 VGND VGND VPWR VPWR _05826_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13545__S net418 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11079_ cpuregs\[20\]\[20\] cpuregs\[21\]\[20\] net657 VGND VGND VPWR VPWR _05759_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07138__B1 net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07689__A1 net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14907_ clknet_leaf_142_clk _01259_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14838_ clknet_leaf_0_clk _01190_ VGND VGND VPWR VPWR cpuregs\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10189__B net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14769_ clknet_leaf_164_clk _00023_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_07310_ net20 _02689_ _02694_ net3 _02812_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__o221a_1
XANTENNA__09330__Y _04292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08374__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08290_ reg_out\[22\] reg_next_pc\[22\] net926 VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07241_ net1064 net1038 _02787_ net1078 _02786_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__a221o_1
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07172_ reg_pc\[2\] decoded_imm\[2\] VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__nand2_1
XFILLER_11_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11945__B1 net866 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07613__A1 net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout304 _03849_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout315 _03836_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout326 net327 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
X_09813_ _04586_ _04436_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__and2b_1
Xfanout337 _03810_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_2
Xfanout348 _03799_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_2
XFILLER_113_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout359 _02914_ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13455__S net426 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09744_ _04534_ _04535_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__nand2_1
X_06956_ genblk2.pcpi_div.quotient\[6\] _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_126_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ _04463_ _04467_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__nand2_1
X_06887_ _02482_ _00814_ _02484_ _02445_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout553_A _03156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08626_ _03996_ _03997_ _03991_ _03994_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__a211o_1
XFILLER_70_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08557_ net1193 net2911 net886 _03939_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__a22o_1
XFILLER_42_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout341_X net341 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout439_X net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net821 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13190__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11703__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07508_ _03033_ _03036_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__or2_1
XANTENNA__08284__S net922 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08488_ genblk1.genblk1.pcpi_mul.next_rs2\[2\] net1101 genblk1.genblk1.pcpi_mul.rd\[1\]
+ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__a21oi_1
X_07439_ net1065 net1012 _02972_ net1078 _02971_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a221o_1
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_X net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11004__A net809 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10450_ net834 _05145_ _05147_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a211o_1
X_09109_ net1475 net339 net504 VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__mux2_1
XANTENNA__11939__A net1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10381_ genblk2.pcpi_div.quotient_msk\[7\] genblk2.pcpi_div.quotient_msk\[6\] genblk2.pcpi_div.quotient_msk\[5\]
+ genblk2.pcpi_div.quotient_msk\[4\] VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__or4_1
XANTENNA__12534__S net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12120_ net3033 net274 _06562_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09409__A net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_X net975 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12051_ net722 _06501_ net1013 VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__a21oi_1
Xhold380 cpuregs\[14\]\[16\] VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 cpuregs\[8\]\[14\] VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11002_ cpuregs\[12\]\[18\] cpuregs\[13\]\[18\] net647 VGND VGND VPWR VPWR _05684_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07907__A2 net228 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout860 _05133_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__buf_4
XANTENNA__10911__B2 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout871 net872 VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__clkbuf_2
Xfanout882 _04421_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__buf_2
Xfanout893 net898 VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__buf_2
X_12953_ net331 net1951 net452 VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__mux2_1
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1080 cpuregs\[9\]\[6\] VGND VGND VPWR VPWR net2394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 cpuregs\[11\]\[3\] VGND VGND VPWR VPWR net2405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11904_ _06373_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__nand2_1
X_12884_ mem_rdata_q\[21\] net14 net962 VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__mux2_1
XFILLER_93_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14623_ clknet_leaf_109_clk net1371 VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_wait
+ sky130_fd_sc_hd__dfxtp_1
X_11835_ genblk2.pcpi_div.divisor\[9\] genblk2.pcpi_div.dividend\[9\] VGND VGND VPWR
+ VPWR _06306_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_25_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_16_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ clknet_leaf_192_clk _00940_ VGND VGND VPWR VPWR cpuregs\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11766_ net1479 net121 net728 VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__mux2_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ net1839 net334 net419 VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _05405_ _05406_ net802 VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__mux2_1
X_14485_ clknet_leaf_95_clk _00874_ VGND VGND VPWR VPWR instr_xori sky130_fd_sc_hd__dfxtp_1
X_11697_ net1978 net348 net373 VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__mux2_1
XFILLER_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13436_ reg_pc\[28\] _05079_ _02339_ _04880_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__a211o_1
X_10648_ cpuregs\[26\]\[8\] net670 VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__or2_1
XFILLER_155_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11388__D1 net793 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13367_ net1012 net755 net558 _02255_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__o211a_1
X_10579_ cpuregs\[17\]\[6\] net627 net608 _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__o211a_1
XFILLER_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07538__S net1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15106_ clknet_leaf_33_clk _01458_ VGND VGND VPWR VPWR cpuregs\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12318_ net1146 decoded_imm_j\[14\] net970 mem_rdata_q\[14\] VGND VGND VPWR VPWR
+ _06638_ sky130_fd_sc_hd__a22o_1
X_13298_ _02407_ net753 VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__nand2_1
XFILLER_114_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15037_ clknet_leaf_135_clk _01389_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_12249_ genblk2.pcpi_div.divisor\[12\] net379 net366 net2677 VGND VGND VPWR VPWR
+ _01118_ sky130_fd_sc_hd__a22o_1
XFILLER_170_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07359__B1 net1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10899__S net796 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06810_ mem_state\[0\] mem_state\[1\] VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__nor2_1
XANTENNA__07781__B net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08369__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07790_ net1172 net1040 VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__nand2_1
XFILLER_111_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12655__B2 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09460_ count_instr\[18\] count_instr\[15\] _04330_ _04336_ VGND VGND VPWR VPWR _04338_
+ sky130_fd_sc_hd__and4_1
X_08411_ reg_pc\[18\] _03813_ reg_pc\[19\] VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_121_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09391_ net1963 net295 net401 VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__mux2_1
XANTENNA__10928__A net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11523__S net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09060__Y _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13304__A _02408_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08342_ _03763_ _03764_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__nor2_1
XANTENNA__15499__Q net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08273_ net1024 _03720_ net980 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__mux2_1
XFILLER_149_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09036__A0 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07224_ net1065 net1040 _02771_ net1078 _02770_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__a221o_1
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07956__B net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07155_ _02383_ net18 _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout301_A _03849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07598__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07086_ net1121 _02647_ genblk2.pcpi_div.dividend\[24\] VGND VGND VPWR VPWR _02648_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_160_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09339__A1 net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1210_A net1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08011__A1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08011__B2 net928 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12894__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06859__Y _02462_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13185__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout389_X net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07988_ net968 _03282_ net934 _03280_ _03499_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__o221a_1
XANTENNA__08279__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09727_ net846 _04519_ _04520_ net876 net2256 VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__a32o_1
X_06939_ genblk2.pcpi_div.dividend\[3\] net1126 _02520_ net949 VGND VGND VPWR VPWR
+ _02522_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout935_A _03459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09658_ decoded_imm_j\[1\] _04422_ _04457_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__a21o_1
XFILLER_70_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ net1203 net2888 net895 _03983_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__a22o_1
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout723_X net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09589_ net1089 net1207 VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__nor2_1
X_11620_ mem_rdata_q\[17\] mem_rdata_q\[16\] mem_rdata_q\[15\] mem_rdata_q\[2\] VGND
+ VGND VPWR VPWR _06209_ sky130_fd_sc_hd__or4_1
XANTENNA__08078__A1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11551_ net1209 net746 VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__nor2_1
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08027__B net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09027__A0 _03749_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10502_ cpuregs\[18\]\[1\] net554 _05200_ net783 VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__o22a_1
XFILLER_156_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14270_ clknet_leaf_129_clk _00724_ VGND VGND VPWR VPWR count_cycle\[15\] sky130_fd_sc_hd__dfxtp_1
X_11482_ net1072 net1089 VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__or2_1
XFILLER_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13221_ _02144_ _02146_ _02150_ net397 net1045 VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__o32a_1
XANTENNA__11669__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10433_ net1083 net1088 net1231 VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__o21a_1
XFILLER_109_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12582__A0 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13152_ net1625 net325 net433 VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__mux2_1
X_10364_ cpuregs\[24\]\[31\] net693 VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__or2_1
XFILLER_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12103_ _06375_ _06546_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__or2_1
XFILLER_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13083_ net334 net1815 net439 VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__mux2_1
X_10295_ decoded_imm\[18\] net1014 VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__nand2_1
XFILLER_78_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_155_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12034_ net861 _06358_ _06488_ _06487_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__a31o_1
XANTENNA__12885__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13095__S net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09750__A1 net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10896__B1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09750__B2 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout690 net691 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output220_A net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13985_ clknet_leaf_42_clk _00439_ VGND VGND VPWR VPWR cpuregs\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12637__B2 net1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12936_ net585 net2415 net453 VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__mux2_1
XFILLER_61_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ net27 net2936 _02450_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_164_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14606_ clknet_leaf_156_clk _00992_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dfxtp_1
X_11818_ _02360_ genblk2.pcpi_div.dividend\[16\] _06288_ VGND VGND VPWR VPWR _06289_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__08069__A1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13062__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15586_ clknet_leaf_53_clk _01922_ VGND VGND VPWR VPWR cpuregs\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12798_ net588 net1938 net465 VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ clknet_leaf_88_clk _00925_ VGND VGND VPWR VPWR is_jalr_addi_slti_sltiu_xori_ori_andi
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11749_ net1890 net102 net727 VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__mux2_1
X_14468_ clknet_leaf_93_clk _00857_ VGND VGND VPWR VPWR instr_beq sky130_fd_sc_hd__dfxtp_1
X_13419_ _02319_ _02320_ _02324_ net398 net1000 VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__o32a_1
X_14399_ clknet_leaf_99_clk _00820_ VGND VGND VPWR VPWR pcpi_timeout_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08241__A1 net251 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08960_ genblk1.genblk1.pcpi_mul.rd\[18\] genblk1.genblk1.pcpi_mul.rd\[50\] net955
+ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12902__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12325__B1 decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07911_ net1171 net1039 VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12876__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08891_ genblk1.genblk1.pcpi_mul.rd\[63\] _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__xor2_1
XANTENNA__11518__S net738 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07842_ _03357_ _03359_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__nand2_2
XANTENNA__10887__B1 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07773_ _03289_ _03290_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__and2_1
XFILLER_37_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09512_ count_instr\[36\] count_instr\[35\] _04363_ _04368_ VGND VGND VPWR VPWR _04372_
+ sky130_fd_sc_hd__and4_1
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07911__A_N net1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09443_ net3065 _04325_ net1226 VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout349_A _03799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09374_ net1920 net406 net400 VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__mux2_1
XANTENNA__13053__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11064__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08325_ net584 net2523 net530 VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__mux2_1
XFILLER_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout516_A net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1160_A net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08256_ reg_out\[5\] reg_next_pc\[5\] net923 VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__mux2_1
X_07207_ net1065 net1042 _02755_ net1079 VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__a22o_1
X_08187_ net1145 _03675_ _03676_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10393__A net1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12564__B1 net719 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07178__S net1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08232__A1 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07138_ net1048 net31 net1057 net1052 VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__o211a_1
XANTENNA__08232__B2 _02690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07069_ net950 _02629_ _02630_ _02632_ _02633_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__o32a_1
XANTENNA__12812__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput260 net260 VGND VGND VPWR VPWR pcpi_rs2[3] sky130_fd_sc_hd__buf_2
XFILLER_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12316__B1 net970 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09393__S net402 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10080_ count_cycle\[29\] count_cycle\[30\] _04816_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__and3_1
XFILLER_0_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout840_X net840 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12619__B2 net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13770_ clknet_leaf_52_clk _00224_ VGND VGND VPWR VPWR cpuregs\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10982_ net822 _05660_ _05662_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__a211o_1
XFILLER_56_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11671__B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ net1335 net883 _02094_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__a21o_1
XFILLER_71_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_154_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11163__S net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15440_ clknet_leaf_3_clk _01779_ VGND VGND VPWR VPWR cpuregs\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_12652_ net1210 net2724 net900 net2971 _02075_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__a221o_1
XANTENNA__13044__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11603_ net1234 mem_rdata_q\[30\] is_alu_reg_reg _06199_ VGND VGND VPWR VPWR _06202_
+ sky130_fd_sc_hd__and4_1
XANTENNA__11055__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15371_ clknet_leaf_20_clk _01710_ VGND VGND VPWR VPWR cpuregs\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12583_ net403 net2023 net467 VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__mux2_1
XFILLER_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_169_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14322_ clknet_leaf_130_clk _06738_ VGND VGND VPWR VPWR reg_out\[2\] sky130_fd_sc_hd__dfxtp_1
X_11534_ mem_rdata_q\[27\] net2875 net736 VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__mux2_1
XANTENNA__07877__A _03368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07274__A2 net1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14771__Q genblk2.pcpi_div.pcpi_rd\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14253_ clknet_leaf_66_clk _00707_ VGND VGND VPWR VPWR reg_next_pc\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11465_ cpuregs\[30\]\[30\] cpuregs\[31\]\[30\] net690 VGND VGND VPWR VPWR _06135_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13204_ net1051 net397 _02130_ _02135_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__o22a_1
XFILLER_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10416_ net1157 _05119_ _05120_ net389 net2455 VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__a32o_1
X_14184_ clknet_leaf_102_clk _00638_ VGND VGND VPWR VPWR count_instr\[55\] sky130_fd_sc_hd__dfxtp_1
X_11396_ net832 _06063_ _06065_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__a211o_1
X_13135_ net1444 net579 net433 VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__mux2_1
X_10347_ cpuregs\[8\]\[31\] net694 VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__or2_1
XFILLER_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10581__A2 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13066_ net586 net2161 net441 VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__mux2_1
X_10278_ _04925_ _04983_ _04926_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12017_ net1025 _06470_ net721 VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__o21a_1
XFILLER_78_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11565__C mem_rdata_q\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07734__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11677__D_N net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13283__A1 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13968_ clknet_leaf_28_clk _00422_ VGND VGND VPWR VPWR cpuregs\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12919_ net309 net2471 net456 VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__mux2_1
X_13899_ clknet_leaf_66_clk _00353_ VGND VGND VPWR VPWR cpuregs\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11073__S net810 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13035__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15638_ clknet_leaf_10_clk _01974_ VGND VGND VPWR VPWR cpuregs\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15569_ clknet_leaf_193_clk _01905_ VGND VGND VPWR VPWR cpuregs\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08110_ _03336_ _03339_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__nand2_1
XFILLER_119_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07787__A net1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09090_ net1545 net285 net511 VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__mux2_1
XANTENNA__08235__X net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08041_ _03432_ _03546_ net988 VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 cpuregs\[18\]\[0\] VGND VGND VPWR VPWR net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 cpuregs\[3\]\[27\] VGND VGND VPWR VPWR net2227 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__A1 _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold924 net177 VGND VGND VPWR VPWR net2238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold935 cpuregs\[7\]\[7\] VGND VGND VPWR VPWR net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold946 cpuregs\[19\]\[20\] VGND VGND VPWR VPWR net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 cpuregs\[24\]\[19\] VGND VGND VPWR VPWR net2271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A3 net720 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold968 cpuregs\[17\]\[9\] VGND VGND VPWR VPWR net2282 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _04452_ _04758_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold979 genblk1.genblk1.pcpi_mul.next_rs1\[24\] VGND VGND VPWR VPWR net2293 sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ net1374 _04248_ net943 VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__mux2_1
XANTENNA__09507__A _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10660__B decoded_imm\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout299_A _03852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08874_ genblk1.genblk1.pcpi_mul.next_rs2\[61\] net1106 _04204_ _04206_ VGND VGND
+ VPWR VPWR _04208_ sky130_fd_sc_hd__and4_1
Xhold1602 _01353_ VGND VGND VPWR VPWR net2916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1613 genblk1.genblk1.pcpi_mul.rd\[55\] VGND VGND VPWR VPWR net2927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 genblk1.genblk1.pcpi_mul.next_rs2\[43\] VGND VGND VPWR VPWR net2938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07725__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1635 genblk1.genblk1.pcpi_mul.rd\[62\] VGND VGND VPWR VPWR net2949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1646 mem_state\[1\] VGND VGND VPWR VPWR net2960 sky130_fd_sc_hd__dlygate4sd3_1
X_07825_ _03341_ _03342_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__nor2_1
XFILLER_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1657 genblk1.genblk1.pcpi_mul.next_rs2\[24\] VGND VGND VPWR VPWR net2971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_A _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1668 count_instr\[3\] VGND VGND VPWR VPWR net2982 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13463__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1679 genblk1.genblk1.pcpi_mul.next_rs2\[13\] VGND VGND VPWR VPWR net2993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07756_ net1176 net1044 VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__nor2_1
XANTENNA__10659__Y _05351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07314__X _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12079__S net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07687_ cpuregs\[10\]\[3\] net661 VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__or2_1
XANTENNA__12478__B1_N net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A net635 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09426_ _04314_ _04315_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__nor2_1
X_09357_ net1562 net299 net478 VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout421_X net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12807__S net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout800_A net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1163_X net1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11711__S net376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout519_X net519 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08308_ reg_out\[31\] reg_next_pc\[31\] net924 VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09388__S net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08292__S net926 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09288_ net1721 net302 net487 VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__mux2_1
XFILLER_100_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08145__X alu_out\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10796__C1 net826 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08239_ net1171 net1158 net940 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__mux2_1
XFILLER_153_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11250_ _05916_ _05925_ _05909_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__a21oi_2
XFILLER_153_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12001__A2 net723 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout790_X net790 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10201_ decoded_imm\[23\] net218 VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__nor2_1
XANTENNA__11947__A net873 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11181_ cpuregs\[30\]\[23\] cpuregs\[31\]\[23\] net697 VGND VGND VPWR VPWR _05858_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12542__S net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10563__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07964__B1 net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10132_ count_cycle\[47\] _04846_ _04852_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__and3_1
XFILLER_79_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11666__B net745 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09705__A1 net1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10063_ net2996 _04806_ net1236 VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__o21ai_1
X_14940_ clknet_leaf_6_clk _01292_ VGND VGND VPWR VPWR cpuregs\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__09705__B2 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input27_A mem_rdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14871_ clknet_leaf_18_clk _01223_ VGND VGND VPWR VPWR cpuregs\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_13822_ clknet_leaf_10_clk _00276_ VGND VGND VPWR VPWR cpuregs\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08467__S net531 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__06776__A net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13753_ clknet_leaf_194_clk _00207_ VGND VGND VPWR VPWR cpuregs\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11276__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10965_ cpuregs\[12\]\[17\] cpuregs\[13\]\[17\] net655 VGND VGND VPWR VPWR _05648_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12704_ net1191 genblk1.genblk1.pcpi_mul.next_rs1\[1\] net916 net1046 VGND VGND VPWR
+ VPWR _02086_ sky130_fd_sc_hd__a22o_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13684_ clknet_leaf_115_clk _00138_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_10896_ net787 _05576_ _05578_ _05580_ net776 VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__o41a_1
X_15423_ clknet_leaf_50_clk _01762_ VGND VGND VPWR VPWR cpuregs\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12635_ net1196 genblk1.genblk1.pcpi_mul.next_rs2\[17\] net914 net1161 VGND VGND
+ VPWR VPWR _02067_ sky130_fd_sc_hd__a22o_1
XFILLER_157_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09298__S net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15354_ clknet_leaf_62_clk _01694_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfxtp_1
XFILLER_156_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12566_ genblk2.pcpi_div.divisor\[61\] _02046_ net874 VGND VGND VPWR VPWR _02047_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12240__A2 net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11517_ mem_rdata_q\[10\] net2042 net737 VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__mux2_1
X_14305_ clknet_leaf_110_clk _00759_ VGND VGND VPWR VPWR count_cycle\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09671__A2_N _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15285_ clknet_leaf_41_clk _01626_ VGND VGND VPWR VPWR cpuregs\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12497_ net240 _05106_ net715 VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_150_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output95_A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14236_ clknet_leaf_177_clk _00690_ VGND VGND VPWR VPWR reg_next_pc\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold209 cpuregs\[31\]\[24\] VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ net817 _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08930__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13548__S net417 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14167_ clknet_leaf_126_clk _00621_ VGND VGND VPWR VPWR count_instr\[38\] sky130_fd_sc_hd__dfxtp_1
X_11379_ net793 _06046_ _06048_ _06050_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__or4_1
XFILLER_4_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13118_ net325 net2424 net437 VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ clknet_leaf_24_clk _00552_ VGND VGND VPWR VPWR cpuregs\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13049_ net1623 net72 net534 VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11592__A mem_rdata_q\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07610_ genblk1.genblk1.pcpi_mul.pcpi_rd\[31\] genblk2.pcpi_div.pcpi_rd\[31\] net1112
+ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__mux2_1
XFILLER_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10700__S net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08590_ net890 _03965_ _03967_ net2567 net1196 VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__a32o_1
XANTENNA__06930__A1 net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11267__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07541_ net1073 _03061_ _03062_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_157_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08683__A1 genblk1.genblk1.pcpi_mul.next_rs2\[32\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07472_ genblk1.genblk1.pcpi_mul.pcpi_rd\[21\] genblk2.pcpi_div.pcpi_rd\[21\] net1112
+ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__mux2_1
XANTENNA__07486__A2 net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09880__B1 net881 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09211_ net1841 net343 net492 VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__mux2_1
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09142_ net1652 net354 net501 VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12231__A2 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09001__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09073_ net1552 net350 net508 VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__mux2_1
XANTENNA__06997__A1 net948 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08024_ _03360_ _03531_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__nor2_1
XFILLER_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11990__B2 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold710 cpuregs\[3\]\[13\] VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 cpuregs\[3\]\[26\] VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 cpuregs\[4\]\[3\] VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13458__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold743 cpuregs\[19\]\[21\] VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10671__A net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold754 cpuregs\[6\]\[20\] VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12362__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1123_A net1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold765 cpuregs\[27\]\[1\] VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A1 net1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold776 cpuregs\[8\]\[27\] VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 net181 VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07456__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09975_ _04450_ _04736_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__and2_1
Xhold798 cpuregs\[2\]\[21\] VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout583_A _03751_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08926_ genblk1.genblk1.pcpi_mul.rd\[1\] genblk1.genblk1.pcpi_mul.rd\[33\] net957
+ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__mux2_1
XFILLER_131_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1410 genblk1.genblk1.pcpi_mul.next_rs2\[25\] VGND VGND VPWR VPWR net2724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_X net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1421 genblk2.pcpi_div.quotient\[17\] VGND VGND VPWR VPWR net2735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1432 genblk2.pcpi_div.quotient\[0\] VGND VGND VPWR VPWR net2746 sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ net901 _04191_ _04193_ net2878 net1213 VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__a32o_1
Xhold1443 _01050_ VGND VGND VPWR VPWR net2757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout371_X net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net751 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1454 reg_sh\[2\] VGND VGND VPWR VPWR net2768 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13193__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net852 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11706__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1465 count_instr\[14\] VGND VGND VPWR VPWR net2779 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ net250 net1006 VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__or2_1
Xhold1476 count_cycle\[9\] VGND VGND VPWR VPWR net2790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1487 genblk2.pcpi_div.quotient\[10\] VGND VGND VPWR VPWR net2801 sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ _04133_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__nand2_1
XFILLER_73_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08287__S net981 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1498 genblk2.pcpi_div.quotient\[19\] VGND VGND VPWR VPWR net2812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11258__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07739_ cpuregs\[16\]\[4\] net698 VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__or2_1
XANTENNA__13206__B net759 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10750_ net828 _05434_ _05436_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__a211o_1
XFILLER_81_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07204__B net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09409_ net1206 _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__nor2_1
X_10681_ _05370_ _05371_ net814 VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout803_X net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12537__S _05082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12758__B1 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13222__A _03227_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12420_ net291 net1966 net473 VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__mux2_1
XFILLER_166_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12351_ decoded_imm\[1\] net745 _06656_ _06657_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__o22a_1
XANTENNA__11430__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11302_ net807 _05973_ _05975_ net836 VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__o211a_1
X_15070_ clknet_leaf_103_clk _01422_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12282_ net1150 net1128 _06618_ mem_rdata_q\[31\] VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__a22o_1
XFILLER_154_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14021_ clknet_leaf_23_clk _00475_ VGND VGND VPWR VPWR cpuregs\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11677__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11233_ net775 _05900_ _05908_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__and3_1
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10536__A2 net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12930__B1 decoded_imm_j\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07219__X _02767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ cpuregs\[24\]\[22\] net683 VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__or2_1
XFILLER_150_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ net2860 _04840_ net1225 VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_73_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ cpuregs\[12\]\[20\] cpuregs\[13\]\[20\] net657 VGND VGND VPWR VPWR _05775_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10046_ _04797_ net1229 _04796_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__and3b_1
X_14923_ clknet_leaf_30_clk _01275_ VGND VGND VPWR VPWR cpuregs\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_output133_A net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07165__A1 net1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold70 cpuregs\[28\]\[29\] VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 cpuregs\[20\]\[22\] VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 decoded_rd\[2\] VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ clknet_leaf_50_clk _01206_ VGND VGND VPWR VPWR cpuregs\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13805_ clknet_leaf_49_clk _00259_ VGND VGND VPWR VPWR cpuregs\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11249__B1 net778 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14785_ clknet_leaf_98_clk _01138_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.instr_mulhu
+ sky130_fd_sc_hd__dfxtp_1
X_11997_ genblk2.pcpi_div.dividend\[10\] net271 _06455_ _06457_ VGND VGND VPWR VPWR
+ _01019_ sky130_fd_sc_hd__o22a_1
XFILLER_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13736_ clknet_leaf_107_clk _00190_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10948_ cpuregs\[25\]\[16\] net621 net605 _05631_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__o211a_1
XANTENNA__08925__S net945 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10879_ net1076 _05563_ net853 VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12447__S net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13667_ clknet_leaf_118_clk _00121_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15406_ clknet_leaf_193_clk _01745_ VGND VGND VPWR VPWR cpuregs\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07401__Y _02938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12618_ net2983 net888 _02058_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__a21o_1
X_13598_ clknet_leaf_21_clk _00053_ VGND VGND VPWR VPWR cpuregs\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11421__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15337_ clknet_leaf_166_clk _01677_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_1
X_12549_ genblk2.pcpi_div.divisor\[57\] _02033_ net874 VGND VGND VPWR VPWR _02034_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10775__A2 net619 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15268_ clknet_leaf_73_clk _01609_ VGND VGND VPWR VPWR cpuregs\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14219_ clknet_leaf_67_clk _00673_ VGND VGND VPWR VPWR reg_pc\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15199_ clknet_leaf_6_clk _01548_ VGND VGND VPWR VPWR cpuregs\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xfanout508 _04278_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkbuf_8
Xfanout519 _04274_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkbuf_4
X_09760_ _04516_ _04432_ _04431_ _04430_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__nand4b_1
XFILLER_101_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07943__A3 net933 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06972_ genblk2.pcpi_div.quotient\[7\] _02544_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__or2_1
XANTENNA__12910__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08711_ _04063_ _04066_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__nand2_1
X_09691_ _04423_ _04424_ _04425_ _04426_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__and4_2
XANTENNA__12685__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07156__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07156__B2 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11526__S net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1090 net1093 VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__buf_2
XFILLER_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08642_ net901 _04009_ _04011_ net2587 net1210 VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__a32o_1
XFILLER_55_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13229__B2 net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08573_ genblk1.genblk1.pcpi_mul.rd\[14\] genblk1.genblk1.pcpi_mul.next_rs2\[15\]
+ net1090 VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__nand3_1
XFILLER_82_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ count_instr\[57\] net1133 net1141 count_cycle\[57\] VGND VGND VPWR VPWR _03052_
+ sky130_fd_sc_hd__a22o_1
X_07455_ count_cycle\[20\] net974 net844 _02987_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout331_A _03818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A net430 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07386_ reg_pc\[16\] decoded_imm\[16\] VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__nand2_1
XANTENNA__13401__A1 net558 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09125_ net1865 net278 net506 VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__mux2_1
XFILLER_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout1240_A net1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09056_ net286 net2348 net514 VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__mux2_1
XFILLER_135_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07631__A2 decoded_imm_j\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08007_ _03354_ _03516_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout798_A net803 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13188__S net429 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold540 cpuregs\[27\]\[5\] VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold551 cpuregs\[21\]\[31\] VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold562 net160 VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold573 cpuregs\[21\]\[13\] VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold584 cpuregs\[25\]\[3\] VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 cpuregs\[27\]\[18\] VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07395__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12820__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09958_ net1129 _04449_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__xor2_1
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08909_ net1210 net2780 net899 _04231_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__a22o_1
XANTENNA__12676__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09889_ _04664_ _04668_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__or2_1
Xhold1240 net171 VGND VGND VPWR VPWR net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1251 reg_next_pc\[21\] VGND VGND VPWR VPWR net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 genblk1.genblk1.pcpi_mul.rd\[48\] VGND VGND VPWR VPWR net2576 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ genblk2.pcpi_div.divisor\[51\] genblk2.pcpi_div.divisor\[50\] genblk2.pcpi_div.divisor\[49\]
+ genblk2.pcpi_div.divisor\[48\] VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__or4_1
XFILLER_46_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1273 genblk1.genblk1.pcpi_mul.rd\[24\] VGND VGND VPWR VPWR net2587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 genblk1.genblk1.pcpi_mul.rd\[40\] VGND VGND VPWR VPWR net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 instr_blt VGND VGND VPWR VPWR net2609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11851_ _06320_ _06321_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__and2_1
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout920_X net920 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10802_ net779 _05480_ _05489_ net776 VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__o211a_1
XFILLER_122_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14570_ clknet_leaf_56_clk _00956_ VGND VGND VPWR VPWR cpuregs\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11782_ net175 net174 VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__nor2_1
XFILLER_13_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11651__A0 decoded_imm_j\[20\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10733_ net1076 _05421_ net853 VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__a21oi_1
X_13521_ net587 net2459 net417 VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__mux2_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11171__S net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13452_ _04879_ _02353_ net394 VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10664_ cpuregs\[4\]\[9\] cpuregs\[5\]\[9\] net666 VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10295__B net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12403_ net356 net2123 net471 VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__mux2_1
XANTENNA__11403__B1 net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13383_ net958 _05012_ _02288_ _02292_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__a31o_1
X_10595_ net829 _05283_ _05287_ net781 VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_11_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15122_ clknet_leaf_183_clk _01474_ VGND VGND VPWR VPWR cpuregs\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07083__B1 net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11954__B2 net873 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12334_ net1148 decoded_imm_j\[7\] net744 VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07622__A2 decoded_imm_j\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15053_ clknet_leaf_102_clk net2479 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12265_ genblk2.pcpi_div.divisor\[28\] net381 net369 net2873 VGND VGND VPWR VPWR
+ _01134_ sky130_fd_sc_hd__a22o_1
XFILLER_107_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10509__A2 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14004_ clknet_leaf_178_clk _00458_ VGND VGND VPWR VPWR cpuregs\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11216_ net250 net859 _05891_ _05892_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__a22o_1
XFILLER_107_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output250_A net250 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12196_ net749 net2714 VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__nor2_1
Xoutput60 net60 VGND VGND VPWR VPWR mem_addr[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput71 net71 VGND VGND VPWR VPWR mem_la_addr[15] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VGND VGND VPWR VPWR mem_la_addr[26] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VGND VGND VPWR VPWR mem_la_addr[7] sky130_fd_sc_hd__buf_2
X_11147_ _05823_ _05824_ net816 VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__mux2_1
XFILLER_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11078_ net824 _05753_ _05755_ _05757_ net788 VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__a2111o_1
XANTENNA__07138__A1 net1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14906_ clknet_leaf_121_clk _01258_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10029_ net2784 _04785_ net1224 VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10693__B2 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14837_ clknet_leaf_195_clk _01189_ VGND VGND VPWR VPWR cpuregs\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13561__S net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14768_ clknet_leaf_163_clk _00022_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07412__X _02948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11642__A0 decoded_imm_j\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13719_ clknet_leaf_151_clk _00173_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14699_ clknet_leaf_152_clk _01084_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11081__S net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07310__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07310__B2 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07240_ genblk1.genblk1.pcpi_mul.pcpi_rd\[6\] genblk2.pcpi_div.pcpi_rd\[6\] net1110
+ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__mux2_1
X_07171_ count_cycle\[2\] net971 net842 _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__o211a_1
XANTENNA__12905__S net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07795__A net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08390__S net1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout305 _03844_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_2
XFILLER_114_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout316 net319 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09812_ _02480_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__nand2_1
Xfanout327 _03823_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout338 _03810_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_2
Xfanout349 _03799_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_2
X_06955_ genblk2.pcpi_div.quotient\[4\] genblk2.pcpi_div.quotient\[5\] _02525_ net1125
+ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__o31a_1
X_09743_ decoded_imm_j\[10\] _04431_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_126_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout281_A _03873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12122__A1 net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net384 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11256__S net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09674_ net2651 net878 _04472_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a21o_1
X_06886_ _02437_ _02438_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_143_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11483__C _02387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08625_ genblk1.genblk1.pcpi_mul.rd\[22\] genblk1.genblk1.pcpi_mul.next_rs2\[23\]
+ net1103 VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__nand3_1
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout1190_A net1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13471__S net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _03741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08556_ _03937_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_59_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08629__A1 net903 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08418__X _03826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07507_ _03034_ _03035_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__nand2_1
XFILLER_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12087__S net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10396__A net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08487_ _03878_ net894 _03880_ net2681 net1199 VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout713_A _02083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08137__Y alu_out\[22\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07438_ genblk1.genblk1.pcpi_mul.pcpi_rd\[19\] genblk2.pcpi_div.pcpi_rd\[19\] net1111
+ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__mux2_1
XFILLER_50_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07369_ _02905_ _02906_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout501_X net501 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__06880__Y _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12815__S net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09108_ net1933 net343 net505 VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__mux2_1
XFILLER_136_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10380_ genblk2.pcpi_div.quotient_msk\[15\] genblk2.pcpi_div.quotient_msk\[14\] genblk2.pcpi_div.quotient_msk\[13\]
+ genblk2.pcpi_div.quotient_msk\[12\] VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__or4_1
XANTENNA__11939__B _02507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09039_ net353 net2298 net512 VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__mux2_1
XANTENNA__10335__S net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11149__C1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12050_ net1013 net722 _06501_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__and3_1
XFILLER_2_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold370 cpuregs\[25\]\[12\] VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08014__C1 net1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold381 cpuregs\[30\]\[9\] VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11001_ net838 _05680_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__o21a_1
Xhold392 cpuregs\[28\]\[3\] VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_X net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10372__A0 net999 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12550__S net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout850 net851 VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10911__A2 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout861 net862 VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__buf_2
Xfanout872 net873 VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__clkbuf_2
Xfanout883 net898 VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__buf_2
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout894 net896 VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__buf_2
XANTENNA__12113__B2 net869 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13310__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12952_ net334 net2178 net452 VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__mux2_1
XFILLER_85_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1070 cpuregs\[7\]\[24\] VGND VGND VPWR VPWR net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 cpuregs\[19\]\[24\] VGND VGND VPWR VPWR net2395 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ genblk2.pcpi_div.dividend\[26\] genblk2.pcpi_div.divisor\[26\] VGND VGND
+ VPWR VPWR _06374_ sky130_fd_sc_hd__nand2b_1
Xhold1092 cpuregs\[18\]\[23\] VGND VGND VPWR VPWR net2406 sky130_fd_sc_hd__dlygate4sd3_1
X_12883_ mem_rdata_q\[20\] net13 net964 VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__mux2_1
XFILLER_46_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14622_ clknet_leaf_108_clk _01008_ VGND VGND VPWR VPWR genblk2.pcpi_div.outsign
+ sky130_fd_sc_hd__dfxtp_1
X_11834_ genblk2.pcpi_div.dividend\[9\] genblk2.pcpi_div.divisor\[9\] VGND VGND VPWR
+ VPWR _06305_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_68_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06784__A net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10427__A1 _02489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14774__Q genblk2.pcpi_div.pcpi_rd\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14553_ clknet_leaf_187_clk _00939_ VGND VGND VPWR VPWR cpuregs\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11765_ net1791 net120 net728 VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__mux2_1
X_10716_ cpuregs\[30\]\[10\] cpuregs\[31\]\[10\] net669 VGND VGND VPWR VPWR _05406_
+ sky130_fd_sc_hd__mux2_1
X_13504_ net1885 net336 net419 VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14484_ clknet_leaf_95_clk _00873_ VGND VGND VPWR VPWR instr_sltiu sky130_fd_sc_hd__dfxtp_1
X_11696_ net2029 net351 net373 VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__mux2_1
XANTENNA__13377__B1 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13435_ is_lui_auipc_jal _06069_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__nor2_1
X_10647_ cpuregs\[25\]\[8\] net627 net608 _05338_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__o211a_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13366_ net1019 net755 _02277_ net710 VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__o211a_1
X_10578_ cpuregs\[16\]\[6\] net671 VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__or2_1
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15105_ clknet_leaf_22_clk _01457_ VGND VGND VPWR VPWR cpuregs\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12317_ net3063 net743 _06632_ _06637_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__o22a_1
XFILLER_114_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13297_ _02404_ net758 VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__nand2_1
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12248_ genblk2.pcpi_div.divisor\[11\] net379 net366 net2704 VGND VGND VPWR VPWR
+ _01117_ sky130_fd_sc_hd__a22o_1
X_15036_ clknet_leaf_135_clk net1338 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_147_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13556__S net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12179_ genblk2.pcpi_div.quotient_msk\[3\] net276 net2694 VGND VGND VPWR VPWR _06582_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07554__S net1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13301__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_160_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08410_ reg_out\[19\] alu_out_q\[19\] net1154 VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__mux2_1
XFILLER_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09390_ net2136 net300 net402 VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08385__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07142__X _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08341_ reg_pc\[5\] _03758_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__and2_1
XFILLER_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11105__A net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08272_ reg_out\[13\] reg_next_pc\[13\] net920 VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__mux2_1
XANTENNA__11091__A1 net798 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07223_ genblk1.genblk1.pcpi_mul.pcpi_rd\[5\] genblk2.pcpi_div.pcpi_rd\[5\] net1111
+ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__mux2_1
XANTENNA__07729__S net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12040__B1 net861 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07154_ net1048 net32 net1057 net1052 VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__o211a_1
XFILLER_146_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07085_ genblk2.pcpi_div.dividend\[23\] _02640_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1036_A net1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13466__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_A net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11775__A _06245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_A mem_rdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07987_ _03283_ net928 VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout663_A net679 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09726_ net1183 _04429_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__or2_1
X_06938_ genblk2.pcpi_div.outsign _02520_ genblk2.pcpi_div.dividend\[3\] VGND VGND
+ VPWR VPWR _02521_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06869_ net2912 _02460_ _02467_ net1057 _02470_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a221o_1
XANTENNA__10657__B2 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A _03137_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_X net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09657_ decoded_imm_j\[2\] _04423_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__xor2_1
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__06875__Y _02474_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11714__S net376 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08608_ _03981_ _03982_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__xnor2_1
X_09588_ net1940 _04418_ _04420_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08295__S net982 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08539_ genblk1.genblk1.pcpi_mul.next_rs2\[10\] net1095 genblk1.genblk1.pcpi_mul.rd\[9\]
+ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__a21o_1
XANTENNA__13214__B _03189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_X net716 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ net1152 net547 _06173_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_46_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13359__B1 net565 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10501_ cpuregs\[19\]\[1\] net636 net598 VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__o21a_1
XFILLER_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11481_ net1072 net1089 VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__nor2_1
XFILLER_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13230__A _03263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13220_ reg_pc\[2\] net565 _02148_ _02149_ net392 VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__a221o_1
XFILLER_155_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10432_ mem_do_wdata _05121_ _05132_ _02453_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__a22o_1
XANTENNA__11669__B net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12031__B1 net862 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13151_ net1493 net328 net431 VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__mux2_1
X_10363_ _05067_ _05068_ net817 VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__mux2_1
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12102_ _06375_ _06546_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__nand2_1
XFILLER_163_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13082_ net337 net2060 net440 VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__mux2_1
X_10294_ decoded_imm\[18\] net1014 VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__and2_1
XFILLER_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13531__A0 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12033_ _06291_ _06355_ _06357_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__nand3_1
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07882__B net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14769__Q genblk2.pcpi_div.pcpi_rd\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10896__A1 net787 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout680 net696 VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__buf_2
XFILLER_120_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout691 net696 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_2
X_13984_ clknet_leaf_0_clk _00438_ VGND VGND VPWR VPWR cpuregs\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input12_X net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09502__A2 _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12935_ net588 net2532 net453 VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__mux2_1
XANTENNA_output213_A net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ net26 net2793 _02450_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__mux2_1
X_14605_ clknet_leaf_118_clk _00991_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfxtp_1
X_11817_ genblk2.pcpi_div.divisor\[17\] genblk2.pcpi_div.dividend\[17\] VGND VGND
+ VPWR VPWR _06288_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_83_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ clknet_leaf_50_clk _01921_ VGND VGND VPWR VPWR cpuregs\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12797_ _03745_ _06663_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_32_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14536_ clknet_leaf_92_clk net2672 VGND VGND VPWR VPWR is_slli_srli_srai sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08933__S net944 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11748_ net1482 net101 net727 VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__mux2_1
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14467_ clknet_leaf_89_clk _00856_ VGND VGND VPWR VPWR instr_jal sky130_fd_sc_hd__dfxtp_2
XANTENNA__12455__S net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11679_ is_sb_sh_sw _06232_ net548 VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__mux2_1
X_13418_ net710 _02301_ _02321_ _02323_ net394 VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__a311o_1
X_14398_ clknet_leaf_99_clk _00819_ VGND VGND VPWR VPWR pcpi_timeout_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13349_ _02408_ net759 VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__nand2_1
XFILLER_143_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12325__A1 is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11595__A mem_rdata_q\[30\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07910_ _03283_ _03427_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__or2_1
X_15019_ clknet_leaf_122_clk net2410 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_08890_ net1107 genblk1.genblk1.pcpi_mul.rs2\[63\] VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__nand2_1
XFILLER_96_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07137__X net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07841_ net1166 net1029 VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__or2_1
X_07772_ net254 net998 VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__or2_1
XFILLER_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09511_ _04370_ _04371_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__nor2_1
XFILLER_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13315__A net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09442_ count_instr\[12\] _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__and2_1
XFILLER_25_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09004__S net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09373_ net2115 net409 net400 VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__mux2_1
XFILLER_80_898 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08128__B net932 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08324_ _03750_ reg_pc\[1\] net768 VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__mux2_4
XANTENNA__12261__B1 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08255_ net1042 _03711_ net981 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__mux2_2
XANTENNA__12365__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A _02358_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A _04278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07206_ genblk1.genblk1.pcpi_mul.pcpi_rd\[4\] genblk2.pcpi_div.pcpi_rd\[4\] net1111
+ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__mux2_1
XANTENNA__12013__B1 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08186_ net990 _03444_ _03446_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__or3_1
XANTENNA__10393__B net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12564__A1 net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07137_ _02689_ net942 _02443_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__a21bo_4
XANTENNA__08232__A2 net1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07068_ genblk2.pcpi_div.dividend\[21\] net1117 _02631_ net947 VGND VGND VPWR VPWR
+ _02633_ sky130_fd_sc_hd__a31o_1
XFILLER_160_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout780_A net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput250 net250 VGND VGND VPWR VPWR pcpi_rs2[23] sky130_fd_sc_hd__buf_2
XANTENNA__13196__S net430 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput261 net261 VGND VGND VPWR VPWR pcpi_rs2[4] sky130_fd_sc_hd__buf_2
XANTENNA__07991__A1 net988 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net882 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11709__S net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12316__B2 mem_rdata_q\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1206_X net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input4_X net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09406__C net1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_X net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07743__A1 net835 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09709_ _04502_ _04503_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__nand2b_1
X_10981_ cpuregs\[18\]\[17\] net552 _05663_ net779 VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__o22a_1
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout833_X net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12720_ net1190 genblk1.genblk1.pcpi_mul.next_rs1\[9\] net914 net1030 VGND VGND VPWR
+ VPWR _02094_ sky130_fd_sc_hd__a22o_1
XANTENNA__11671__C net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ _02396_ net913 VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__nor2_1
XFILLER_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11602_ net2400 net563 _06175_ _06201_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__a22o_1
XANTENNA__12252__B1 net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12582_ net408 net2402 net468 VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__mux2_1
X_15370_ clknet_leaf_180_clk _01709_ VGND VGND VPWR VPWR cpuregs\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10802__A1 net779 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14321_ clknet_leaf_131_clk _06727_ VGND VGND VPWR VPWR reg_out\[1\] sky130_fd_sc_hd__dfxtp_1
X_11533_ mem_rdata_q\[26\] net2684 net736 VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__mux2_1
XFILLER_156_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11464_ cpuregs\[28\]\[30\] cpuregs\[29\]\[30\] net690 VGND VGND VPWR VPWR _06134_
+ sky130_fd_sc_hd__mux2_1
X_14252_ clknet_leaf_66_clk _00706_ VGND VGND VPWR VPWR reg_next_pc\[29\] sky130_fd_sc_hd__dfxtp_1
X_10415_ net1214 _05083_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__nor2_2
X_13203_ net755 _02134_ _02132_ net393 VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__a211o_1
X_14183_ clknet_leaf_102_clk _00637_ VGND VGND VPWR VPWR count_instr\[54\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08223__A2 net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11395_ cpuregs\[18\]\[28\] net554 _06066_ net783 VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__o22a_1
XANTENNA__10566__B1 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10346_ net817 _05049_ _05051_ net833 VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__o211a_1
XFILLER_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13134_ net1484 net583 net433 VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__mux2_1
XANTENNA__12307__A1 mem_rdata_q\[31\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13065_ _03745_ _04272_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__or2_1
XFILLER_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10277_ _04978_ _04982_ _04928_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12016_ net3020 _06473_ net269 VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__mux2_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08928__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13967_ clknet_leaf_45_clk _00421_ VGND VGND VPWR VPWR cpuregs\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10759__A net800 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11354__S net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12918_ net314 net2437 net457 VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__mux2_1
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13898_ clknet_leaf_51_clk _00352_ VGND VGND VPWR VPWR cpuregs\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09239__A1 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15637_ clknet_leaf_199_clk _01973_ VGND VGND VPWR VPWR cpuregs\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12849_ net328 net2147 net459 VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__mux2_1
XFILLER_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12243__B1 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15568_ clknet_leaf_193_clk _01904_ VGND VGND VPWR VPWR cpuregs\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14519_ clknet_leaf_65_clk _00908_ VGND VGND VPWR VPWR decoded_imm_j\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15499_ clknet_leaf_133_clk _01835_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dfxtp_2
X_08040_ _03360_ _03364_ _03543_ _03545_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__o31a_1
XANTENNA__07670__B1 net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11349__A2 net639 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold903 cpuregs\[18\]\[26\] VGND VGND VPWR VPWR net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 cpuregs\[17\]\[17\] VGND VGND VPWR VPWR net2228 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12913__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08214__A2 net1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold925 cpuregs\[11\]\[12\] VGND VGND VPWR VPWR net2239 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10557__B1 net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 cpuregs\[21\]\[0\] VGND VGND VPWR VPWR net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 cpuregs\[3\]\[7\] VGND VGND VPWR VPWR net2261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__X net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold958 cpuregs\[17\]\[25\] VGND VGND VPWR VPWR net2272 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net1129 _04452_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold969 cpuregs\[5\]\[3\] VGND VGND VPWR VPWR net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11529__S net742 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08942_ genblk1.genblk1.pcpi_mul.rd\[9\] genblk1.genblk1.pcpi_mul.rd\[41\] net954
+ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__mux2_1
XFILLER_69_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08873_ genblk1.genblk1.pcpi_mul.next_rs2\[61\] net1106 _04204_ _04206_ VGND VGND
+ VPWR VPWR _04207_ sky130_fd_sc_hd__a22o_1
Xhold1603 genblk1.genblk1.pcpi_mul.rd\[59\] VGND VGND VPWR VPWR net2917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1614 genblk1.genblk1.pcpi_mul.next_rs2\[49\] VGND VGND VPWR VPWR net2928 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1625 genblk1.genblk1.pcpi_mul.next_rs2\[33\] VGND VGND VPWR VPWR net2939 sky130_fd_sc_hd__dlygate4sd3_1
X_07824_ net1161 net1018 VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__nor2_1
Xhold1636 genblk1.genblk1.pcpi_mul.next_rs2\[4\] VGND VGND VPWR VPWR net2950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1647 genblk2.pcpi_div.quotient\[12\] VGND VGND VPWR VPWR net2961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1658 count_cycle\[21\] VGND VGND VPWR VPWR net2972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1669 genblk1.genblk1.pcpi_mul.next_rs2\[7\] VGND VGND VPWR VPWR net2983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07755_ net1176 net1044 VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout361_A net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A _02118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07686_ cpuregs\[9\]\[3\] net623 net606 _03205_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__o211a_1
XFILLER_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09425_ net3053 _04313_ net1225 VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09356_ net1356 net303 net478 VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__mux2_1
XANTENNA__06882__A net1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08307_ net992 _03737_ net982 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__mux2_1
XFILLER_21_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09287_ net1970 _03844_ net487 VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__mux2_1
XFILLER_139_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout414_X net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10608__S net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_X net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08238_ net1172 net248 net940 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__mux2_1
XFILLER_166_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08169_ _03271_ _03294_ _03648_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__and3_1
XANTENNA__12823__S net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10200_ decoded_imm\[23\] net1006 VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__and2_1
X_11180_ net1158 net856 _05856_ _05857_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout783_X net783 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10131_ count_cycle\[48\] count_cycle\[49\] VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__and2_1
XANTENNA__11666__C _06223_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10062_ count_cycle\[23\] count_cycle\[24\] _04804_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__and3_1
XANTENNA__07218__A net1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14870_ clknet_leaf_7_clk _01222_ VGND VGND VPWR VPWR cpuregs\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13821_ clknet_leaf_198_clk _00275_ VGND VGND VPWR VPWR cpuregs\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13752_ clknet_leaf_193_clk _00206_ VGND VGND VPWR VPWR cpuregs\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10964_ net825 _05642_ _05646_ net779 VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__a211o_1
XFILLER_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10298__B net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12703_ net1191 genblk1.genblk1.pcpi_mul.next_rs1\[0\] net2409 net897 _02085_ VGND
+ VGND VPWR VPWR _01371_ sky130_fd_sc_hd__a221o_1
XFILLER_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13683_ clknet_leaf_117_clk _00137_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_10895_ cpuregs\[11\]\[15\] net618 net589 _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_80_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15422_ clknet_leaf_57_clk _01761_ VGND VGND VPWR VPWR cpuregs\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11028__A1 net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12634_ net2814 net890 _02066_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__a21o_1
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11579__A2 net740 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14782__Q genblk2.pcpi_div.pcpi_rd\[29\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15353_ clknet_leaf_55_clk _01693_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfxtp_1
X_12565_ _02398_ _02045_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09641__B2 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14304_ clknet_leaf_110_clk _00758_ VGND VGND VPWR VPWR count_cycle\[49\] sky130_fd_sc_hd__dfxtp_1
X_11516_ mem_rdata_q\[9\] net1863 net738 VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__mux2_1
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15284_ clknet_leaf_2_clk _01625_ VGND VGND VPWR VPWR cpuregs\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12496_ _01991_ _01992_ net2536 net387 VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_156_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12523__B1_N net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14235_ clknet_leaf_177_clk _00689_ VGND VGND VPWR VPWR reg_next_pc\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_150_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11447_ cpuregs\[14\]\[30\] cpuregs\[15\]\[30\] net689 VGND VGND VPWR VPWR _06117_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output88_A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11378_ cpuregs\[11\]\[28\] net637 net598 _06049_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__o211a_1
XFILLER_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14166_ clknet_leaf_126_clk _00620_ VGND VGND VPWR VPWR count_instr\[37\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10761__B net666 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07955__A1 net771 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10329_ net1188 decoded_imm\[31\] VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__or2_1
XFILLER_3_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13117_ net329 net2464 net435 VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ clknet_leaf_179_clk _00551_ VGND VGND VPWR VPWR cpuregs\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_13048_ net1681 net71 net534 VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__mux2_1
XANTENNA__13564__S net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11592__B mem_rdata_q\[28\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14999_ clknet_leaf_150_clk _01351_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07540_ _02702_ _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_12_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10475__C1 net839 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07471_ count_cycle\[21\] net973 net844 _03002_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__o211a_1
XANTENNA__12908__S net455 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09880__A1 net851 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09210_ net1453 net347 net492 VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__mux2_1
XANTENNA__11019__A1 net822 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08246__X net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09141_ net1564 net406 net501 VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__mux2_1
XANTENNA__11424__D1 net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09072_ net1728 net354 net509 VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__mux2_1
XANTENNA__07643__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08023_ _03529_ _03530_ net1143 VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold700 cpuregs\[2\]\[20\] VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10952__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold711 cpuregs\[10\]\[19\] VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 cpuregs\[3\]\[4\] VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07737__S net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold733 cpuregs\[21\]\[2\] VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 cpuregs\[6\]\[24\] VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 cpuregs\[6\]\[21\] VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_153_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold766 cpuregs\[14\]\[11\] VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 genblk1.genblk1.pcpi_mul.pcpi_rd\[17\] VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold788 cpuregs\[7\]\[8\] VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09974_ _04450_ _04736_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__nor2_1
Xhold799 cpuregs\[15\]\[1\] VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10950__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08925_ net1393 _04239_ net945 VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__mux2_1
Xhold1400 _06590_ VGND VGND VPWR VPWR net2714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout576_A _03756_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13474__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1411 genblk2.pcpi_div.quotient\[24\] VGND VGND VPWR VPWR net2725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _06596_ VGND VGND VPWR VPWR net2736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 count_cycle\[28\] VGND VGND VPWR VPWR net2747 sky130_fd_sc_hd__dlygate4sd3_1
X_08856_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__inv_2
Xhold1444 count_cycle\[56\] VGND VGND VPWR VPWR net2758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07472__S net1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1455 genblk2.pcpi_div.divisor\[18\] VGND VGND VPWR VPWR net2769 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ net250 net1006 VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__nand2_1
Xhold1466 genblk1.genblk1.pcpi_mul.rdx\[32\] VGND VGND VPWR VPWR net2780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1477 genblk2.pcpi_div.quotient_msk\[25\] VGND VGND VPWR VPWR net2791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1488 instr_slti VGND VGND VPWR VPWR net2802 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout364_X net364 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08787_ genblk1.genblk1.pcpi_mul.next_rs2\[48\] net1095 genblk1.genblk1.pcpi_mul.rd\[47\]
+ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__a21o_1
XANTENNA__10399__A net1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1499 _06598_ VGND VGND VPWR VPWR net2813 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_40_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07738_ _03255_ _03256_ net807 VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__mux2_1
XFILLER_169_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10466__C1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout910_A _03879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_X net531 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12818__S net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07669_ net1080 _03189_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout629_X net629 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09408_ cpu_state\[1\] count_instr\[1\] count_instr\[0\] net1186 VGND VGND VPWR VPWR
+ _04303_ sky130_fd_sc_hd__and4_1
XFILLER_158_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10680_ cpuregs\[28\]\[9\] cpuregs\[29\]\[9\] net670 VGND VGND VPWR VPWR _05371_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12758__B2 net995 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09339_ net1805 net522 net475 VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__mux2_1
XANTENNA__13222__B net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10769__B1 net860 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09623__B2 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07634__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12350_ net1151 decoded_imm_j\[1\] _06223_ mem_rdata_q\[21\] net734 VGND VGND VPWR
+ VPWR _06657_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout998_X net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11301_ net820 _05974_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__or2_1
XFILLER_153_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12281_ _06223_ _06617_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__or2_1
XANTENNA__12553__S net874 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13183__A1 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14020_ clknet_leaf_43_clk _00474_ VGND VGND VPWR VPWR cpuregs\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11232_ net835 _05903_ _05905_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__a211o_1
XANTENNA__11194__B1 net595 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11733__A2 _06242_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12930__A1 net1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11163_ _05839_ _05840_ net816 VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__mux2_1
XFILLER_122_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10941__B1 net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10114_ count_cycle\[41\] count_cycle\[42\] count_cycle\[43\] _04836_ VGND VGND VPWR
+ VPWR _04841_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_73_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _05771_ _05773_ net782 VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__a21o_1
X_10045_ count_cycle\[18\] _04791_ _04795_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__and3_1
X_14922_ clknet_leaf_108_clk _01274_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06787__A net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold60 genblk1.genblk1.pcpi_mul.pcpi_rd\[9\] VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 cpuregs\[22\]\[20\] VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 cpuregs\[12\]\[29\] VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14777__Q genblk2.pcpi_div.pcpi_rd\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14853_ clknet_leaf_54_clk _01205_ VGND VGND VPWR VPWR cpuregs\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold93 cpuregs\[14\]\[28\] VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output126_A net1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ clknet_leaf_52_clk _00258_ VGND VGND VPWR VPWR cpuregs\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11249__A1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14784_ clknet_leaf_149_clk _00040_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_11996_ net867 _06456_ net271 VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__o21ai_1
XFILLER_16_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12997__A1 net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13735_ clknet_leaf_113_clk _00189_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10947_ cpuregs\[24\]\[16\] net656 VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__or2_1
XANTENNA__13413__A net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13666_ clknet_leaf_118_clk _00120_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_10878_ net1075 decoded_imm\[14\] VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__or2_1
XANTENNA__09102__S net505 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15405_ clknet_leaf_181_clk _01744_ VGND VGND VPWR VPWR cpuregs\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12617_ net1195 genblk1.genblk1.pcpi_mul.next_rs2\[8\] net915 net1169 VGND VGND VPWR
+ VPWR _02058_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_152_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12029__A net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13597_ clknet_leaf_28_clk _00052_ VGND VGND VPWR VPWR cpuregs\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15336_ clknet_leaf_149_clk _01676_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08941__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12548_ net252 _02032_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13559__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12463__S net383 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15267_ clknet_leaf_47_clk _01608_ VGND VGND VPWR VPWR cpuregs\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12479_ genblk2.pcpi_div.divisor\[42\] net870 VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__nor2_1
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14218_ clknet_leaf_68_clk _00672_ VGND VGND VPWR VPWR reg_pc\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_144_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15198_ clknet_leaf_6_clk _01547_ VGND VGND VPWR VPWR cpuregs\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07928__A1 _02397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11185__B1 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14149_ clknet_leaf_97_clk _00603_ VGND VGND VPWR VPWR count_instr\[20\] sky130_fd_sc_hd__dfxtp_1
Xfanout509 _04278_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_2
X_06971_ genblk2.pcpi_div.dividend\[8\] _02548_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08710_ _04067_ _04068_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__nand2_1
XANTENNA__11488__A1 net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11488__B2 net1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08388__S net766 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09690_ _04474_ _04484_ _04485_ net984 VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a31o_1
Xfanout1080 net1081 VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__buf_2
XANTENNA__07156__A2 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1091 net1093 VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__buf_2
X_08641_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__inv_2
XFILLER_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09504__C _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07305__B decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08572_ genblk1.genblk1.pcpi_mul.next_rs2\[15\] net1090 genblk1.genblk1.pcpi_mul.rd\[14\]
+ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__a21o_1
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07523_ net18 net938 net937 VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_25_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13323__A net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07454_ count_instr\[52\] net1134 net978 _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__a211o_1
XANTENNA__10463__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11660__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09012__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07385_ reg_pc\[16\] decoded_imm\[16\] VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__or2_1
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09605__B2 net846 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_A net1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09124_ net2244 net283 net506 VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__mux2_1
XFILLER_109_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10953__Y _05637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13469__S net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09055_ net291 net2413 net514 VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__mux2_1
XFILLER_136_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12373__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout1233_A net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08006_ _03431_ _03515_ net988 VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__mux2_1
Xhold530 cpuregs\[16\]\[1\] VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold541 cpuregs\[15\]\[22\] VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold552 cpuregs\[4\]\[7\] VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _00973_ VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold574 cpuregs\[27\]\[20\] VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1021_X net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold585 cpuregs\[25\]\[11\] VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold596 cpuregs\[5\]\[0\] VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07395__A2 net939 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09957_ net2597 net880 _04731_ net850 VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout481_X net481 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A _05133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net959 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06878__Y _02477_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08908_ _04046_ _04048_ _04045_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11479__A1 net1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08298__S net924 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09888_ _04664_ _04668_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__nand2_1
Xhold1230 genblk1.genblk1.pcpi_mul.next_rs1\[3\] VGND VGND VPWR VPWR net2544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 _00822_ VGND VGND VPWR VPWR net2555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1252 genblk2.pcpi_div.divisor\[39\] VGND VGND VPWR VPWR net2566 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ genblk1.genblk1.pcpi_mul.next_rs2\[56\] net1104 genblk1.genblk1.pcpi_mul.rd\[55\]
+ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__a21o_1
Xhold1263 genblk1.genblk1.pcpi_mul.rd\[28\] VGND VGND VPWR VPWR net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 net195 VGND VGND VPWR VPWR net2588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout746_X net746 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1285 genblk2.pcpi_div.divisor\[40\] VGND VGND VPWR VPWR net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 genblk1.genblk1.pcpi_mul.rd\[52\] VGND VGND VPWR VPWR net2610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12428__B1 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ genblk2.pcpi_div.divisor\[1\] genblk2.pcpi_div.dividend\[1\] VGND VGND VPWR
+ VPWR _06321_ sky130_fd_sc_hd__xnor2_1
X_10801_ net787 _05484_ _05486_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__or4_1
X_11781_ net2817 _06254_ net536 VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout913_X net913 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11100__B1 net605 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13520_ _03742_ _04273_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__or2_4
XANTENNA__13233__A net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11651__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10732_ net1076 decoded_imm\[10\] VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__or2_1
XFILLER_159_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07377__B1_N net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13451_ reg_pc\[30\] _05079_ _06143_ is_lui_auipc_jal VGND VGND VPWR VPWR _02353_
+ sky130_fd_sc_hd__o2bb2a_1
X_10663_ cpuregs\[6\]\[9\] cpuregs\[7\]\[9\] net671 VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13520__X _02357_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12402_ net403 net2043 net471 VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__mux2_1
X_10594_ cpuregs\[3\]\[7\] net630 net595 _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__o211a_1
X_13382_ net558 _02270_ _02289_ _02291_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__a31o_1
XFILLER_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15121_ clknet_leaf_182_clk _01473_ VGND VGND VPWR VPWR cpuregs\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12333_ decoded_imm\[8\] net735 _06643_ mem_rdata_q\[28\] _06646_ VGND VGND VPWR
+ VPWR _01166_ sky130_fd_sc_hd__a221o_1
XFILLER_127_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15052_ clknet_leaf_102_clk net2502 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12264_ net2743 net381 net369 net2903 VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__a22o_1
XANTENNA__11167__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14003_ clknet_leaf_25_clk _00457_ VGND VGND VPWR VPWR cpuregs\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08032__B1 net770 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11215_ net1082 decoded_imm\[23\] _05133_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__o21a_1
X_12195_ genblk2.pcpi_div.quotient_msk\[11\] net272 net2713 VGND VGND VPWR VPWR _06590_
+ sky130_fd_sc_hd__a21oi_1
Xoutput50 net50 VGND VGND VPWR VPWR mem_addr[25] sky130_fd_sc_hd__buf_2
Xoutput61 net61 VGND VGND VPWR VPWR mem_addr[6] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VGND VGND VPWR VPWR mem_la_addr[16] sky130_fd_sc_hd__buf_2
Xoutput83 net83 VGND VGND VPWR VPWR mem_la_addr[27] sky130_fd_sc_hd__buf_2
X_11146_ cpuregs\[4\]\[22\] cpuregs\[5\]\[22\] net686 VGND VGND VPWR VPWR _05824_
+ sky130_fd_sc_hd__mux2_1
Xoutput94 net94 VGND VGND VPWR VPWR mem_la_addr[8] sky130_fd_sc_hd__buf_2
XANTENNA_output243_A net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__06788__Y _02396_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13408__A net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11077_ cpuregs\[27\]\[20\] net622 net591 _05756_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__o211a_1
XFILLER_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07138__A2 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10678__C1 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14905_ clknet_leaf_142_clk _01257_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_10028_ count_cycle\[10\] count_cycle\[11\] count_cycle\[12\] _04781_ VGND VGND VPWR
+ VPWR _04786_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_196_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_196_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_37_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14836_ clknet_leaf_195_clk _01188_ VGND VGND VPWR VPWR cpuregs\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10693__A2 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08936__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11494__C_N net267 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08099__B1 net967 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14767_ clknet_leaf_163_clk _00021_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11979_ net865 _06439_ _06441_ _06442_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__a22o_1
X_13718_ clknet_leaf_138_clk _00172_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11642__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14698_ clknet_leaf_152_clk _01083_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07141__A _02383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13649_ clknet_leaf_118_clk _00103_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07170_ net1139 count_cycle\[34\] net976 _02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a211o_1
XFILLER_157_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15319_ clknet_leaf_7_clk _01659_ VGND VGND VPWR VPWR cpuregs\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08271__A0 net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11945__A2 _02443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07795__B net994 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10706__S net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_117_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11158__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12921__S net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout306 net307 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09811_ _04592_ _04597_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout317 net318 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_2
Xfanout328 _03818_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 _03807_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkload11_A clknet_4_11_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09742_ decoded_imm_j\[10\] _04431_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__nand2_1
XANTENNA__12222__A net749 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06954_ _02532_ _02534_ net949 VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__mux2_1
XFILLER_67_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09007__S net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09523__B1 net1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09673_ _02481_ _04469_ _04471_ _02489_ _04470_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__o221a_1
X_06885_ net961 _02483_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_187_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_187_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_143_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout274_A net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08624_ genblk1.genblk1.pcpi_mul.next_rs2\[23\] net1104 genblk1.genblk1.pcpi_mul.rd\[22\]
+ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_6_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13083__A0 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08555_ _03931_ _03934_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__nand2_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout441_A net442 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10677__A net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12368__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07506_ reg_pc\[24\] decoded_imm\[24\] VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08486_ genblk1.genblk1.pcpi_mul.next_rs2\[1\] net1102 genblk1.genblk1.pcpi_mul.rd\[0\]
+ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a21o_1
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10396__B net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07437_ count_cycle\[19\] net973 net843 _02970_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout706_A net707 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_X net1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12189__A2 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13386__A1 net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07368_ reg_pc\[15\] decoded_imm\[15\] VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__nand2_1
XANTENNA__08434__X _03839_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09107_ net1887 net347 net504 VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__mux2_1
XANTENNA__10616__S net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07299_ net1139 count_cycle\[42\] net976 _02841_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_111_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_92_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11301__A net820 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09038_ net356 net2312 net512 VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout696_X net696 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold360 cpuregs\[29\]\[30\] VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12831__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold371 cpuregs\[8\]\[8\] VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold382 cpuregs\[27\]\[2\] VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 cpuregs\[15\]\[14\] VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ cpuregs\[1\]\[18\] net549 _05681_ net796 net823 VGND VGND VPWR VPWR _05682_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_53_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09762__B1 _02380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10372__A1 net992 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout840 _03136_ VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__buf_2
Xfanout851 net852 VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__clkbuf_4
Xfanout862 net865 VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__clkbuf_4
Xfanout873 net874 VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__clkbuf_2
Xfanout884 net898 VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13310__B2 net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout895 net896 VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__buf_2
X_12951_ net338 net2155 net452 VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__mux2_1
XANTENNA__15216__Q cpu_state\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_178_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_178_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11321__B1 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1060 cpuregs\[17\]\[21\] VGND VGND VPWR VPWR net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 cpuregs\[2\]\[14\] VGND VGND VPWR VPWR net2385 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ genblk2.pcpi_div.divisor\[26\] genblk2.pcpi_div.dividend\[26\] VGND VGND
+ VPWR VPWR _06373_ sky130_fd_sc_hd__nand2b_1
Xhold1082 cpuregs\[17\]\[7\] VGND VGND VPWR VPWR net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12882_ mem_rdata_q\[19\] net11 net962 VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__mux2_1
Xhold1093 cpuregs\[17\]\[22\] VGND VGND VPWR VPWR net2407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07660__S net701 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14621_ clknet_leaf_109_clk _01007_ VGND VGND VPWR VPWR genblk2.pcpi_div.instr_div
+ sky130_fd_sc_hd__dfxtp_1
X_11833_ genblk2.pcpi_div.divisor\[10\] genblk2.pcpi_div.dividend\[10\] VGND VGND
+ VPWR VPWR _06304_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14552_ clknet_leaf_184_clk _00938_ VGND VGND VPWR VPWR cpuregs\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11764_ net1673 net118 net729 VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13503_ net1776 net341 net419 VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__mux2_1
X_10715_ cpuregs\[28\]\[10\] cpuregs\[29\]\[10\] net669 VGND VGND VPWR VPWR _05405_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ clknet_leaf_94_clk _00872_ VGND VGND VPWR VPWR instr_slti sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ net2033 net355 net373 VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__mux2_1
X_13434_ net998 net756 _02133_ _02315_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__o211a_1
X_10646_ cpuregs\[24\]\[8\] net670 VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__or2_1
XFILLER_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output193_A net193 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08253__A0 net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_8
X_13365_ net1004 net760 VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__or2_1
XFILLER_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10577_ _05269_ _05270_ net814 VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__mux2_1
XANTENNA__11211__A net788 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15104_ clknet_leaf_36_clk _01456_ VGND VGND VPWR VPWR cpuregs\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12316_ net1146 decoded_imm_j\[15\] net970 mem_rdata_q\[15\] VGND VGND VPWR VPWR
+ _06637_ sky130_fd_sc_hd__a22o_1
X_13296_ net567 _05491_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__nor2_1
XFILLER_170_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15035_ clknet_leaf_135_clk _01387_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12888__A0 mem_rdata_q\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12247_ net2742 net379 net366 net2853 VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output70_A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12178_ net751 _06581_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__nor2_1
XFILLER_122_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11129_ cpuregs\[26\]\[21\] net681 VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13301__B2 net1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_169_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_169_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_160_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13572__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14819_ clknet_leaf_82_clk _01171_ VGND VGND VPWR VPWR decoded_imm\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08340_ reg_pc\[5\] _03758_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__nor2_1
X_08271_ net1026 _03719_ net980 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__mux2_1
XFILLER_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12916__S net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07222_ count_cycle\[5\] net971 net841 _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__o211a_1
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07153_ net1073 decoded_imm\[0\] _02698_ _02705_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__a211o_1
XANTENNA__12040__A1 net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10051__B1 net1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07084_ _02645_ _02646_ _02643_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__o21ai_1
XFILLER_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12879__A0 mem_rdata_q\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1029_A net1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__C1 net823 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout391_A net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_A _04287_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07986_ _03493_ _03498_ VGND VGND VPWR VPWR alu_out\[5\] sky130_fd_sc_hd__nand2_1
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09725_ net1149 _04515_ _04518_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__a21o_1
X_06937_ genblk2.pcpi_div.dividend\[2\] genblk2.pcpi_div.dividend\[1\] genblk2.pcpi_div.dividend\[0\]
+ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout277_X net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A net663 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13482__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10657__A2 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09656_ decoded_imm_j\[2\] _04423_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__and2_1
XANTENNA__06885__A net961 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06868_ instr_lbu instr_lb net410 VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _03975_ _03978_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nand2_1
X_09587_ net1940 _04418_ net1238 VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout823_A net826 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06799_ net1018 VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout444_X net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_X net1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08538_ net887 _03921_ _03923_ net2592 net1193 VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__a32o_1
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10200__A decoded_imm\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08469_ reg_pc\[30\] _03863_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout611_X net611 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08483__B1 net916 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12826__S net466 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13359__A1 net557 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_X net709 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10500_ cpuregs\[17\]\[1\] net636 net612 _05198_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__o211a_1
X_11480_ _02436_ _02438_ net1084 VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__o21a_1
XFILLER_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09200__S net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08235__A0 net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10431_ mem_do_wdata _02702_ _05124_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__and3b_1
XANTENNA__12031__A1 net1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13230__B net568 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13150_ net1664 net334 net431 VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__mux2_1
X_10362_ cpuregs\[28\]\[31\] cpuregs\[29\]\[31\] net694 VGND VGND VPWR VPWR _05068_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout980_X net980 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12101_ _06369_ _06380_ _06377_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__a21o_1
X_13081_ net341 net1628 net439 VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__mux2_1
X_10293_ decoded_imm\[19\] net1012 VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__nor2_1
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12032_ _06485_ _06486_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__nor2_1
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold190 genblk1.genblk1.pcpi_mul.pcpi_rd\[29\] VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout670 net671 VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 net696 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12098__A1 net1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout692 net695 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__clkbuf_4
X_13983_ clknet_leaf_0_clk _00437_ VGND VGND VPWR VPWR cpuregs\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12934_ _03744_ _04283_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06795__A net1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15653_ clknet_leaf_49_clk _01989_ VGND VGND VPWR VPWR cpuregs\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_103_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ net23 mem_rdata_q\[2\] _02450_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__mux2_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output206_A net1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14604_ clknet_leaf_118_clk _00990_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfxtp_1
X_11816_ genblk2.pcpi_div.dividend\[17\] genblk2.pcpi_div.divisor\[17\] VGND VGND
+ VPWR VPWR _06287_ sky130_fd_sc_hd__and2b_1
XANTENNA__07403__B decoded_imm\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15584_ clknet_leaf_57_clk _01920_ VGND VGND VPWR VPWR cpuregs\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_83_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _02414_ _02115_ _02116_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__o21a_1
XFILLER_61_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14535_ clknet_leaf_88_clk _00923_ VGND VGND VPWR VPWR is_lb_lh_lw_lbu_lhu sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ net1965 net100 net730 VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__mux2_1
XANTENNA__11640__S net546 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14466_ clknet_leaf_89_clk _00855_ VGND VGND VPWR VPWR instr_auipc sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_78_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11678_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__inv_2
XANTENNA__09110__S net504 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13417_ net558 _02299_ _02322_ net566 reg_pc\[26\] VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__a32o_1
XANTENNA__08226__B1 net1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10629_ _05319_ _05320_ net815 VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__mux2_1
X_14397_ clknet_leaf_102_clk _00818_ VGND VGND VPWR VPWR pcpi_timeout_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13348_ net1007 net759 VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__or2_1
XANTENNA__11781__B1 net536 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13567__S net411 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13279_ net959 _04976_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__and3_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15018_ clknet_leaf_121_clk _01370_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rs1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12325__A2 mem_rdata_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11533__A0 mem_rdata_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07840_ net1166 net1029 VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_87_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07771_ net254 net998 VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__06960__B1 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09510_ net2992 _04369_ net1226 VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11297__C1 net836 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08396__S net1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09441_ _04325_ net1226 _04324_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__and3b_1
XANTENNA__09512__C _04363_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09372_ net1928 net522 net400 VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__mux2_1
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08323_ reg_out\[1\] alu_out_q\[1\] net1154 VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__mux2_1
XANTENNA__07268__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11064__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07268__B2 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13331__A net1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08254_ reg_out\[4\] reg_next_pc\[4\] net923 VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__mux2_1
XFILLER_166_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09020__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07205_ net27 net130 _02695_ net13 _02753_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__a221o_1
XANTENNA__08217__B1 net265 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12013__A1 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08185_ _03291_ _03297_ _03663_ _03674_ _03290_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__a32oi_2
XANTENNA_fanout404_A _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10393__C net1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09965__B1 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07136_ net1054 net1057 VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__nand2b_2
XFILLER_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13477__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07067_ net1117 _02631_ genblk2.pcpi_div.dividend\[21\] VGND VGND VPWR VPWR _02632_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07440__A1 net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12381__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput240 net240 VGND VGND VPWR VPWR pcpi_rs2[14] sky130_fd_sc_hd__buf_2
Xoutput251 net251 VGND VGND VPWR VPWR pcpi_rs2[24] sky130_fd_sc_hd__buf_2
XFILLER_160_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput262 net262 VGND VGND VPWR VPWR pcpi_rs2[5] sky130_fd_sc_hd__buf_2
XFILLER_88_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12316__A2 decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11524__A0 mem_rdata_q\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _03170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13277__B1 net395 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07969_ _03275_ _03482_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout940_A _02693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09262__Y _04288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09708_ decoded_imm_j\[7\] _04428_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__or2_1
X_10980_ cpuregs\[19\]\[17\] net617 net589 VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__o21a_1
XFILLER_56_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09639_ reg_pc\[25\] net879 _04446_ net849 VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_X net826 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12650_ net1210 net2971 net899 net3002 _02074_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__a221o_1
X_11601_ net1234 is_alu_reg_reg _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__and3_2
XANTENNA__07259__A1 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11055__A2 net632 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12581_ net521 net1911 net467 VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__mux2_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13241__A net1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14320_ clknet_leaf_128_clk _06716_ VGND VGND VPWR VPWR reg_out\[0\] sky130_fd_sc_hd__dfxtp_1
X_11532_ mem_rdata_q\[25\] net2680 net736 VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__mux2_1
XFILLER_168_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14251_ clknet_leaf_68_clk _00705_ VGND VGND VPWR VPWR reg_next_pc\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08208__B1 net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11463_ net832 _06128_ _06130_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__a211o_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ net1042 net709 net557 net1047 VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__a22o_1
XANTENNA__10015__B1 net1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10414_ net258 _05118_ _02507_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11212__C1 net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14182_ clknet_leaf_109_clk net2591 VGND VGND VPWR VPWR count_instr\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11394_ cpuregs\[19\]\[28\] net636 net598 VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__o21a_1
XANTENNA__10566__A1 net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13133_ net1535 net588 net433 VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__mux2_1
X_10345_ net806 _05050_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__or2_1
XANTENNA__07893__B net1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13064_ net2258 net88 net534 VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__mux2_1
XANTENNA__11515__A0 mem_rdata_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10276_ _04935_ _04936_ _04973_ _04980_ _04934_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__a311o_1
XANTENNA__08070__A net968 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12015_ net867 _06468_ _06469_ _06472_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__o31ai_1
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07734__A2 net631 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06796__Y _02404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13416__A net1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ clknet_leaf_36_clk _00420_ VGND VGND VPWR VPWR cpuregs\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08069__X alu_out\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09105__S net505 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12917_ net317 net2336 net457 VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__mux2_1
XANTENNA__07498__A1 genblk2.pcpi_div.pcpi_rd\[23\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13897_ clknet_leaf_56_clk _00351_ VGND VGND VPWR VPWR cpuregs\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12848_ net333 net2522 net459 VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__mux2_1
X_15636_ clknet_leaf_191_clk _01972_ VGND VGND VPWR VPWR cpuregs\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08944__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15567_ clknet_leaf_182_clk _01903_ VGND VGND VPWR VPWR cpuregs\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12466__S net868 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12779_ net1221 net2233 net2489 net909 net765 VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__a221o_1
XFILLER_9_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ clknet_leaf_28_clk _00907_ VGND VGND VPWR VPWR decoded_imm_j\[19\] sky130_fd_sc_hd__dfxtp_1
X_15498_ clknet_leaf_132_clk _01834_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dfxtp_2
XFILLER_147_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14449_ clknet_leaf_55_clk _00838_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold904 cpuregs\[4\]\[18\] VGND VGND VPWR VPWR net2218 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold915 cpuregs\[1\]\[16\] VGND VGND VPWR VPWR net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold926 cpuregs\[19\]\[9\] VGND VGND VPWR VPWR net2240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold937 cpuregs\[17\]\[26\] VGND VGND VPWR VPWR net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 cpuregs\[25\]\[1\] VGND VGND VPWR VPWR net2262 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _04751_ _04753_ _04752_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__a21bo_1
Xhold959 cpuregs\[9\]\[28\] VGND VGND VPWR VPWR net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08941_ net1831 _04247_ net943 VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__mux2_1
XFILLER_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08872_ genblk1.genblk1.pcpi_mul.rd\[60\] genblk1.genblk1.pcpi_mul.rdx\[60\] VGND
+ VGND VPWR VPWR _04206_ sky130_fd_sc_hd__or2_1
XFILLER_111_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1604 genblk1.genblk1.pcpi_mul.rd\[33\] VGND VGND VPWR VPWR net2918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09363__X _04293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1615 _01355_ VGND VGND VPWR VPWR net2929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07725__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1626 count_cycle\[34\] VGND VGND VPWR VPWR net2940 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09804__A decoded_imm_j\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07823_ _02395_ _02407_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__nor2_1
Xhold1637 _01310_ VGND VGND VPWR VPWR net2951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1648 _06591_ VGND VGND VPWR VPWR net2962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06933__B1 net953 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1659 count_instr\[7\] VGND VGND VPWR VPWR net2973 sky130_fd_sc_hd__dlygate4sd3_1
X_07754_ _03269_ _03270_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__nand2_1
XANTENNA__12230__A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09015__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07685_ cpuregs\[8\]\[3\] net662 VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_91_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1096_A net1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09424_ count_instr\[6\] _04313_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__and2_1
XFILLER_53_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09355_ net1358 net307 net477 VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__mux2_1
XANTENNA__12376__S net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A net522 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11280__S net706 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06882__B net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_A net620 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08306_ reg_out\[30\] reg_next_pc\[30\] net924 VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09286_ net1612 net308 net486 VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__mux2_1
XANTENNA__10796__A1 net812 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08237_ net1175 net247 net940 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__mux2_1
XFILLER_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout1051_X net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1149_X net1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08168_ net966 _03296_ _03297_ net929 _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout988_A net990 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07119_ genblk2.pcpi_div.dividend\[29\] net1123 _02669_ net948 VGND VGND VPWR VPWR
+ _02676_ sky130_fd_sc_hd__a31o_1
XANTENNA__07413__A1 genblk2.pcpi_div.pcpi_rd\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08099_ net1159 net1012 net967 VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__o21a_1
XFILLER_122_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10130_ count_cycle\[47\] count_cycle\[48\] _04846_ count_cycle\[49\] VGND VGND VPWR
+ VPWR _04851_ sky130_fd_sc_hd__a31o_1
XANTENNA__07964__A2 net930 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout776_X net776 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10061_ _04806_ _04807_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__nor2_1
XANTENNA__07218__B net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout943_X net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_197_clk _00274_ VGND VGND VPWR VPWR cpuregs\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12140__A net1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13751_ clknet_leaf_181_clk _00205_ VGND VGND VPWR VPWR cpuregs\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10963_ cpuregs\[3\]\[17\] net623 net592 _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__o211a_1
XANTENNA__11276__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12702_ _02383_ net912 VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13682_ clknet_leaf_117_clk _00136_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10894_ cpuregs\[10\]\[15\] net647 VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15421_ clknet_leaf_57_clk _01760_ VGND VGND VPWR VPWR cpuregs\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__08991__C _03743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ net1198 genblk1.genblk1.pcpi_mul.next_rs2\[16\] net915 net1162 VGND VGND
+ VPWR VPWR _02066_ sky130_fd_sc_hd__a22o_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15352_ clknet_leaf_62_clk _01692_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12564_ net255 _05117_ net719 VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__o21a_1
XANTENNA__09641__A2 net879 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14303_ clknet_leaf_110_clk _00757_ VGND VGND VPWR VPWR count_cycle\[48\] sky130_fd_sc_hd__dfxtp_1
X_11515_ mem_rdata_q\[8\] net1924 net736 VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__mux2_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15283_ clknet_leaf_2_clk _01624_ VGND VGND VPWR VPWR cpuregs\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12495_ net871 _06715_ _01990_ net387 VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__a31o_1
XFILLER_138_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14234_ clknet_leaf_177_clk _00688_ VGND VGND VPWR VPWR reg_next_pc\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11446_ cpuregs\[12\]\[30\] cpuregs\[13\]\[30\] net689 VGND VGND VPWR VPWR _06116_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14165_ clknet_leaf_126_clk _00619_ VGND VGND VPWR VPWR count_instr\[36\] sky130_fd_sc_hd__dfxtp_1
X_11377_ cpuregs\[10\]\[28\] net689 VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__or2_1
XFILLER_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13116_ net334 net2354 net435 VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__mux2_1
X_10328_ _04893_ _04894_ _05032_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__nor3_1
XANTENNA__07409__A net358 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14096_ clknet_leaf_32_clk _00550_ VGND VGND VPWR VPWR cpuregs\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13047_ net1363 net70 net535 VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__mux2_1
X_10259_ _04937_ _04939_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__nor2_1
XFILLER_39_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08939__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07168__B1 _02695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1240 net1241 VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__buf_1
XFILLER_94_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11365__S net692 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12050__A net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14998_ clknet_leaf_149_clk net2827 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_13949_ clknet_leaf_198_clk _00403_ VGND VGND VPWR VPWR cpuregs\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13580__S net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07470_ count_instr\[21\] net1138 net978 _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__a211o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15619_ clknet_4_11_0_clk _01955_ VGND VGND VPWR VPWR cpuregs\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_09140_ net1867 net409 net500 VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10778__A1 net826 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09071_ net1534 net405 net509 VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__mux2_1
XANTENNA__12924__S net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08022_ _03356_ _03431_ _03414_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__o21bai_1
Xhold701 cpuregs\[4\]\[9\] VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__D1 net792 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold712 cpuregs\[6\]\[9\] VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 cpuregs\[2\]\[15\] VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 cpuregs\[13\]\[31\] VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 cpuregs\[13\]\[0\] VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold756 cpuregs\[16\]\[13\] VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 cpuregs\[8\]\[9\] VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold778 cpuregs\[25\]\[6\] VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _04741_ _04744_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__a21o_1
Xhold789 cpuregs\[20\]\[19\] VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_168_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07876__A_N net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ genblk1.genblk1.pcpi_mul.rd\[0\] genblk1.genblk1.pcpi_mul.rd\[32\] net956
+ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__mux2_1
XFILLER_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1401 genblk2.pcpi_div.divisor\[7\] VGND VGND VPWR VPWR net2715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 _06603_ VGND VGND VPWR VPWR net2726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08855_ _04183_ _04186_ _04188_ _04190_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__o211a_1
Xhold1423 net199 VGND VGND VPWR VPWR net2737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout471_A net472 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1434 genblk1.genblk1.pcpi_mul.rd\[21\] VGND VGND VPWR VPWR net2748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout569_A net570 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1445 genblk1.genblk1.pcpi_mul.next_rs2\[1\] VGND VGND VPWR VPWR net2759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 _01123_ VGND VGND VPWR VPWR net2770 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07806_ _03320_ _03322_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_146_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08786_ genblk1.genblk1.pcpi_mul.rd\[47\] genblk1.genblk1.pcpi_mul.next_rs2\[48\]
+ net1094 VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__nand3_1
Xhold1467 genblk1.genblk1.pcpi_mul.rd\[25\] VGND VGND VPWR VPWR net2781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1478 _01066_ VGND VGND VPWR VPWR net2792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10399__B net1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1489 genblk2.pcpi_div.quotient_msk\[12\] VGND VGND VPWR VPWR net2803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07737_ cpuregs\[22\]\[4\] cpuregs\[23\]\[4\] net701 VGND VGND VPWR VPWR _03256_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11258__A2 net642 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout736_A net738 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout357_X net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13490__S net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06893__A instr_jal VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07668_ net775 _03180_ _03188_ _03172_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__a31o_1
XFILLER_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09407_ _04302_ net1231 _04301_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__and3b_1
XANTENNA__13404__B1 net958 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07599_ count_cycle\[30\] net974 net843 _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout903_A _03879_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_X net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09338_ net1847 net525 net475 VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__mux2_1
XFILLER_138_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09623__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11023__B net647 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09269_ net1643 net539 net484 VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__mux2_1
XANTENNA__12834__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11430__A2 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11300_ cpuregs\[14\]\[26\] cpuregs\[15\]\[26\] net704 VGND VGND VPWR VPWR _05974_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12280_ is_beq_bne_blt_bge_bltu_bgeu is_sb_sh_sw VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__or2_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11231_ cpuregs\[18\]\[24\] net555 _05906_ net786 VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__o22a_1
XANTENNA__11677__C net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07937__A2 _03389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11162_ cpuregs\[28\]\[22\] cpuregs\[29\]\[22\] net683 VGND VGND VPWR VPWR _05840_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09139__A1 net523 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10113_ _04840_ net1225 _04839_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__and3b_1
XFILLER_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ cpuregs\[1\]\[20\] net549 _05772_ net799 net825 VGND VGND VPWR VPWR _05773_
+ sky130_fd_sc_hd__a221o_1
XFILLER_96_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12143__B1 net372 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input32_A mem_rdata[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10044_ _04791_ _04795_ count_cycle\[18\] VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__a21o_1
X_14921_ clknet_leaf_109_clk _01273_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[60\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold50 genblk1.genblk1.pcpi_mul.next_rs1\[6\] VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold61 cpuregs\[12\]\[27\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold72 cpuregs\[20\]\[4\] VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ clknet_leaf_69_clk _01204_ VGND VGND VPWR VPWR cpuregs\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold83 cpuregs\[30\]\[0\] VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 cpuregs\[30\]\[28\] VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13803_ clknet_leaf_72_clk _00257_ VGND VGND VPWR VPWR cpuregs\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14783_ clknet_leaf_149_clk _00039_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[30\]
+ sky130_fd_sc_hd__dfxtp_2
X_11995_ _06304_ _06339_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_55_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_output119_A net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13734_ clknet_leaf_113_clk _00188_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10946_ _05628_ _05629_ net810 VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13665_ clknet_leaf_119_clk _00119_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_10877_ _05536_ _05545_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__a21oi_2
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11214__A net1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11406__C1 net837 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15404_ clknet_leaf_182_clk _01743_ VGND VGND VPWR VPWR cpuregs\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12616_ net2902 net892 _02057_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__a21o_1
XANTENNA__12749__A2 net897 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ clknet_leaf_45_clk _00051_ VGND VGND VPWR VPWR cpuregs\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15335_ clknet_leaf_145_clk _01675_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_1
X_12547_ net251 _05114_ net719 VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11421__A2 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15266_ clknet_leaf_38_clk _01607_ VGND VGND VPWR VPWR cpuregs\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12478_ _05102_ net718 net1166 VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_113_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14217_ clknet_leaf_75_clk _00671_ VGND VGND VPWR VPWR reg_pc\[25\] sky130_fd_sc_hd__dfxtp_1
X_11429_ cpuregs\[17\]\[29\] net644 net615 _06099_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__o211a_1
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15197_ clknet_leaf_18_clk _01546_ VGND VGND VPWR VPWR cpuregs\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07928__A2 net998 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14148_ clknet_leaf_97_clk _00602_ VGND VGND VPWR VPWR count_instr\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13575__S net413 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14079_ clknet_leaf_2_clk _00533_ VGND VGND VPWR VPWR cpuregs\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_06970_ genblk2.pcpi_div.dividend\[7\] _02541_ net1118 VGND VGND VPWR VPWR _02548_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_67_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07426__X _02961_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12685__A1 net1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1070 cpu_state\[5\] VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_163_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1081 net1087 VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08640_ genblk1.genblk1.pcpi_mul.next_rs2\[25\] net1103 _04006_ _04008_ VGND VGND
+ VPWR VPWR _04010_ sky130_fd_sc_hd__and4_1
Xfanout1092 net1093 VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08571_ net885 _03949_ _03951_ net2765 net1192 VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__a32o_1
XANTENNA__12919__S net456 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07522_ _03035_ _03037_ _03048_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__nand3_1
XANTENNA__08257__X net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07453_ count_instr\[20\] net1138 count_cycle\[52\] net1142 VGND VGND VPWR VPWR _02986_
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07384_ _02920_ _02921_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__or2_1
XANTENNA__09605__A2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09123_ net1992 net285 net507 VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__mux2_1
XFILLER_148_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07616__A1 net986 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09054_ net293 net2418 net514 VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__mux2_1
XFILLER_129_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08005_ _03315_ _03508_ _03317_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__a21oi_1
Xhold520 net65 VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 cpuregs\[22\]\[3\] VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11176__A1 net831 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold542 cpuregs\[15\]\[5\] VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold553 cpuregs\[31\]\[9\] VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold564 cpuregs\[16\]\[22\] VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold575 cpuregs\[21\]\[3\] VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 cpuregs\[2\]\[0\] VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13485__S net425 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold597 cpuregs\[5\]\[8\] VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09956_ _04448_ _04730_ net1185 VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__mux2_1
XANTENNA__06888__A net1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_X net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08907_ net1212 net2625 net904 _04230_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__a22o_1
XANTENNA__07336__X _06719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09887_ _04621_ _04665_ _04667_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout474_X net474 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1220 genblk2.pcpi_div.divisor\[53\] VGND VGND VPWR VPWR net2534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 genblk2.pcpi_div.divisor\[35\] VGND VGND VPWR VPWR net2545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 net216 VGND VGND VPWR VPWR net2556 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ genblk1.genblk1.pcpi_mul.rd\[55\] genblk1.genblk1.pcpi_mul.next_rs2\[56\]
+ net1103 VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1253 genblk1.genblk1.pcpi_mul.rd\[16\] VGND VGND VPWR VPWR net2567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 reg_next_pc\[19\] VGND VGND VPWR VPWR net2578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07552__B1 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1275 genblk2.pcpi_div.divisor\[61\] VGND VGND VPWR VPWR net2589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1286 genblk2.pcpi_div.divisor\[50\] VGND VGND VPWR VPWR net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1297 net180 VGND VGND VPWR VPWR net2611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08769_ genblk1.genblk1.pcpi_mul.next_rs2\[45\] net1090 _04116_ _04118_ VGND VGND
+ VPWR VPWR _04119_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout641_X net641 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12829__S net466 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_X net739 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_10800_ cpuregs\[11\]\[12\] net619 net589 _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__o211a_1
XANTENNA__10439__B1 net597 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11780_ _02448_ _06238_ _06252_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__a211o_1
XANTENNA__09203__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10731_ net773 _05412_ _05420_ _05404_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__a31oi_4
XFILLER_15_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13450_ _04879_ _02349_ _02350_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__or4_1
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10662_ net1168 net853 _05352_ _05353_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12401_ net408 net2015 net472 VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__mux2_1
XANTENNA__11403__A2 net644 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13381_ net710 _02271_ _02290_ _04879_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__a31o_1
X_10593_ cpuregs\[2\]\[7\] net673 VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15120_ clknet_leaf_184_clk _01472_ VGND VGND VPWR VPWR cpuregs\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__10611__B1 net593 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12332_ net1148 decoded_imm_j\[8\] net744 VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__and3_1
XFILLER_166_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15051_ clknet_leaf_102_clk _01403_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12263_ genblk2.pcpi_div.divisor\[26\] net381 net369 net2743 VGND VGND VPWR VPWR
+ _01132_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14002_ clknet_leaf_29_clk _00456_ VGND VGND VPWR VPWR cpuregs\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11214_ net1082 _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__nand2_1
X_12194_ net749 _06589_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__nor2_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput40 net40 VGND VGND VPWR VPWR mem_addr[15] sky130_fd_sc_hd__buf_2
Xoutput51 net51 VGND VGND VPWR VPWR mem_addr[26] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VGND VGND VPWR VPWR mem_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_122_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput73 net73 VGND VGND VPWR VPWR mem_la_addr[17] sky130_fd_sc_hd__buf_2
X_11145_ cpuregs\[6\]\[22\] cpuregs\[7\]\[22\] net686 VGND VGND VPWR VPWR _05823_
+ sky130_fd_sc_hd__mux2_1
Xoutput84 net84 VGND VGND VPWR VPWR mem_la_addr[28] sky130_fd_sc_hd__buf_2
XANTENNA__06798__A net1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12116__B1 net997 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput95 net95 VGND VGND VPWR VPWR mem_la_addr[9] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_14_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11076_ cpuregs\[26\]\[20\] net658 VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__or2_1
XANTENNA__13408__B net760 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output236_A net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14904_ clknet_leaf_144_clk _01256_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_10027_ _04785_ net1224 _04784_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__and3b_1
XFILLER_91_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14835_ clknet_leaf_3_clk _01187_ VGND VGND VPWR VPWR cpuregs\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_106_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11643__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08099__A1 net1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14766_ clknet_leaf_163_clk _00020_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_11978_ net1036 _06440_ net868 VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__o21a_1
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09113__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_152_clk_A clknet_4_5_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13717_ clknet_leaf_151_clk _00171_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_10929_ net810 _05610_ _05612_ net824 VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__o211a_1
X_14697_ clknet_leaf_152_clk _01082_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10850__B1 net781 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08952__S net954 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13648_ clknet_leaf_144_clk _00102_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_9_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09599__B2 net847 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13395__A2 net397 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13579_ net301 net2272 net414 VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__mux2_1
XFILLER_157_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_167_clk_A clknet_4_4_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15318_ clknet_leaf_9_clk _01658_ VGND VGND VPWR VPWR cpuregs\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11945__A3 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15249_ clknet_leaf_32_clk _01590_ VGND VGND VPWR VPWR cpuregs\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12355__B1 net956 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09810_ _04571_ _04595_ _04596_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__o21ba_1
Xfanout307 _03844_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout318 net319 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_2
Xfanout329 _03818_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_1
XANTENNA__08399__S net528 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09741_ net845 _04532_ _04533_ net875 net2638 VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__a32o_1
X_06953_ genblk2.pcpi_div.quotient\[5\] _02533_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_15_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09672_ _04423_ _04424_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__nand2_1
X_06884_ mem_do_prefetch _02452_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09812__A _02480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08623_ net900 _03993_ _03995_ net2748 net1202 VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_19_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_08554_ _03935_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__nand2_1
XFILLER_36_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09023__S net518 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07505_ reg_pc\[24\] decoded_imm\[24\] VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__or2_1
XANTENNA__11094__B1 net782 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08485_ genblk1.genblk1.pcpi_mul.mul_waiting net1216 VGND VGND VPWR VPWR _03879_
+ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_18_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1176_A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07436_ count_instr\[19\] net1138 net978 _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__a211o_1
XFILLER_149_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13386__A2 net393 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12384__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07367_ reg_pc\[15\] decoded_imm\[15\] VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout601_A _03153_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11397__A1 net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09106_ net1744 net350 net504 VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__mux2_1
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07298_ count_instr\[42\] net1131 net1135 count_instr\[10\] VGND VGND VPWR VPWR _02841_
+ sky130_fd_sc_hd__a22o_1
X_09037_ net403 net2266 net513 VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11149__B2 net804 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08014__A1 net1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold350 cpuregs\[12\]\[17\] VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__X _03852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout591_X net591 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold361 cpuregs\[28\]\[22\] VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 cpuregs\[16\]\[26\] VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold383 cpuregs\[29\]\[15\] VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__A1 net984 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold394 cpuregs\[14\]\[14\] VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout830 _03137_ VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout841 net842 VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__buf_2
XFILLER_120_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout852 _02468_ VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__buf_2
X_09939_ net1127 _04447_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__xor2_1
Xfanout863 net865 VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__buf_2
XANTENNA_fanout856_X net856 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout874 _05082_ VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__clkbuf_4
Xfanout885 net891 VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__buf_2
XANTENNA__11029__A net1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ net342 net1944 net452 VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__mux2_1
Xfanout896 net897 VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07525__B1 net979 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1050 genblk1.genblk1.pcpi_mul.next_rs1\[17\] VGND VGND VPWR VPWR net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 genblk1.genblk1.pcpi_mul.next_rs1\[53\] VGND VGND VPWR VPWR net2375 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _06370_ _06371_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__nand2b_1
XFILLER_18_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1072 cpuregs\[10\]\[29\] VGND VGND VPWR VPWR net2386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__B net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12881_ mem_rdata_q\[18\] net10 net962 VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__mux2_1
Xhold1083 cpuregs\[5\]\[26\] VGND VGND VPWR VPWR net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 cpuregs\[11\]\[8\] VGND VGND VPWR VPWR net2408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14620_ clknet_leaf_93_clk _01006_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
X_11832_ genblk2.pcpi_div.divisor\[10\] genblk2.pcpi_div.dividend\[10\] VGND VGND
+ VPWR VPWR _06303_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_116_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09817__A2 net876 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ clknet_leaf_184_clk _00937_ VGND VGND VPWR VPWR cpuregs\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11763_ net1761 net117 net730 VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__mux2_1
XFILLER_26_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10714_ net780 _05394_ _05403_ net777 VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__o211a_1
X_13502_ net1707 net345 net420 VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__mux2_1
X_14482_ clknet_leaf_93_clk _00871_ VGND VGND VPWR VPWR instr_addi sky130_fd_sc_hd__dfxtp_1
X_11694_ net1747 net406 net373 VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__mux2_1
XFILLER_41_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13433_ net1005 net756 _02336_ net710 VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__o211a_1
X_10645_ _05335_ _05336_ net814 VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__mux2_1
XANTENNA__11388__A1 net832 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13364_ net569 _05784_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__nor2_1
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10576_ cpuregs\[20\]\[6\] cpuregs\[21\]\[6\] net670 VGND VGND VPWR VPWR _05270_
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15103_ clknet_leaf_16_clk _01455_ VGND VGND VPWR VPWR cpuregs\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12315_ net3055 net743 _06632_ _06636_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_125_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13295_ net960 _04983_ _02214_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__nor3_1
X_15034_ clknet_leaf_135_clk _01386_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12246_ net2661 net379 net366 net2742 VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__a22o_1
XFILLER_107_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12888__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12177_ net2750 net276 net2908 VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09108__S net505 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11128_ cpuregs\[25\]\[21\] net622 net605 _05806_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__o211a_1
XFILLER_111_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11059_ cpuregs\[28\]\[19\] cpuregs\[29\]\[19\] net681 VGND VGND VPWR VPWR _05740_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07136__B net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08947__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14818_ clknet_leaf_82_clk _01170_ VGND VGND VPWR VPWR decoded_imm\[4\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_121_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14749_ clknet_leaf_155_clk net2874 VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08270_ reg_out\[12\] reg_next_pc\[12\] net920 VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__mux2_1
XFILLER_33_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07221_ net1139 count_cycle\[37\] net976 _02768_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__a211o_1
XANTENNA__13368__A2 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10717__S net802 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08244__A1 net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07152_ _02700_ net842 _02704_ _02696_ net1060 VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__a32o_1
XANTENNA__12040__A2 net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07083_ net1121 genblk2.pcpi_div.quotient\[23\] _02644_ net953 VGND VGND VPWR VPWR
+ _02646_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_8_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12879__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13329__A net960 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09018__S net519 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07985_ _03311_ _03496_ _03497_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout384_A net390 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09724_ net984 _04516_ _04517_ _02380_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__a31o_1
X_06936_ _02516_ _02517_ _02519_ net953 VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09655_ net848 _04454_ _04455_ net878 net1330 VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__a32o_1
X_06867_ net2132 _02467_ _02469_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__a21o_1
XANTENNA__12379__S net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout649_A net654 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08606_ _03979_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__nand2_1
X_09586_ _04418_ _04419_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__nor2_1
XANTENNA__13056__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_06798_ net1024 VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__inv_2
XFILLER_169_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08537_ _03922_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1081_X net1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10200__B net1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_964 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout816_A net818 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1179_X net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08468_ reg_out\[30\] alu_out_q\[30\] net1156 VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__mux2_1
XFILLER_24_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08483__B2 net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ _02923_ _02941_ _02939_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__o21ai_1
X_08399_ net336 net2315 net528 VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__mux2_1
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13003__S net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10430_ net3008 _05121_ net410 VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__a21o_1
XANTENNA__08235__A1 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ cpuregs\[30\]\[31\] cpuregs\[31\]\[31\] net694 VGND VGND VPWR VPWR _05067_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12842__S net460 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12100_ genblk2.pcpi_div.dividend\[25\] net273 _06545_ VGND VGND VPWR VPWR _01034_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13080_ net346 net1682 net440 VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__mux2_1
X_10292_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__inv_2
XFILLER_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11458__S net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12031_ net1019 net722 _06484_ net862 VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__a31o_1
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold180 net42 VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 cpuregs\[24\]\[12\] VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout660 net663 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkbuf_2
Xfanout671 net672 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__buf_2
XANTENNA__11982__A net1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout682 net683 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__buf_2
Xfanout693 net694 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__buf_2
X_13982_ clknet_leaf_10_clk _00436_ VGND VGND VPWR VPWR cpuregs\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_92_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12933_ _03192_ _05204_ _02121_ _02502_ net2170 VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__o32a_1
XANTENNA__10598__A net815 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15652_ clknet_leaf_53_clk _01988_ VGND VGND VPWR VPWR cpuregs\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__13047__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ net12 net2645 _02450_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__mux2_1
X_14603_ clknet_leaf_117_clk _00989_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dfxtp_1
X_11815_ _06283_ _06285_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__nor2_1
X_12795_ _02414_ _02115_ net918 VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__a21oi_1
X_15583_ clknet_leaf_58_clk _01919_ VGND VGND VPWR VPWR cpuregs\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10805__B1 net854 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14534_ clknet_leaf_87_clk _00001_ VGND VGND VPWR VPWR is_lui_auipc_jal sky130_fd_sc_hd__dfxtp_2
X_11746_ net1642 net99 net730 VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__mux2_1
X_11677_ net29 _06226_ net27 net28 VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__or4b_1
X_14465_ clknet_leaf_89_clk _00854_ VGND VGND VPWR VPWR instr_lui sky130_fd_sc_hd__dfxtp_1
XFILLER_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12558__B1 net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13416_ net1002 net757 VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__or2_1
XANTENNA__08226__A1 net1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10628_ cpuregs\[4\]\[8\] cpuregs\[5\]\[8\] net677 VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__mux2_1
X_14396_ clknet_leaf_102_clk _00817_ VGND VGND VPWR VPWR pcpi_timeout_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08226__B2 net942 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13347_ net568 _05710_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__nor2_1
XANTENNA__11230__B1 net601 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10559_ cpuregs\[12\]\[6\] cpuregs\[13\]\[6\] net673 VGND VGND VPWR VPWR _05253_
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13278_ _04933_ _04975_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__nand2_1
XFILLER_170_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15017_ clknet_leaf_106_clk net2528 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rs2\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12229_ genblk2.pcpi_div.quotient_msk\[28\] net274 net2806 VGND VGND VPWR VPWR _06607_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_96_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12730__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13583__S net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_142_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07770_ _03286_ _03287_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__and2_2
X_09440_ count_instr\[11\] count_instr\[10\] count_instr\[9\] _04318_ VGND VGND VPWR
+ VPWR _04325_ sky130_fd_sc_hd__and4_1
XANTENNA__13038__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11049__B1 _03171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09371_ net1823 net524 net399 VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__mux2_1
XFILLER_52_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12927__S net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08322_ net587 net2216 net530 VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__mux2_1
XANTENNA__08265__X net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12261__A2 net381 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_151_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09301__S net480 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13331__B net759 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08253_ net1044 _03710_ net981 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__mux2_2
XFILLER_165_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12228__A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07204_ net203 net1057 _02752_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__and3_1
XANTENNA__08217__A1 net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08184_ _03289_ _03295_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__nand2_1
XANTENNA__08217__B2 net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13210__A1 net1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09965__A1 net1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10393__D net1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11221__B1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07135_ net1048 net1054 VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__nand2_4
XANTENNA__11772__A1 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07066_ genblk2.pcpi_div.dividend\[20\] _02622_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__or2_1
XFILLER_160_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput230 net1041 VGND VGND VPWR VPWR pcpi_rs1[5] sky130_fd_sc_hd__buf_2
Xoutput241 net1162 VGND VGND VPWR VPWR pcpi_rs2[15] sky130_fd_sc_hd__buf_2
XFILLER_88_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput252 net252 VGND VGND VPWR VPWR pcpi_rs2[25] sky130_fd_sc_hd__buf_2
XANTENNA_fanout599_A net600 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput263 net263 VGND VGND VPWR VPWR pcpi_rs2[6] sky130_fd_sc_hd__buf_2
XFILLER_160_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_160_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13493__S net419 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A _03747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07968_ _03275_ _03482_ _03465_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06919_ genblk2.pcpi_div.instr_div genblk2.pcpi_div.instr_rem VGND VGND VPWR VPWR
+ _02507_ sky130_fd_sc_hd__or2_2
XFILLER_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09707_ decoded_imm_j\[7\] _04428_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__and2_1
X_07899_ net1165 _02404_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout554_X net554 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11307__A net794 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09638_ _03845_ reg_next_pc\[25\] net924 VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__mux2_2
XANTENNA__10211__A decoded_imm\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ net2889 _04406_ net1240 VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout721_X net721 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12837__S net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_X net819 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11600_ is_alu_reg_imm _06183_ _06200_ net741 instr_srli VGND VGND VPWR VPWR _00879_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__11741__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12580_ net527 net1922 net467 VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__mux2_1
XANTENNA__07259__A2 _02799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12252__A2 net377 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10865__B net664 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09211__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11531_ mem_rdata_q\[24\] net1589 net737 VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_129_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11460__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11042__A net816 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14250_ clknet_leaf_68_clk _00704_ VGND VGND VPWR VPWR reg_next_pc\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11462_ cpuregs\[18\]\[30\] net554 _06131_ net783 VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__o22a_1
X_13201_ net1063 _02474_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__and2_2
X_10413_ net256 net255 _05117_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__or3_1
X_14181_ clknet_leaf_109_clk _00635_ VGND VGND VPWR VPWR count_instr\[52\] sky130_fd_sc_hd__dfxtp_1
X_11393_ cpuregs\[17\]\[28\] net636 net612 _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__o211a_1
X_13132_ _04273_ _02127_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__nor2_1
XFILLER_125_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10344_ cpuregs\[12\]\[31\] cpuregs\[13\]\[31\] net694 VGND VGND VPWR VPWR _05050_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13063_ net1439 net87 net533 VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__mux2_1
XFILLER_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10275_ _04934_ _04935_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__and2b_1
X_12014_ net1025 net721 _06470_ _06471_ net862 VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__a311o_1
XANTENNA__12712__B1 net914 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07195__A1 net1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 _04287_ VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_8
XFILLER_94_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__06942__B2 net949 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13416__B net757 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13965_ clknet_leaf_56_clk _00419_ VGND VGND VPWR VPWR cpuregs\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12916_ net323 net2034 net456 VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload8_A clknet_4_8_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_59_clk _00350_ VGND VGND VPWR VPWR cpuregs\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15635_ clknet_leaf_196_clk _01971_ VGND VGND VPWR VPWR cpuregs\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12847_ net337 net2306 net459 VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__mux2_1
XFILLER_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15566_ clknet_leaf_182_clk _01902_ VGND VGND VPWR VPWR cpuregs\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__12243__A2 net382 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12778_ net1221 genblk1.genblk1.pcpi_mul.next_rs1\[46\] net2233 net909 net765 VGND
+ VGND VPWR VPWR _01417_ sky130_fd_sc_hd__a221o_1
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09121__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11451__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14517_ clknet_leaf_77_clk _00906_ VGND VGND VPWR VPWR decoded_imm_j\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_155_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ latched_rd\[0\] _06242_ _06243_ net1740 VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a22o_1
X_15497_ clknet_leaf_132_clk _01833_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dfxtp_2
XANTENNA__08960__S net955 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14448_ clknet_leaf_42_clk _00837_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dfxtp_1
XANTENNA__13578__S net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07407__C1 net991 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09947__B2 net849 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold905 cpuregs\[21\]\[26\] VGND VGND VPWR VPWR net2219 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ clknet_leaf_131_clk _00800_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dfxtp_4
Xhold916 cpuregs\[17\]\[23\] VGND VGND VPWR VPWR net2230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07958__B1 net1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold927 cpuregs\[2\]\[23\] VGND VGND VPWR VPWR net2241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold938 cpuregs\[19\]\[26\] VGND VGND VPWR VPWR net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold949 cpuregs\[25\]\[30\] VGND VGND VPWR VPWR net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_08940_ genblk1.genblk1.pcpi_mul.rd\[8\] genblk1.genblk1.pcpi_mul.rd\[40\] net954
+ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__mux2_1
X_08871_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__inv_2
XANTENNA__10714__C1 net777 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1605 genblk1.genblk1.pcpi_mul.rd\[31\] VGND VGND VPWR VPWR net2919 sky130_fd_sc_hd__dlygate4sd3_1
X_07822_ _03336_ _03339_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__or2_1
Xhold1616 instr_lbu VGND VGND VPWR VPWR net2930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1627 genblk1.genblk1.pcpi_mul.rd\[63\] VGND VGND VPWR VPWR net2941 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13259__A1 net1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1638 genblk1.genblk1.pcpi_mul.next_rs2\[56\] VGND VGND VPWR VPWR net2952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1649 genblk1.genblk1.pcpi_mul.next_rs2\[60\] VGND VGND VPWR VPWR net2963 sky130_fd_sc_hd__dlygate4sd3_1
X_07753_ _03269_ _03270_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__and2_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07324__B decoded_imm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07684_ net810 _03201_ _03203_ net825 VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__o211a_1
X_09423_ _04313_ net1231 _04311_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__and3b_1
XFILLER_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13342__A net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_A cpu_state\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09354_ net1378 net310 net477 VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__mux2_1
X_08305_ net994 _03736_ net982 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09031__S net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11442__B1 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09285_ net2177 net312 net486 VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__mux2_1
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout514_A net515 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08236_ net1176 net1159 net940 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__mux2_1
XANTENNA__10650__D1 net789 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13488__S net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08167_ _03295_ net935 VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__nor2_1
XANTENNA__12392__S net474 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout1044_X net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07118_ net1123 _02669_ genblk2.pcpi_div.dividend\[29\] VGND VGND VPWR VPWR _02675_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08098_ _03337_ net932 _03588_ _03597_ VGND VGND VPWR VPWR alu_out\[18\] sky130_fd_sc_hd__a211o_1
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout883_A net898 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07049_ _02615_ _02616_ _02613_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13498__A1 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10060_ net3038 _04804_ net1236 VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11736__S net729 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09206__S net492 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__15505__Q net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__15732__A net1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13750_ clknet_leaf_182_clk _00204_ VGND VGND VPWR VPWR cpuregs\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10962_ cpuregs\[2\]\[17\] net659 VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__or2_1
XFILLER_83_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09730__A decoded_imm_j\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12701_ net1199 net1098 net897 net2772 _02084_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__a221o_1
XFILLER_43_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12567__S net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10876__A net772 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10893_ cpuregs\[9\]\[15\] net618 net603 _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__o211a_1
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13681_ clknet_leaf_118_clk _00135_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15420_ clknet_leaf_35_clk _01759_ VGND VGND VPWR VPWR cpuregs\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12632_ net1192 net2814 net885 genblk1.genblk1.pcpi_mul.next_rs2\[14\] _02065_ VGND
+ VGND VPWR VPWR _01320_ sky130_fd_sc_hd__a221o_1
XANTENNA__12225__A2 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12563_ _02044_ net2627 net390 VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__mux2_1
X_15351_ clknet_leaf_43_clk _01691_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11514_ mem_rdata_q\[7\] net2055 net736 VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__mux2_1
X_14302_ clknet_leaf_110_clk _00756_ VGND VGND VPWR VPWR count_cycle\[47\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11984__B2 net867 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15282_ clknet_leaf_7_clk _01623_ VGND VGND VPWR VPWR cpuregs\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12494_ genblk2.pcpi_div.divisor\[45\] net871 VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__nor2_1
XFILLER_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11445_ net832 _06110_ _06114_ net783 VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__a211o_1
X_14233_ clknet_leaf_173_clk _00687_ VGND VGND VPWR VPWR reg_next_pc\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11736__A1 net1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14164_ clknet_leaf_126_clk _00618_ VGND VGND VPWR VPWR count_instr\[35\] sky130_fd_sc_hd__dfxtp_1
X_11376_ cpuregs\[9\]\[28\] net637 net612 _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__o211a_1
XFILLER_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output266_A net1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10327_ _04894_ _04895_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__nor2_1
X_13115_ net337 net2213 net436 VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__mux2_1
XFILLER_124_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14095_ clknet_leaf_47_clk _00549_ VGND VGND VPWR VPWR cpuregs\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ net1352 net69 net534 VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__mux2_1
XFILLER_3_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09905__A net1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10258_ decoded_imm\[6\] net1038 _04940_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__nand3_1
XANTENNA__07168__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout1230 net1241 VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11646__S net545 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07168__B2 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1241 net34 VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__buf_2
X_10189_ decoded_imm\[29\] net994 VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__and2_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09116__S net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14997_ clknet_leaf_148_clk _01349_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs2\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13948_ clknet_leaf_191_clk _00402_ VGND VGND VPWR VPWR cpuregs\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_47_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08955__S net943 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10475__A1 net806 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13879_ clknet_leaf_185_clk _00333_ VGND VGND VPWR VPWR cpuregs\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15618_ clknet_leaf_46_clk _01954_ VGND VGND VPWR VPWR cpuregs\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__07628__C1 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15549_ clknet_leaf_17_clk _01885_ VGND VGND VPWR VPWR cpuregs\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_170_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09070_ net1930 net407 net509 VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08021_ _03522_ _03528_ _03349_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10725__S net814 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap410 _02455_ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11410__A net808 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold702 cpuregs\[6\]\[22\] VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13101__S net437 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold713 cpuregs\[5\]\[23\] VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 cpuregs\[7\]\[6\] VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 cpuregs\[19\]\[10\] VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 cpuregs\[10\]\[16\] VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 cpuregs\[31\]\[0\] VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 cpuregs\[23\]\[26\] VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 cpuregs\[31\]\[26\] VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _04741_ _04744_ net1152 VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12940__S net454 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08923_ net1213 net2665 net901 _04238_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__a22o_1
XFILLER_131_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12688__C1 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A _03852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09093__Y _04279_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1402 _01112_ VGND VGND VPWR VPWR net2716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 instr_or VGND VGND VPWR VPWR net2727 sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ _04188_ _04190_ _04183_ _04186_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__a211o_1
Xhold1424 _00828_ VGND VGND VPWR VPWR net2738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout1004_A net1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06906__B2 net1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1435 genblk1.genblk1.pcpi_mul.rd\[9\] VGND VGND VPWR VPWR net2749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 mem_state\[0\] VGND VGND VPWR VPWR net2760 sky130_fd_sc_hd__dlygate4sd3_1
X_07805_ _03319_ _03321_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__nor2_1
Xhold1457 genblk2.pcpi_div.divisor\[32\] VGND VGND VPWR VPWR net2771 sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ net885 _04130_ _04132_ net2697 net1194 VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__a32o_1
Xhold1468 genblk2.pcpi_div.divisor\[26\] VGND VGND VPWR VPWR net2782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08108__B1 net969 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1479 mem_rdata_q\[3\] VGND VGND VPWR VPWR net2793 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout464_A _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07736_ cpuregs\[20\]\[4\] cpuregs\[21\]\[4\] net701 VGND VGND VPWR VPWR _03255_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07622__X _03143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11663__A0 decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12387__S net362 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07667_ net837 _03183_ _03185_ _03187_ net794 VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__a2111o_1
XFILLER_41_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout631_A net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06893__B _02479_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout729_A net730 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09406_ net1089 count_instr\[0\] net1184 VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__and3_1
X_07598_ count_instr\[30\] net1137 net978 _03120_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__a211o_1
XFILLER_125_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12207__A2 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11415__B1 net602 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09337_ net1617 net539 net475 VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1161_X net1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_X net517 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10769__A2 decoded_imm\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07095__B1 net952 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09268_ net2087 net543 net487 VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__mux2_1
XANTENNA__08831__A1 net900 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07634__A2 net640 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08219_ net1058 net1179 net266 net1054 VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__a22o_1
XFILLER_153_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09199_ net2007 net582 net494 VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__mux2_1
XFILLER_147_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13011__S net443 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11230_ cpuregs\[19\]\[24\] net640 net601 VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__o21a_1
XFILLER_153_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11194__A2 net630 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__15727__A net1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11161_ cpuregs\[30\]\[22\] cpuregs\[31\]\[22\] net683 VGND VGND VPWR VPWR _05839_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07229__B decoded_imm\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12850__S net461 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10112_ count_cycle\[41\] count_cycle\[42\] _04836_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__and3_1
XFILLER_161_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12679__C1 net711 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11092_ cpuregs\[2\]\[20\] cpuregs\[3\]\[20\] net661 VGND VGND VPWR VPWR _05772_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11466__S net805 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10043_ _04791_ _04795_ _04794_ net1206 VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a211oi_1
X_14920_ clknet_leaf_109_clk _01272_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13247__A net1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold40 genblk1.genblk1.pcpi_mul.next_rs1\[7\] VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold51 _01376_ VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 cpuregs\[26\]\[3\] VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A mem_rdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14851_ clknet_leaf_51_clk _01203_ VGND VGND VPWR VPWR cpuregs\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold73 cpuregs\[26\]\[2\] VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold84 net145 VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold95 cpuregs\[12\]\[11\] VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_47_clk _00256_ VGND VGND VPWR VPWR cpuregs\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_14782_ clknet_leaf_155_clk _00037_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[29\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__10877__Y _05563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11994_ net862 _06454_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__nor2_1
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10457__B2 net784 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13733_ clknet_leaf_112_clk _00187_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10945_ cpuregs\[28\]\[16\] cpuregs\[29\]\[16\] net656 VGND VGND VPWR VPWR _05629_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13664_ clknet_leaf_119_clk _00118_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_10876_ net772 _05553_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__and3_1
XFILLER_71_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15403_ clknet_leaf_20_clk _01742_ VGND VGND VPWR VPWR cpuregs\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12615_ net1201 genblk1.genblk1.pcpi_mul.next_rs2\[7\] net916 net125 VGND VGND VPWR
+ VPWR _02057_ sky130_fd_sc_hd__a22o_1
XANTENNA__11214__B _05890_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ clknet_leaf_39_clk _00050_ VGND VGND VPWR VPWR cpuregs\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11957__A1 net726 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15334_ clknet_leaf_156_clk _01674_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_1
X_12546_ _02031_ net2722 net390 VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__mux2_1
X_15265_ clknet_leaf_57_clk _01606_ VGND VGND VPWR VPWR cpuregs\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12477_ net1166 net715 _05102_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_113_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12906__A0 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output93_A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14216_ clknet_leaf_75_clk _00670_ VGND VGND VPWR VPWR reg_pc\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11428_ cpuregs\[16\]\[29\] net706 VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__or2_1
XFILLER_125_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15196_ clknet_leaf_6_clk _01545_ VGND VGND VPWR VPWR cpuregs\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11185__A2 net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14147_ clknet_leaf_97_clk _00601_ VGND VGND VPWR VPWR count_instr\[18\] sky130_fd_sc_hd__dfxtp_1
X_11359_ cpuregs\[18\]\[27\] net554 _06031_ net784 VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__o22a_1
XFILLER_125_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_956 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14078_ clknet_leaf_7_clk _00532_ VGND VGND VPWR VPWR cpuregs\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_13029_ net299 net2510 net445 VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__mux2_1
XFILLER_112_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1060 net1062 VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__buf_2
XFILLER_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1071 net1074 VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_2_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1082 net1086 VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1109 VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__clkbuf_2
XFILLER_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08570_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__inv_2
XFILLER_82_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07521_ _03035_ _03037_ _03048_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__a21o_1
XANTENNA__11645__A0 decoded_imm_j\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07452_ net13 net939 net936 VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__a21oi_1
XFILLER_168_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07383_ net842 _02917_ _02918_ _02909_ net1071 VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__a32o_1
XANTENNA__12935__S net453 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09122_ net2373 net289 net506 VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__mux2_1
XANTENNA__07616__A2 decoded_imm_j\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08273__X net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09053_ net297 net2457 net514 VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__mux2_1
XANTENNA__12236__A net750 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08004_ net967 _03353_ _03354_ net928 _03513_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__a221o_1
XANTENNA__11140__A net774 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold510 cpuregs\[13\]\[9\] VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 cpuregs\[21\]\[18\] VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 cpuregs\[6\]\[6\] VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 cpuregs\[13\]\[14\] VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold554 cpuregs\[16\]\[25\] VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold565 cpuregs\[4\]\[12\] VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold576 net140 VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 cpuregs\[8\]\[24\] VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 cpuregs\[21\]\[16\] VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _04726_ _04727_ _04728_ _04729_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout581_A _03753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__06888__B is_beq_bne_blt_bge_bltu_bgeu VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A _03139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08906_ _04024_ _04026_ _04023_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__a21bo_1
X_09886_ _04638_ _04653_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1007_X net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1210 cpuregs\[1\]\[2\] VGND VGND VPWR VPWR net2524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11333__C1 net833 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1221 genblk2.pcpi_div.divisor\[57\] VGND VGND VPWR VPWR net2535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 genblk2.pcpi_div.divisor\[37\] VGND VGND VPWR VPWR net2546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 instr_lui VGND VGND VPWR VPWR net2557 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net900 _04174_ _04176_ net2755 net1211 VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_51_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout467_X net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1254 genblk1.genblk1.pcpi_mul.pcpi_rd\[15\] VGND VGND VPWR VPWR net2568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout846_A net852 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10203__B net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1265 genblk2.pcpi_div.divisor\[0\] VGND VGND VPWR VPWR net2579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 count_instr\[53\] VGND VGND VPWR VPWR net2590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 genblk1.genblk1.pcpi_mul.pcpi_rd\[14\] VGND VGND VPWR VPWR net2601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 net196 VGND VGND VPWR VPWR net2612 sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ genblk1.genblk1.pcpi_mul.rd\[44\] genblk1.genblk1.pcpi_mul.rdx\[44\] VGND
+ VGND VPWR VPWR _04118_ sky130_fd_sc_hd__or2_1
X_07719_ cpuregs\[14\]\[4\] cpuregs\[15\]\[4\] net698 VGND VGND VPWR VPWR _03238_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout634_X net634 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08699_ _04051_ _04054_ _04056_ _04058_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__o211a_1
XANTENNA__13006__S net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10730_ net827 _05415_ _05417_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__a211o_1
XFILLER_159_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10661_ net1076 _05351_ net853 VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12845__S net460 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout801_X net801 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07068__B1 net947 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12400_ net522 net2135 net471 VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__mux2_1
XFILLER_167_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13380_ net1000 net760 VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__or2_1
X_10592_ cpuregs\[1\]\[7\] net630 net609 _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__o211a_1
XANTENNA__11969__B net1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12331_ decoded_imm\[9\] net735 _06643_ mem_rdata_q\[29\] _06645_ VGND VGND VPWR
+ VPWR _01165_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_58_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15050_ clknet_leaf_102_clk net2338 VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.next_rs1\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_12262_ net2775 net381 net369 net2782 VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13561__A0 net524 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12364__A1 net540 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14001_ clknet_leaf_21_clk _00455_ VGND VGND VPWR VPWR cpuregs\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11213_ net774 _05865_ _05873_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__a31oi_4
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12193_ net2798 net272 net2801 VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12580__S net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10375__B1 net566 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput41 net41 VGND VGND VPWR VPWR mem_addr[16] sky130_fd_sc_hd__buf_2
Xoutput52 net52 VGND VGND VPWR VPWR mem_addr[27] sky130_fd_sc_hd__buf_2
XFILLER_150_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11144_ net248 net859 _05821_ _05822_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__a22o_1
XFILLER_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput63 net63 VGND VGND VPWR VPWR mem_addr[8] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VGND VGND VPWR VPWR mem_la_addr[18] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VGND VGND VPWR VPWR mem_la_addr[29] sky130_fd_sc_hd__buf_2
Xoutput96 net96 VGND VGND VPWR VPWR mem_la_read sky130_fd_sc_hd__buf_2
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11075_ cpuregs\[25\]\[20\] net622 net605 _05754_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__o211a_1
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10678__A1 net780 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14903_ clknet_leaf_143_clk _01255_ VGND VGND VPWR VPWR genblk2.pcpi_div.divisor\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10026_ count_cycle\[10\] count_cycle\[11\] _04781_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__and3_1
XANTENNA_input28_X net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output131_A net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07543__A1 net1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07543__B2 net978 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output229_A net229 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14834_ clknet_leaf_192_clk _01186_ VGND VGND VPWR VPWR cpuregs\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ clknet_leaf_163_clk _00019_ VGND VGND VPWR VPWR genblk2.pcpi_div.pcpi_rd\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08099__A2 net1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11977_ net1036 _06440_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__nand2_1
XFILLER_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13716_ clknet_leaf_140_clk _00170_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.pcpi_rd\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10928_ net798 _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__or2_1
X_14696_ clknet_leaf_152_clk _01081_ VGND VGND VPWR VPWR genblk2.pcpi_div.quotient\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13647_ clknet_leaf_143_clk _00101_ VGND VGND VPWR VPWR genblk1.genblk1.pcpi_mul.rd\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10859_ net787 _05540_ _05542_ _05544_ net777 VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__o41a_1
XANTENNA__09599__A2 net877 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13578_ net306 net2359 net414 VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__mux2_1
X_15317_ clknet_leaf_11_clk _01657_ VGND VGND VPWR VPWR cpuregs\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12529_ genblk2.pcpi_div.divisor\[52\] _02018_ net872 VGND VGND VPWR VPWR _02019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15248_ clknet_leaf_16_clk _01589_ VGND VGND VPWR VPWR cpuregs\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12355__B2 net917 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15179_ clknet_leaf_91_clk _01528_ VGND VGND VPWR VPWR mem_rdata_q\[30\] sky130_fd_sc_hd__dfxtp_4
XFILLER_126_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07437__X _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout308 net311 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_2
Xfanout319 _03831_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09508__C1 net1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09740_ net1183 _04430_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__or2_1
X_06952_ genblk2.pcpi_div.quotient\[4\] _02525_ net1125 VGND VGND VPWR VPWR _02533_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__14421__D alu_out\[21\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

