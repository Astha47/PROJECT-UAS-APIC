module picorv32 (clk,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    pcpi_ready,
    pcpi_valid,
    pcpi_wait,
    pcpi_wr,
    resetn,
    trace_valid,
    trap,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    pcpi_insn,
    pcpi_rd,
    pcpi_rs1,
    pcpi_rs2,
    trace_data);
 input clk;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input pcpi_ready;
 output pcpi_valid;
 input pcpi_wait;
 input pcpi_wr;
 input resetn;
 output trace_valid;
 output trap;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [31:0] pcpi_insn;
 input [31:0] pcpi_rd;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 output [35:0] trace_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire \alu_out[0] ;
 wire \alu_out[10] ;
 wire \alu_out[11] ;
 wire \alu_out[12] ;
 wire \alu_out[13] ;
 wire \alu_out[14] ;
 wire \alu_out[15] ;
 wire \alu_out[16] ;
 wire \alu_out[17] ;
 wire \alu_out[18] ;
 wire \alu_out[19] ;
 wire \alu_out[1] ;
 wire \alu_out[20] ;
 wire \alu_out[21] ;
 wire \alu_out[22] ;
 wire \alu_out[23] ;
 wire \alu_out[24] ;
 wire \alu_out[25] ;
 wire \alu_out[26] ;
 wire \alu_out[27] ;
 wire \alu_out[28] ;
 wire \alu_out[29] ;
 wire \alu_out[2] ;
 wire \alu_out[30] ;
 wire \alu_out[31] ;
 wire \alu_out[3] ;
 wire \alu_out[4] ;
 wire \alu_out[5] ;
 wire \alu_out[6] ;
 wire \alu_out[7] ;
 wire \alu_out[8] ;
 wire \alu_out[9] ;
 wire \alu_out_q[0] ;
 wire \alu_out_q[10] ;
 wire \alu_out_q[11] ;
 wire \alu_out_q[12] ;
 wire \alu_out_q[13] ;
 wire \alu_out_q[14] ;
 wire \alu_out_q[15] ;
 wire \alu_out_q[16] ;
 wire \alu_out_q[17] ;
 wire \alu_out_q[18] ;
 wire \alu_out_q[19] ;
 wire \alu_out_q[1] ;
 wire \alu_out_q[20] ;
 wire \alu_out_q[21] ;
 wire \alu_out_q[22] ;
 wire \alu_out_q[23] ;
 wire \alu_out_q[24] ;
 wire \alu_out_q[25] ;
 wire \alu_out_q[26] ;
 wire \alu_out_q[27] ;
 wire \alu_out_q[28] ;
 wire \alu_out_q[29] ;
 wire \alu_out_q[2] ;
 wire \alu_out_q[30] ;
 wire \alu_out_q[31] ;
 wire \alu_out_q[3] ;
 wire \alu_out_q[4] ;
 wire \alu_out_q[5] ;
 wire \alu_out_q[6] ;
 wire \alu_out_q[7] ;
 wire \alu_out_q[8] ;
 wire \alu_out_q[9] ;
 wire \count_cycle[0] ;
 wire \count_cycle[10] ;
 wire \count_cycle[11] ;
 wire \count_cycle[12] ;
 wire \count_cycle[13] ;
 wire \count_cycle[14] ;
 wire \count_cycle[15] ;
 wire \count_cycle[16] ;
 wire \count_cycle[17] ;
 wire \count_cycle[18] ;
 wire \count_cycle[19] ;
 wire \count_cycle[1] ;
 wire \count_cycle[20] ;
 wire \count_cycle[21] ;
 wire \count_cycle[22] ;
 wire \count_cycle[23] ;
 wire \count_cycle[24] ;
 wire \count_cycle[25] ;
 wire \count_cycle[26] ;
 wire \count_cycle[27] ;
 wire \count_cycle[28] ;
 wire \count_cycle[29] ;
 wire \count_cycle[2] ;
 wire \count_cycle[30] ;
 wire \count_cycle[31] ;
 wire \count_cycle[32] ;
 wire \count_cycle[33] ;
 wire \count_cycle[34] ;
 wire \count_cycle[35] ;
 wire \count_cycle[36] ;
 wire \count_cycle[37] ;
 wire \count_cycle[38] ;
 wire \count_cycle[39] ;
 wire \count_cycle[3] ;
 wire \count_cycle[40] ;
 wire \count_cycle[41] ;
 wire \count_cycle[42] ;
 wire \count_cycle[43] ;
 wire \count_cycle[44] ;
 wire \count_cycle[45] ;
 wire \count_cycle[46] ;
 wire \count_cycle[47] ;
 wire \count_cycle[48] ;
 wire \count_cycle[49] ;
 wire \count_cycle[4] ;
 wire \count_cycle[50] ;
 wire \count_cycle[51] ;
 wire \count_cycle[52] ;
 wire \count_cycle[53] ;
 wire \count_cycle[54] ;
 wire \count_cycle[55] ;
 wire \count_cycle[56] ;
 wire \count_cycle[57] ;
 wire \count_cycle[58] ;
 wire \count_cycle[59] ;
 wire \count_cycle[5] ;
 wire \count_cycle[60] ;
 wire \count_cycle[61] ;
 wire \count_cycle[62] ;
 wire \count_cycle[63] ;
 wire \count_cycle[6] ;
 wire \count_cycle[7] ;
 wire \count_cycle[8] ;
 wire \count_cycle[9] ;
 wire \count_instr[0] ;
 wire \count_instr[10] ;
 wire \count_instr[11] ;
 wire \count_instr[12] ;
 wire \count_instr[13] ;
 wire \count_instr[14] ;
 wire \count_instr[15] ;
 wire \count_instr[16] ;
 wire \count_instr[17] ;
 wire \count_instr[18] ;
 wire \count_instr[19] ;
 wire \count_instr[1] ;
 wire \count_instr[20] ;
 wire \count_instr[21] ;
 wire \count_instr[22] ;
 wire \count_instr[23] ;
 wire \count_instr[24] ;
 wire \count_instr[25] ;
 wire \count_instr[26] ;
 wire \count_instr[27] ;
 wire \count_instr[28] ;
 wire \count_instr[29] ;
 wire \count_instr[2] ;
 wire \count_instr[30] ;
 wire \count_instr[31] ;
 wire \count_instr[32] ;
 wire \count_instr[33] ;
 wire \count_instr[34] ;
 wire \count_instr[35] ;
 wire \count_instr[36] ;
 wire \count_instr[37] ;
 wire \count_instr[38] ;
 wire \count_instr[39] ;
 wire \count_instr[3] ;
 wire \count_instr[40] ;
 wire \count_instr[41] ;
 wire \count_instr[42] ;
 wire \count_instr[43] ;
 wire \count_instr[44] ;
 wire \count_instr[45] ;
 wire \count_instr[46] ;
 wire \count_instr[47] ;
 wire \count_instr[48] ;
 wire \count_instr[49] ;
 wire \count_instr[4] ;
 wire \count_instr[50] ;
 wire \count_instr[51] ;
 wire \count_instr[52] ;
 wire \count_instr[53] ;
 wire \count_instr[54] ;
 wire \count_instr[55] ;
 wire \count_instr[56] ;
 wire \count_instr[57] ;
 wire \count_instr[58] ;
 wire \count_instr[59] ;
 wire \count_instr[5] ;
 wire \count_instr[60] ;
 wire \count_instr[61] ;
 wire \count_instr[62] ;
 wire \count_instr[63] ;
 wire \count_instr[6] ;
 wire \count_instr[7] ;
 wire \count_instr[8] ;
 wire \count_instr[9] ;
 wire \cpu_state[0] ;
 wire \cpu_state[1] ;
 wire \cpu_state[2] ;
 wire \cpu_state[3] ;
 wire \cpu_state[4] ;
 wire \cpu_state[5] ;
 wire \cpu_state[6] ;
 wire \cpu_state[7] ;
 wire \cpuregs[0][0] ;
 wire \cpuregs[0][16] ;
 wire \cpuregs[0][17] ;
 wire \cpuregs[0][19] ;
 wire \cpuregs[0][25] ;
 wire \cpuregs[0][2] ;
 wire \cpuregs[0][30] ;
 wire \cpuregs[0][31] ;
 wire \cpuregs[0][7] ;
 wire \cpuregs[10][0] ;
 wire \cpuregs[10][10] ;
 wire \cpuregs[10][11] ;
 wire \cpuregs[10][12] ;
 wire \cpuregs[10][13] ;
 wire \cpuregs[10][14] ;
 wire \cpuregs[10][15] ;
 wire \cpuregs[10][16] ;
 wire \cpuregs[10][17] ;
 wire \cpuregs[10][18] ;
 wire \cpuregs[10][19] ;
 wire \cpuregs[10][1] ;
 wire \cpuregs[10][20] ;
 wire \cpuregs[10][21] ;
 wire \cpuregs[10][22] ;
 wire \cpuregs[10][23] ;
 wire \cpuregs[10][24] ;
 wire \cpuregs[10][25] ;
 wire \cpuregs[10][26] ;
 wire \cpuregs[10][27] ;
 wire \cpuregs[10][28] ;
 wire \cpuregs[10][29] ;
 wire \cpuregs[10][2] ;
 wire \cpuregs[10][30] ;
 wire \cpuregs[10][31] ;
 wire \cpuregs[10][3] ;
 wire \cpuregs[10][4] ;
 wire \cpuregs[10][5] ;
 wire \cpuregs[10][6] ;
 wire \cpuregs[10][7] ;
 wire \cpuregs[10][8] ;
 wire \cpuregs[10][9] ;
 wire \cpuregs[11][0] ;
 wire \cpuregs[11][10] ;
 wire \cpuregs[11][11] ;
 wire \cpuregs[11][12] ;
 wire \cpuregs[11][13] ;
 wire \cpuregs[11][14] ;
 wire \cpuregs[11][15] ;
 wire \cpuregs[11][16] ;
 wire \cpuregs[11][17] ;
 wire \cpuregs[11][18] ;
 wire \cpuregs[11][19] ;
 wire \cpuregs[11][1] ;
 wire \cpuregs[11][20] ;
 wire \cpuregs[11][21] ;
 wire \cpuregs[11][22] ;
 wire \cpuregs[11][23] ;
 wire \cpuregs[11][24] ;
 wire \cpuregs[11][25] ;
 wire \cpuregs[11][26] ;
 wire \cpuregs[11][27] ;
 wire \cpuregs[11][28] ;
 wire \cpuregs[11][29] ;
 wire \cpuregs[11][2] ;
 wire \cpuregs[11][30] ;
 wire \cpuregs[11][31] ;
 wire \cpuregs[11][3] ;
 wire \cpuregs[11][4] ;
 wire \cpuregs[11][5] ;
 wire \cpuregs[11][6] ;
 wire \cpuregs[11][7] ;
 wire \cpuregs[11][8] ;
 wire \cpuregs[11][9] ;
 wire \cpuregs[12][0] ;
 wire \cpuregs[12][10] ;
 wire \cpuregs[12][11] ;
 wire \cpuregs[12][12] ;
 wire \cpuregs[12][13] ;
 wire \cpuregs[12][14] ;
 wire \cpuregs[12][15] ;
 wire \cpuregs[12][16] ;
 wire \cpuregs[12][17] ;
 wire \cpuregs[12][18] ;
 wire \cpuregs[12][19] ;
 wire \cpuregs[12][1] ;
 wire \cpuregs[12][20] ;
 wire \cpuregs[12][21] ;
 wire \cpuregs[12][22] ;
 wire \cpuregs[12][23] ;
 wire \cpuregs[12][24] ;
 wire \cpuregs[12][25] ;
 wire \cpuregs[12][26] ;
 wire \cpuregs[12][27] ;
 wire \cpuregs[12][28] ;
 wire \cpuregs[12][29] ;
 wire \cpuregs[12][2] ;
 wire \cpuregs[12][30] ;
 wire \cpuregs[12][31] ;
 wire \cpuregs[12][3] ;
 wire \cpuregs[12][4] ;
 wire \cpuregs[12][5] ;
 wire \cpuregs[12][6] ;
 wire \cpuregs[12][7] ;
 wire \cpuregs[12][8] ;
 wire \cpuregs[12][9] ;
 wire \cpuregs[13][0] ;
 wire \cpuregs[13][10] ;
 wire \cpuregs[13][11] ;
 wire \cpuregs[13][12] ;
 wire \cpuregs[13][13] ;
 wire \cpuregs[13][14] ;
 wire \cpuregs[13][15] ;
 wire \cpuregs[13][16] ;
 wire \cpuregs[13][17] ;
 wire \cpuregs[13][18] ;
 wire \cpuregs[13][19] ;
 wire \cpuregs[13][1] ;
 wire \cpuregs[13][20] ;
 wire \cpuregs[13][21] ;
 wire \cpuregs[13][22] ;
 wire \cpuregs[13][23] ;
 wire \cpuregs[13][24] ;
 wire \cpuregs[13][25] ;
 wire \cpuregs[13][26] ;
 wire \cpuregs[13][27] ;
 wire \cpuregs[13][28] ;
 wire \cpuregs[13][29] ;
 wire \cpuregs[13][2] ;
 wire \cpuregs[13][30] ;
 wire \cpuregs[13][31] ;
 wire \cpuregs[13][3] ;
 wire \cpuregs[13][4] ;
 wire \cpuregs[13][5] ;
 wire \cpuregs[13][6] ;
 wire \cpuregs[13][7] ;
 wire \cpuregs[13][8] ;
 wire \cpuregs[13][9] ;
 wire \cpuregs[14][0] ;
 wire \cpuregs[14][10] ;
 wire \cpuregs[14][11] ;
 wire \cpuregs[14][12] ;
 wire \cpuregs[14][13] ;
 wire \cpuregs[14][14] ;
 wire \cpuregs[14][15] ;
 wire \cpuregs[14][16] ;
 wire \cpuregs[14][17] ;
 wire \cpuregs[14][18] ;
 wire \cpuregs[14][19] ;
 wire \cpuregs[14][1] ;
 wire \cpuregs[14][20] ;
 wire \cpuregs[14][21] ;
 wire \cpuregs[14][22] ;
 wire \cpuregs[14][23] ;
 wire \cpuregs[14][24] ;
 wire \cpuregs[14][25] ;
 wire \cpuregs[14][26] ;
 wire \cpuregs[14][27] ;
 wire \cpuregs[14][28] ;
 wire \cpuregs[14][29] ;
 wire \cpuregs[14][2] ;
 wire \cpuregs[14][30] ;
 wire \cpuregs[14][31] ;
 wire \cpuregs[14][3] ;
 wire \cpuregs[14][4] ;
 wire \cpuregs[14][5] ;
 wire \cpuregs[14][6] ;
 wire \cpuregs[14][7] ;
 wire \cpuregs[14][8] ;
 wire \cpuregs[14][9] ;
 wire \cpuregs[15][0] ;
 wire \cpuregs[15][10] ;
 wire \cpuregs[15][11] ;
 wire \cpuregs[15][12] ;
 wire \cpuregs[15][13] ;
 wire \cpuregs[15][14] ;
 wire \cpuregs[15][15] ;
 wire \cpuregs[15][16] ;
 wire \cpuregs[15][17] ;
 wire \cpuregs[15][18] ;
 wire \cpuregs[15][19] ;
 wire \cpuregs[15][1] ;
 wire \cpuregs[15][20] ;
 wire \cpuregs[15][21] ;
 wire \cpuregs[15][22] ;
 wire \cpuregs[15][23] ;
 wire \cpuregs[15][24] ;
 wire \cpuregs[15][25] ;
 wire \cpuregs[15][26] ;
 wire \cpuregs[15][27] ;
 wire \cpuregs[15][28] ;
 wire \cpuregs[15][29] ;
 wire \cpuregs[15][2] ;
 wire \cpuregs[15][30] ;
 wire \cpuregs[15][31] ;
 wire \cpuregs[15][3] ;
 wire \cpuregs[15][4] ;
 wire \cpuregs[15][5] ;
 wire \cpuregs[15][6] ;
 wire \cpuregs[15][7] ;
 wire \cpuregs[15][8] ;
 wire \cpuregs[15][9] ;
 wire \cpuregs[16][0] ;
 wire \cpuregs[16][10] ;
 wire \cpuregs[16][11] ;
 wire \cpuregs[16][12] ;
 wire \cpuregs[16][13] ;
 wire \cpuregs[16][14] ;
 wire \cpuregs[16][15] ;
 wire \cpuregs[16][16] ;
 wire \cpuregs[16][17] ;
 wire \cpuregs[16][18] ;
 wire \cpuregs[16][19] ;
 wire \cpuregs[16][1] ;
 wire \cpuregs[16][20] ;
 wire \cpuregs[16][21] ;
 wire \cpuregs[16][22] ;
 wire \cpuregs[16][23] ;
 wire \cpuregs[16][24] ;
 wire \cpuregs[16][25] ;
 wire \cpuregs[16][26] ;
 wire \cpuregs[16][27] ;
 wire \cpuregs[16][28] ;
 wire \cpuregs[16][29] ;
 wire \cpuregs[16][2] ;
 wire \cpuregs[16][30] ;
 wire \cpuregs[16][31] ;
 wire \cpuregs[16][3] ;
 wire \cpuregs[16][4] ;
 wire \cpuregs[16][5] ;
 wire \cpuregs[16][6] ;
 wire \cpuregs[16][7] ;
 wire \cpuregs[16][8] ;
 wire \cpuregs[16][9] ;
 wire \cpuregs[17][0] ;
 wire \cpuregs[17][10] ;
 wire \cpuregs[17][11] ;
 wire \cpuregs[17][12] ;
 wire \cpuregs[17][13] ;
 wire \cpuregs[17][14] ;
 wire \cpuregs[17][15] ;
 wire \cpuregs[17][16] ;
 wire \cpuregs[17][17] ;
 wire \cpuregs[17][18] ;
 wire \cpuregs[17][19] ;
 wire \cpuregs[17][1] ;
 wire \cpuregs[17][20] ;
 wire \cpuregs[17][21] ;
 wire \cpuregs[17][22] ;
 wire \cpuregs[17][23] ;
 wire \cpuregs[17][24] ;
 wire \cpuregs[17][25] ;
 wire \cpuregs[17][26] ;
 wire \cpuregs[17][27] ;
 wire \cpuregs[17][28] ;
 wire \cpuregs[17][29] ;
 wire \cpuregs[17][2] ;
 wire \cpuregs[17][30] ;
 wire \cpuregs[17][31] ;
 wire \cpuregs[17][3] ;
 wire \cpuregs[17][4] ;
 wire \cpuregs[17][5] ;
 wire \cpuregs[17][6] ;
 wire \cpuregs[17][7] ;
 wire \cpuregs[17][8] ;
 wire \cpuregs[17][9] ;
 wire \cpuregs[18][0] ;
 wire \cpuregs[18][10] ;
 wire \cpuregs[18][11] ;
 wire \cpuregs[18][12] ;
 wire \cpuregs[18][13] ;
 wire \cpuregs[18][14] ;
 wire \cpuregs[18][15] ;
 wire \cpuregs[18][16] ;
 wire \cpuregs[18][17] ;
 wire \cpuregs[18][18] ;
 wire \cpuregs[18][19] ;
 wire \cpuregs[18][1] ;
 wire \cpuregs[18][20] ;
 wire \cpuregs[18][21] ;
 wire \cpuregs[18][22] ;
 wire \cpuregs[18][23] ;
 wire \cpuregs[18][24] ;
 wire \cpuregs[18][25] ;
 wire \cpuregs[18][26] ;
 wire \cpuregs[18][27] ;
 wire \cpuregs[18][28] ;
 wire \cpuregs[18][29] ;
 wire \cpuregs[18][2] ;
 wire \cpuregs[18][30] ;
 wire \cpuregs[18][31] ;
 wire \cpuregs[18][3] ;
 wire \cpuregs[18][4] ;
 wire \cpuregs[18][5] ;
 wire \cpuregs[18][6] ;
 wire \cpuregs[18][7] ;
 wire \cpuregs[18][8] ;
 wire \cpuregs[18][9] ;
 wire \cpuregs[19][0] ;
 wire \cpuregs[19][10] ;
 wire \cpuregs[19][11] ;
 wire \cpuregs[19][12] ;
 wire \cpuregs[19][13] ;
 wire \cpuregs[19][14] ;
 wire \cpuregs[19][15] ;
 wire \cpuregs[19][16] ;
 wire \cpuregs[19][17] ;
 wire \cpuregs[19][18] ;
 wire \cpuregs[19][19] ;
 wire \cpuregs[19][1] ;
 wire \cpuregs[19][20] ;
 wire \cpuregs[19][21] ;
 wire \cpuregs[19][22] ;
 wire \cpuregs[19][23] ;
 wire \cpuregs[19][24] ;
 wire \cpuregs[19][25] ;
 wire \cpuregs[19][26] ;
 wire \cpuregs[19][27] ;
 wire \cpuregs[19][28] ;
 wire \cpuregs[19][29] ;
 wire \cpuregs[19][2] ;
 wire \cpuregs[19][30] ;
 wire \cpuregs[19][31] ;
 wire \cpuregs[19][3] ;
 wire \cpuregs[19][4] ;
 wire \cpuregs[19][5] ;
 wire \cpuregs[19][6] ;
 wire \cpuregs[19][7] ;
 wire \cpuregs[19][8] ;
 wire \cpuregs[19][9] ;
 wire \cpuregs[1][0] ;
 wire \cpuregs[1][10] ;
 wire \cpuregs[1][11] ;
 wire \cpuregs[1][12] ;
 wire \cpuregs[1][13] ;
 wire \cpuregs[1][14] ;
 wire \cpuregs[1][15] ;
 wire \cpuregs[1][16] ;
 wire \cpuregs[1][17] ;
 wire \cpuregs[1][18] ;
 wire \cpuregs[1][19] ;
 wire \cpuregs[1][1] ;
 wire \cpuregs[1][20] ;
 wire \cpuregs[1][21] ;
 wire \cpuregs[1][22] ;
 wire \cpuregs[1][23] ;
 wire \cpuregs[1][24] ;
 wire \cpuregs[1][25] ;
 wire \cpuregs[1][26] ;
 wire \cpuregs[1][27] ;
 wire \cpuregs[1][28] ;
 wire \cpuregs[1][29] ;
 wire \cpuregs[1][2] ;
 wire \cpuregs[1][30] ;
 wire \cpuregs[1][31] ;
 wire \cpuregs[1][3] ;
 wire \cpuregs[1][4] ;
 wire \cpuregs[1][5] ;
 wire \cpuregs[1][6] ;
 wire \cpuregs[1][7] ;
 wire \cpuregs[1][8] ;
 wire \cpuregs[1][9] ;
 wire \cpuregs[20][0] ;
 wire \cpuregs[20][10] ;
 wire \cpuregs[20][11] ;
 wire \cpuregs[20][12] ;
 wire \cpuregs[20][13] ;
 wire \cpuregs[20][14] ;
 wire \cpuregs[20][15] ;
 wire \cpuregs[20][16] ;
 wire \cpuregs[20][17] ;
 wire \cpuregs[20][18] ;
 wire \cpuregs[20][19] ;
 wire \cpuregs[20][1] ;
 wire \cpuregs[20][20] ;
 wire \cpuregs[20][21] ;
 wire \cpuregs[20][22] ;
 wire \cpuregs[20][23] ;
 wire \cpuregs[20][24] ;
 wire \cpuregs[20][25] ;
 wire \cpuregs[20][26] ;
 wire \cpuregs[20][27] ;
 wire \cpuregs[20][28] ;
 wire \cpuregs[20][29] ;
 wire \cpuregs[20][2] ;
 wire \cpuregs[20][30] ;
 wire \cpuregs[20][31] ;
 wire \cpuregs[20][3] ;
 wire \cpuregs[20][4] ;
 wire \cpuregs[20][5] ;
 wire \cpuregs[20][6] ;
 wire \cpuregs[20][7] ;
 wire \cpuregs[20][8] ;
 wire \cpuregs[20][9] ;
 wire \cpuregs[21][0] ;
 wire \cpuregs[21][10] ;
 wire \cpuregs[21][11] ;
 wire \cpuregs[21][12] ;
 wire \cpuregs[21][13] ;
 wire \cpuregs[21][14] ;
 wire \cpuregs[21][15] ;
 wire \cpuregs[21][16] ;
 wire \cpuregs[21][17] ;
 wire \cpuregs[21][18] ;
 wire \cpuregs[21][19] ;
 wire \cpuregs[21][1] ;
 wire \cpuregs[21][20] ;
 wire \cpuregs[21][21] ;
 wire \cpuregs[21][22] ;
 wire \cpuregs[21][23] ;
 wire \cpuregs[21][24] ;
 wire \cpuregs[21][25] ;
 wire \cpuregs[21][26] ;
 wire \cpuregs[21][27] ;
 wire \cpuregs[21][28] ;
 wire \cpuregs[21][29] ;
 wire \cpuregs[21][2] ;
 wire \cpuregs[21][30] ;
 wire \cpuregs[21][31] ;
 wire \cpuregs[21][3] ;
 wire \cpuregs[21][4] ;
 wire \cpuregs[21][5] ;
 wire \cpuregs[21][6] ;
 wire \cpuregs[21][7] ;
 wire \cpuregs[21][8] ;
 wire \cpuregs[21][9] ;
 wire \cpuregs[22][0] ;
 wire \cpuregs[22][10] ;
 wire \cpuregs[22][11] ;
 wire \cpuregs[22][12] ;
 wire \cpuregs[22][13] ;
 wire \cpuregs[22][14] ;
 wire \cpuregs[22][15] ;
 wire \cpuregs[22][16] ;
 wire \cpuregs[22][17] ;
 wire \cpuregs[22][18] ;
 wire \cpuregs[22][19] ;
 wire \cpuregs[22][1] ;
 wire \cpuregs[22][20] ;
 wire \cpuregs[22][21] ;
 wire \cpuregs[22][22] ;
 wire \cpuregs[22][23] ;
 wire \cpuregs[22][24] ;
 wire \cpuregs[22][25] ;
 wire \cpuregs[22][26] ;
 wire \cpuregs[22][27] ;
 wire \cpuregs[22][28] ;
 wire \cpuregs[22][29] ;
 wire \cpuregs[22][2] ;
 wire \cpuregs[22][30] ;
 wire \cpuregs[22][31] ;
 wire \cpuregs[22][3] ;
 wire \cpuregs[22][4] ;
 wire \cpuregs[22][5] ;
 wire \cpuregs[22][6] ;
 wire \cpuregs[22][7] ;
 wire \cpuregs[22][8] ;
 wire \cpuregs[22][9] ;
 wire \cpuregs[23][0] ;
 wire \cpuregs[23][10] ;
 wire \cpuregs[23][11] ;
 wire \cpuregs[23][12] ;
 wire \cpuregs[23][13] ;
 wire \cpuregs[23][14] ;
 wire \cpuregs[23][15] ;
 wire \cpuregs[23][16] ;
 wire \cpuregs[23][17] ;
 wire \cpuregs[23][18] ;
 wire \cpuregs[23][19] ;
 wire \cpuregs[23][1] ;
 wire \cpuregs[23][20] ;
 wire \cpuregs[23][21] ;
 wire \cpuregs[23][22] ;
 wire \cpuregs[23][23] ;
 wire \cpuregs[23][24] ;
 wire \cpuregs[23][25] ;
 wire \cpuregs[23][26] ;
 wire \cpuregs[23][27] ;
 wire \cpuregs[23][28] ;
 wire \cpuregs[23][29] ;
 wire \cpuregs[23][2] ;
 wire \cpuregs[23][30] ;
 wire \cpuregs[23][31] ;
 wire \cpuregs[23][3] ;
 wire \cpuregs[23][4] ;
 wire \cpuregs[23][5] ;
 wire \cpuregs[23][6] ;
 wire \cpuregs[23][7] ;
 wire \cpuregs[23][8] ;
 wire \cpuregs[23][9] ;
 wire \cpuregs[24][0] ;
 wire \cpuregs[24][10] ;
 wire \cpuregs[24][11] ;
 wire \cpuregs[24][12] ;
 wire \cpuregs[24][13] ;
 wire \cpuregs[24][14] ;
 wire \cpuregs[24][15] ;
 wire \cpuregs[24][16] ;
 wire \cpuregs[24][17] ;
 wire \cpuregs[24][18] ;
 wire \cpuregs[24][19] ;
 wire \cpuregs[24][1] ;
 wire \cpuregs[24][20] ;
 wire \cpuregs[24][21] ;
 wire \cpuregs[24][22] ;
 wire \cpuregs[24][23] ;
 wire \cpuregs[24][24] ;
 wire \cpuregs[24][25] ;
 wire \cpuregs[24][26] ;
 wire \cpuregs[24][27] ;
 wire \cpuregs[24][28] ;
 wire \cpuregs[24][29] ;
 wire \cpuregs[24][2] ;
 wire \cpuregs[24][30] ;
 wire \cpuregs[24][31] ;
 wire \cpuregs[24][3] ;
 wire \cpuregs[24][4] ;
 wire \cpuregs[24][5] ;
 wire \cpuregs[24][6] ;
 wire \cpuregs[24][7] ;
 wire \cpuregs[24][8] ;
 wire \cpuregs[24][9] ;
 wire \cpuregs[25][0] ;
 wire \cpuregs[25][10] ;
 wire \cpuregs[25][11] ;
 wire \cpuregs[25][12] ;
 wire \cpuregs[25][13] ;
 wire \cpuregs[25][14] ;
 wire \cpuregs[25][15] ;
 wire \cpuregs[25][16] ;
 wire \cpuregs[25][17] ;
 wire \cpuregs[25][18] ;
 wire \cpuregs[25][19] ;
 wire \cpuregs[25][1] ;
 wire \cpuregs[25][20] ;
 wire \cpuregs[25][21] ;
 wire \cpuregs[25][22] ;
 wire \cpuregs[25][23] ;
 wire \cpuregs[25][24] ;
 wire \cpuregs[25][25] ;
 wire \cpuregs[25][26] ;
 wire \cpuregs[25][27] ;
 wire \cpuregs[25][28] ;
 wire \cpuregs[25][29] ;
 wire \cpuregs[25][2] ;
 wire \cpuregs[25][30] ;
 wire \cpuregs[25][31] ;
 wire \cpuregs[25][3] ;
 wire \cpuregs[25][4] ;
 wire \cpuregs[25][5] ;
 wire \cpuregs[25][6] ;
 wire \cpuregs[25][7] ;
 wire \cpuregs[25][8] ;
 wire \cpuregs[25][9] ;
 wire \cpuregs[26][0] ;
 wire \cpuregs[26][10] ;
 wire \cpuregs[26][11] ;
 wire \cpuregs[26][12] ;
 wire \cpuregs[26][13] ;
 wire \cpuregs[26][14] ;
 wire \cpuregs[26][15] ;
 wire \cpuregs[26][16] ;
 wire \cpuregs[26][17] ;
 wire \cpuregs[26][18] ;
 wire \cpuregs[26][19] ;
 wire \cpuregs[26][1] ;
 wire \cpuregs[26][20] ;
 wire \cpuregs[26][21] ;
 wire \cpuregs[26][22] ;
 wire \cpuregs[26][23] ;
 wire \cpuregs[26][24] ;
 wire \cpuregs[26][25] ;
 wire \cpuregs[26][26] ;
 wire \cpuregs[26][27] ;
 wire \cpuregs[26][28] ;
 wire \cpuregs[26][29] ;
 wire \cpuregs[26][2] ;
 wire \cpuregs[26][30] ;
 wire \cpuregs[26][31] ;
 wire \cpuregs[26][3] ;
 wire \cpuregs[26][4] ;
 wire \cpuregs[26][5] ;
 wire \cpuregs[26][6] ;
 wire \cpuregs[26][7] ;
 wire \cpuregs[26][8] ;
 wire \cpuregs[26][9] ;
 wire \cpuregs[27][0] ;
 wire \cpuregs[27][10] ;
 wire \cpuregs[27][11] ;
 wire \cpuregs[27][12] ;
 wire \cpuregs[27][13] ;
 wire \cpuregs[27][14] ;
 wire \cpuregs[27][15] ;
 wire \cpuregs[27][16] ;
 wire \cpuregs[27][17] ;
 wire \cpuregs[27][18] ;
 wire \cpuregs[27][19] ;
 wire \cpuregs[27][1] ;
 wire \cpuregs[27][20] ;
 wire \cpuregs[27][21] ;
 wire \cpuregs[27][22] ;
 wire \cpuregs[27][23] ;
 wire \cpuregs[27][24] ;
 wire \cpuregs[27][25] ;
 wire \cpuregs[27][26] ;
 wire \cpuregs[27][27] ;
 wire \cpuregs[27][28] ;
 wire \cpuregs[27][29] ;
 wire \cpuregs[27][2] ;
 wire \cpuregs[27][30] ;
 wire \cpuregs[27][31] ;
 wire \cpuregs[27][3] ;
 wire \cpuregs[27][4] ;
 wire \cpuregs[27][5] ;
 wire \cpuregs[27][6] ;
 wire \cpuregs[27][7] ;
 wire \cpuregs[27][8] ;
 wire \cpuregs[27][9] ;
 wire \cpuregs[28][0] ;
 wire \cpuregs[28][10] ;
 wire \cpuregs[28][11] ;
 wire \cpuregs[28][12] ;
 wire \cpuregs[28][13] ;
 wire \cpuregs[28][14] ;
 wire \cpuregs[28][15] ;
 wire \cpuregs[28][16] ;
 wire \cpuregs[28][17] ;
 wire \cpuregs[28][18] ;
 wire \cpuregs[28][19] ;
 wire \cpuregs[28][1] ;
 wire \cpuregs[28][20] ;
 wire \cpuregs[28][21] ;
 wire \cpuregs[28][22] ;
 wire \cpuregs[28][23] ;
 wire \cpuregs[28][24] ;
 wire \cpuregs[28][25] ;
 wire \cpuregs[28][26] ;
 wire \cpuregs[28][27] ;
 wire \cpuregs[28][28] ;
 wire \cpuregs[28][29] ;
 wire \cpuregs[28][2] ;
 wire \cpuregs[28][30] ;
 wire \cpuregs[28][31] ;
 wire \cpuregs[28][3] ;
 wire \cpuregs[28][4] ;
 wire \cpuregs[28][5] ;
 wire \cpuregs[28][6] ;
 wire \cpuregs[28][7] ;
 wire \cpuregs[28][8] ;
 wire \cpuregs[28][9] ;
 wire \cpuregs[29][0] ;
 wire \cpuregs[29][10] ;
 wire \cpuregs[29][11] ;
 wire \cpuregs[29][12] ;
 wire \cpuregs[29][13] ;
 wire \cpuregs[29][14] ;
 wire \cpuregs[29][15] ;
 wire \cpuregs[29][16] ;
 wire \cpuregs[29][17] ;
 wire \cpuregs[29][18] ;
 wire \cpuregs[29][19] ;
 wire \cpuregs[29][1] ;
 wire \cpuregs[29][20] ;
 wire \cpuregs[29][21] ;
 wire \cpuregs[29][22] ;
 wire \cpuregs[29][23] ;
 wire \cpuregs[29][24] ;
 wire \cpuregs[29][25] ;
 wire \cpuregs[29][26] ;
 wire \cpuregs[29][27] ;
 wire \cpuregs[29][28] ;
 wire \cpuregs[29][29] ;
 wire \cpuregs[29][2] ;
 wire \cpuregs[29][30] ;
 wire \cpuregs[29][31] ;
 wire \cpuregs[29][3] ;
 wire \cpuregs[29][4] ;
 wire \cpuregs[29][5] ;
 wire \cpuregs[29][6] ;
 wire \cpuregs[29][7] ;
 wire \cpuregs[29][8] ;
 wire \cpuregs[29][9] ;
 wire \cpuregs[2][0] ;
 wire \cpuregs[2][10] ;
 wire \cpuregs[2][11] ;
 wire \cpuregs[2][12] ;
 wire \cpuregs[2][13] ;
 wire \cpuregs[2][14] ;
 wire \cpuregs[2][15] ;
 wire \cpuregs[2][16] ;
 wire \cpuregs[2][17] ;
 wire \cpuregs[2][18] ;
 wire \cpuregs[2][19] ;
 wire \cpuregs[2][1] ;
 wire \cpuregs[2][20] ;
 wire \cpuregs[2][21] ;
 wire \cpuregs[2][22] ;
 wire \cpuregs[2][23] ;
 wire \cpuregs[2][24] ;
 wire \cpuregs[2][25] ;
 wire \cpuregs[2][26] ;
 wire \cpuregs[2][27] ;
 wire \cpuregs[2][28] ;
 wire \cpuregs[2][29] ;
 wire \cpuregs[2][2] ;
 wire \cpuregs[2][30] ;
 wire \cpuregs[2][31] ;
 wire \cpuregs[2][3] ;
 wire \cpuregs[2][4] ;
 wire \cpuregs[2][5] ;
 wire \cpuregs[2][6] ;
 wire \cpuregs[2][7] ;
 wire \cpuregs[2][8] ;
 wire \cpuregs[2][9] ;
 wire \cpuregs[30][0] ;
 wire \cpuregs[30][10] ;
 wire \cpuregs[30][11] ;
 wire \cpuregs[30][12] ;
 wire \cpuregs[30][13] ;
 wire \cpuregs[30][14] ;
 wire \cpuregs[30][15] ;
 wire \cpuregs[30][16] ;
 wire \cpuregs[30][17] ;
 wire \cpuregs[30][18] ;
 wire \cpuregs[30][19] ;
 wire \cpuregs[30][1] ;
 wire \cpuregs[30][20] ;
 wire \cpuregs[30][21] ;
 wire \cpuregs[30][22] ;
 wire \cpuregs[30][23] ;
 wire \cpuregs[30][24] ;
 wire \cpuregs[30][25] ;
 wire \cpuregs[30][26] ;
 wire \cpuregs[30][27] ;
 wire \cpuregs[30][28] ;
 wire \cpuregs[30][29] ;
 wire \cpuregs[30][2] ;
 wire \cpuregs[30][30] ;
 wire \cpuregs[30][31] ;
 wire \cpuregs[30][3] ;
 wire \cpuregs[30][4] ;
 wire \cpuregs[30][5] ;
 wire \cpuregs[30][6] ;
 wire \cpuregs[30][7] ;
 wire \cpuregs[30][8] ;
 wire \cpuregs[30][9] ;
 wire \cpuregs[31][0] ;
 wire \cpuregs[31][10] ;
 wire \cpuregs[31][11] ;
 wire \cpuregs[31][12] ;
 wire \cpuregs[31][13] ;
 wire \cpuregs[31][14] ;
 wire \cpuregs[31][15] ;
 wire \cpuregs[31][16] ;
 wire \cpuregs[31][17] ;
 wire \cpuregs[31][18] ;
 wire \cpuregs[31][19] ;
 wire \cpuregs[31][1] ;
 wire \cpuregs[31][20] ;
 wire \cpuregs[31][21] ;
 wire \cpuregs[31][22] ;
 wire \cpuregs[31][23] ;
 wire \cpuregs[31][24] ;
 wire \cpuregs[31][25] ;
 wire \cpuregs[31][26] ;
 wire \cpuregs[31][27] ;
 wire \cpuregs[31][28] ;
 wire \cpuregs[31][29] ;
 wire \cpuregs[31][2] ;
 wire \cpuregs[31][30] ;
 wire \cpuregs[31][31] ;
 wire \cpuregs[31][3] ;
 wire \cpuregs[31][4] ;
 wire \cpuregs[31][5] ;
 wire \cpuregs[31][6] ;
 wire \cpuregs[31][7] ;
 wire \cpuregs[31][8] ;
 wire \cpuregs[31][9] ;
 wire \cpuregs[3][0] ;
 wire \cpuregs[3][10] ;
 wire \cpuregs[3][11] ;
 wire \cpuregs[3][12] ;
 wire \cpuregs[3][13] ;
 wire \cpuregs[3][14] ;
 wire \cpuregs[3][15] ;
 wire \cpuregs[3][16] ;
 wire \cpuregs[3][17] ;
 wire \cpuregs[3][18] ;
 wire \cpuregs[3][19] ;
 wire \cpuregs[3][1] ;
 wire \cpuregs[3][20] ;
 wire \cpuregs[3][21] ;
 wire \cpuregs[3][22] ;
 wire \cpuregs[3][23] ;
 wire \cpuregs[3][24] ;
 wire \cpuregs[3][25] ;
 wire \cpuregs[3][26] ;
 wire \cpuregs[3][27] ;
 wire \cpuregs[3][28] ;
 wire \cpuregs[3][29] ;
 wire \cpuregs[3][2] ;
 wire \cpuregs[3][30] ;
 wire \cpuregs[3][31] ;
 wire \cpuregs[3][3] ;
 wire \cpuregs[3][4] ;
 wire \cpuregs[3][5] ;
 wire \cpuregs[3][6] ;
 wire \cpuregs[3][7] ;
 wire \cpuregs[3][8] ;
 wire \cpuregs[3][9] ;
 wire \cpuregs[4][0] ;
 wire \cpuregs[4][10] ;
 wire \cpuregs[4][11] ;
 wire \cpuregs[4][12] ;
 wire \cpuregs[4][13] ;
 wire \cpuregs[4][14] ;
 wire \cpuregs[4][15] ;
 wire \cpuregs[4][16] ;
 wire \cpuregs[4][17] ;
 wire \cpuregs[4][18] ;
 wire \cpuregs[4][19] ;
 wire \cpuregs[4][1] ;
 wire \cpuregs[4][20] ;
 wire \cpuregs[4][21] ;
 wire \cpuregs[4][22] ;
 wire \cpuregs[4][23] ;
 wire \cpuregs[4][24] ;
 wire \cpuregs[4][25] ;
 wire \cpuregs[4][26] ;
 wire \cpuregs[4][27] ;
 wire \cpuregs[4][28] ;
 wire \cpuregs[4][29] ;
 wire \cpuregs[4][2] ;
 wire \cpuregs[4][30] ;
 wire \cpuregs[4][31] ;
 wire \cpuregs[4][3] ;
 wire \cpuregs[4][4] ;
 wire \cpuregs[4][5] ;
 wire \cpuregs[4][6] ;
 wire \cpuregs[4][7] ;
 wire \cpuregs[4][8] ;
 wire \cpuregs[4][9] ;
 wire \cpuregs[5][0] ;
 wire \cpuregs[5][10] ;
 wire \cpuregs[5][11] ;
 wire \cpuregs[5][12] ;
 wire \cpuregs[5][13] ;
 wire \cpuregs[5][14] ;
 wire \cpuregs[5][15] ;
 wire \cpuregs[5][16] ;
 wire \cpuregs[5][17] ;
 wire \cpuregs[5][18] ;
 wire \cpuregs[5][19] ;
 wire \cpuregs[5][1] ;
 wire \cpuregs[5][20] ;
 wire \cpuregs[5][21] ;
 wire \cpuregs[5][22] ;
 wire \cpuregs[5][23] ;
 wire \cpuregs[5][24] ;
 wire \cpuregs[5][25] ;
 wire \cpuregs[5][26] ;
 wire \cpuregs[5][27] ;
 wire \cpuregs[5][28] ;
 wire \cpuregs[5][29] ;
 wire \cpuregs[5][2] ;
 wire \cpuregs[5][30] ;
 wire \cpuregs[5][31] ;
 wire \cpuregs[5][3] ;
 wire \cpuregs[5][4] ;
 wire \cpuregs[5][5] ;
 wire \cpuregs[5][6] ;
 wire \cpuregs[5][7] ;
 wire \cpuregs[5][8] ;
 wire \cpuregs[5][9] ;
 wire \cpuregs[6][0] ;
 wire \cpuregs[6][10] ;
 wire \cpuregs[6][11] ;
 wire \cpuregs[6][12] ;
 wire \cpuregs[6][13] ;
 wire \cpuregs[6][14] ;
 wire \cpuregs[6][15] ;
 wire \cpuregs[6][16] ;
 wire \cpuregs[6][17] ;
 wire \cpuregs[6][18] ;
 wire \cpuregs[6][19] ;
 wire \cpuregs[6][1] ;
 wire \cpuregs[6][20] ;
 wire \cpuregs[6][21] ;
 wire \cpuregs[6][22] ;
 wire \cpuregs[6][23] ;
 wire \cpuregs[6][24] ;
 wire \cpuregs[6][25] ;
 wire \cpuregs[6][26] ;
 wire \cpuregs[6][27] ;
 wire \cpuregs[6][28] ;
 wire \cpuregs[6][29] ;
 wire \cpuregs[6][2] ;
 wire \cpuregs[6][30] ;
 wire \cpuregs[6][31] ;
 wire \cpuregs[6][3] ;
 wire \cpuregs[6][4] ;
 wire \cpuregs[6][5] ;
 wire \cpuregs[6][6] ;
 wire \cpuregs[6][7] ;
 wire \cpuregs[6][8] ;
 wire \cpuregs[6][9] ;
 wire \cpuregs[7][0] ;
 wire \cpuregs[7][10] ;
 wire \cpuregs[7][11] ;
 wire \cpuregs[7][12] ;
 wire \cpuregs[7][13] ;
 wire \cpuregs[7][14] ;
 wire \cpuregs[7][15] ;
 wire \cpuregs[7][16] ;
 wire \cpuregs[7][17] ;
 wire \cpuregs[7][18] ;
 wire \cpuregs[7][19] ;
 wire \cpuregs[7][1] ;
 wire \cpuregs[7][20] ;
 wire \cpuregs[7][21] ;
 wire \cpuregs[7][22] ;
 wire \cpuregs[7][23] ;
 wire \cpuregs[7][24] ;
 wire \cpuregs[7][25] ;
 wire \cpuregs[7][26] ;
 wire \cpuregs[7][27] ;
 wire \cpuregs[7][28] ;
 wire \cpuregs[7][29] ;
 wire \cpuregs[7][2] ;
 wire \cpuregs[7][30] ;
 wire \cpuregs[7][31] ;
 wire \cpuregs[7][3] ;
 wire \cpuregs[7][4] ;
 wire \cpuregs[7][5] ;
 wire \cpuregs[7][6] ;
 wire \cpuregs[7][7] ;
 wire \cpuregs[7][8] ;
 wire \cpuregs[7][9] ;
 wire \cpuregs[8][0] ;
 wire \cpuregs[8][10] ;
 wire \cpuregs[8][11] ;
 wire \cpuregs[8][12] ;
 wire \cpuregs[8][13] ;
 wire \cpuregs[8][14] ;
 wire \cpuregs[8][15] ;
 wire \cpuregs[8][16] ;
 wire \cpuregs[8][17] ;
 wire \cpuregs[8][18] ;
 wire \cpuregs[8][19] ;
 wire \cpuregs[8][1] ;
 wire \cpuregs[8][20] ;
 wire \cpuregs[8][21] ;
 wire \cpuregs[8][22] ;
 wire \cpuregs[8][23] ;
 wire \cpuregs[8][24] ;
 wire \cpuregs[8][25] ;
 wire \cpuregs[8][26] ;
 wire \cpuregs[8][27] ;
 wire \cpuregs[8][28] ;
 wire \cpuregs[8][29] ;
 wire \cpuregs[8][2] ;
 wire \cpuregs[8][30] ;
 wire \cpuregs[8][31] ;
 wire \cpuregs[8][3] ;
 wire \cpuregs[8][4] ;
 wire \cpuregs[8][5] ;
 wire \cpuregs[8][6] ;
 wire \cpuregs[8][7] ;
 wire \cpuregs[8][8] ;
 wire \cpuregs[8][9] ;
 wire \cpuregs[9][0] ;
 wire \cpuregs[9][10] ;
 wire \cpuregs[9][11] ;
 wire \cpuregs[9][12] ;
 wire \cpuregs[9][13] ;
 wire \cpuregs[9][14] ;
 wire \cpuregs[9][15] ;
 wire \cpuregs[9][16] ;
 wire \cpuregs[9][17] ;
 wire \cpuregs[9][18] ;
 wire \cpuregs[9][19] ;
 wire \cpuregs[9][1] ;
 wire \cpuregs[9][20] ;
 wire \cpuregs[9][21] ;
 wire \cpuregs[9][22] ;
 wire \cpuregs[9][23] ;
 wire \cpuregs[9][24] ;
 wire \cpuregs[9][25] ;
 wire \cpuregs[9][26] ;
 wire \cpuregs[9][27] ;
 wire \cpuregs[9][28] ;
 wire \cpuregs[9][29] ;
 wire \cpuregs[9][2] ;
 wire \cpuregs[9][30] ;
 wire \cpuregs[9][31] ;
 wire \cpuregs[9][3] ;
 wire \cpuregs[9][4] ;
 wire \cpuregs[9][5] ;
 wire \cpuregs[9][6] ;
 wire \cpuregs[9][7] ;
 wire \cpuregs[9][8] ;
 wire \cpuregs[9][9] ;
 wire \decoded_imm[0] ;
 wire \decoded_imm[10] ;
 wire \decoded_imm[11] ;
 wire \decoded_imm[12] ;
 wire \decoded_imm[13] ;
 wire \decoded_imm[14] ;
 wire \decoded_imm[15] ;
 wire \decoded_imm[16] ;
 wire \decoded_imm[17] ;
 wire \decoded_imm[18] ;
 wire \decoded_imm[19] ;
 wire \decoded_imm[1] ;
 wire \decoded_imm[20] ;
 wire \decoded_imm[21] ;
 wire \decoded_imm[22] ;
 wire \decoded_imm[23] ;
 wire \decoded_imm[24] ;
 wire \decoded_imm[25] ;
 wire \decoded_imm[26] ;
 wire \decoded_imm[27] ;
 wire \decoded_imm[28] ;
 wire \decoded_imm[29] ;
 wire \decoded_imm[2] ;
 wire \decoded_imm[30] ;
 wire \decoded_imm[31] ;
 wire \decoded_imm[3] ;
 wire \decoded_imm[4] ;
 wire \decoded_imm[5] ;
 wire \decoded_imm[6] ;
 wire \decoded_imm[7] ;
 wire \decoded_imm[8] ;
 wire \decoded_imm[9] ;
 wire \decoded_imm_j[10] ;
 wire \decoded_imm_j[11] ;
 wire \decoded_imm_j[12] ;
 wire \decoded_imm_j[13] ;
 wire \decoded_imm_j[14] ;
 wire \decoded_imm_j[15] ;
 wire \decoded_imm_j[16] ;
 wire \decoded_imm_j[17] ;
 wire \decoded_imm_j[18] ;
 wire \decoded_imm_j[19] ;
 wire \decoded_imm_j[1] ;
 wire \decoded_imm_j[20] ;
 wire \decoded_imm_j[2] ;
 wire \decoded_imm_j[3] ;
 wire \decoded_imm_j[4] ;
 wire \decoded_imm_j[5] ;
 wire \decoded_imm_j[6] ;
 wire \decoded_imm_j[7] ;
 wire \decoded_imm_j[8] ;
 wire \decoded_imm_j[9] ;
 wire \decoded_rd[0] ;
 wire \decoded_rd[1] ;
 wire \decoded_rd[2] ;
 wire \decoded_rd[3] ;
 wire \decoded_rd[4] ;
 wire decoder_pseudo_trigger;
 wire decoder_trigger;
 wire net1243;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1244;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1245;
 wire net1273;
 wire net1274;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire \genblk1.genblk1.pcpi_mul.instr_any_mul ;
 wire \genblk1.genblk1.pcpi_mul.instr_mul ;
 wire \genblk1.genblk1.pcpi_mul.instr_mulh ;
 wire \genblk1.genblk1.pcpi_mul.instr_mulhsu ;
 wire \genblk1.genblk1.pcpi_mul.instr_mulhu ;
 wire \genblk1.genblk1.pcpi_mul.mul_counter[0] ;
 wire \genblk1.genblk1.pcpi_mul.mul_counter[1] ;
 wire \genblk1.genblk1.pcpi_mul.mul_counter[2] ;
 wire \genblk1.genblk1.pcpi_mul.mul_counter[3] ;
 wire \genblk1.genblk1.pcpi_mul.mul_counter[4] ;
 wire \genblk1.genblk1.pcpi_mul.mul_counter[5] ;
 wire \genblk1.genblk1.pcpi_mul.mul_counter[6] ;
 wire \genblk1.genblk1.pcpi_mul.mul_finish ;
 wire \genblk1.genblk1.pcpi_mul.mul_waiting ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[0] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[10] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[11] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[12] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[13] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[14] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[15] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[16] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[17] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[18] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[19] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[1] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[20] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[21] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[22] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[23] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[24] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[25] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[26] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[27] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[28] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[29] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[2] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[30] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[31] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[32] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[33] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[34] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[35] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[36] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[37] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[38] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[39] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[3] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[40] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[41] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[42] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[43] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[44] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[45] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[46] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[47] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[48] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[49] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[4] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[50] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[51] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[52] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[53] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[54] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[55] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[56] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[57] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[58] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[59] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[5] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[60] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[61] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[62] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[6] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[7] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[8] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs1[9] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[10] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[11] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[12] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[13] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[14] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[15] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[16] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[17] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[18] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[19] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[1] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[20] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[21] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[22] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[23] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[24] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[25] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[26] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[27] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[28] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[29] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[2] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[30] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[31] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[32] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[33] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[34] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[35] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[36] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[37] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[38] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[39] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[3] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[40] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[41] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[42] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[43] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[44] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[45] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[46] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[47] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[48] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[49] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[4] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[50] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[51] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[52] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[53] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[54] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[55] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[56] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[57] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[58] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[59] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[5] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[60] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[61] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[62] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[63] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[6] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[7] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[8] ;
 wire \genblk1.genblk1.pcpi_mul.next_rs2[9] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[0] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[10] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[11] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[12] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[13] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[14] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[15] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[16] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[17] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[18] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[19] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[1] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[20] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[21] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[22] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[23] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[24] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[25] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[26] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[27] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[28] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[29] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[2] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[30] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[31] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[3] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[4] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[5] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[6] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[7] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[8] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_rd[9] ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_ready ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_wait ;
 wire \genblk1.genblk1.pcpi_mul.pcpi_wait_q ;
 wire \genblk1.genblk1.pcpi_mul.rd[0] ;
 wire \genblk1.genblk1.pcpi_mul.rd[10] ;
 wire \genblk1.genblk1.pcpi_mul.rd[11] ;
 wire \genblk1.genblk1.pcpi_mul.rd[12] ;
 wire \genblk1.genblk1.pcpi_mul.rd[13] ;
 wire \genblk1.genblk1.pcpi_mul.rd[14] ;
 wire \genblk1.genblk1.pcpi_mul.rd[15] ;
 wire \genblk1.genblk1.pcpi_mul.rd[16] ;
 wire \genblk1.genblk1.pcpi_mul.rd[17] ;
 wire \genblk1.genblk1.pcpi_mul.rd[18] ;
 wire \genblk1.genblk1.pcpi_mul.rd[19] ;
 wire \genblk1.genblk1.pcpi_mul.rd[1] ;
 wire \genblk1.genblk1.pcpi_mul.rd[20] ;
 wire \genblk1.genblk1.pcpi_mul.rd[21] ;
 wire \genblk1.genblk1.pcpi_mul.rd[22] ;
 wire \genblk1.genblk1.pcpi_mul.rd[23] ;
 wire \genblk1.genblk1.pcpi_mul.rd[24] ;
 wire \genblk1.genblk1.pcpi_mul.rd[25] ;
 wire \genblk1.genblk1.pcpi_mul.rd[26] ;
 wire \genblk1.genblk1.pcpi_mul.rd[27] ;
 wire \genblk1.genblk1.pcpi_mul.rd[28] ;
 wire \genblk1.genblk1.pcpi_mul.rd[29] ;
 wire \genblk1.genblk1.pcpi_mul.rd[2] ;
 wire \genblk1.genblk1.pcpi_mul.rd[30] ;
 wire \genblk1.genblk1.pcpi_mul.rd[31] ;
 wire \genblk1.genblk1.pcpi_mul.rd[32] ;
 wire \genblk1.genblk1.pcpi_mul.rd[33] ;
 wire \genblk1.genblk1.pcpi_mul.rd[34] ;
 wire \genblk1.genblk1.pcpi_mul.rd[35] ;
 wire \genblk1.genblk1.pcpi_mul.rd[36] ;
 wire \genblk1.genblk1.pcpi_mul.rd[37] ;
 wire \genblk1.genblk1.pcpi_mul.rd[38] ;
 wire \genblk1.genblk1.pcpi_mul.rd[39] ;
 wire \genblk1.genblk1.pcpi_mul.rd[3] ;
 wire \genblk1.genblk1.pcpi_mul.rd[40] ;
 wire \genblk1.genblk1.pcpi_mul.rd[41] ;
 wire \genblk1.genblk1.pcpi_mul.rd[42] ;
 wire \genblk1.genblk1.pcpi_mul.rd[43] ;
 wire \genblk1.genblk1.pcpi_mul.rd[44] ;
 wire \genblk1.genblk1.pcpi_mul.rd[45] ;
 wire \genblk1.genblk1.pcpi_mul.rd[46] ;
 wire \genblk1.genblk1.pcpi_mul.rd[47] ;
 wire \genblk1.genblk1.pcpi_mul.rd[48] ;
 wire \genblk1.genblk1.pcpi_mul.rd[49] ;
 wire \genblk1.genblk1.pcpi_mul.rd[4] ;
 wire \genblk1.genblk1.pcpi_mul.rd[50] ;
 wire \genblk1.genblk1.pcpi_mul.rd[51] ;
 wire \genblk1.genblk1.pcpi_mul.rd[52] ;
 wire \genblk1.genblk1.pcpi_mul.rd[53] ;
 wire \genblk1.genblk1.pcpi_mul.rd[54] ;
 wire \genblk1.genblk1.pcpi_mul.rd[55] ;
 wire \genblk1.genblk1.pcpi_mul.rd[56] ;
 wire \genblk1.genblk1.pcpi_mul.rd[57] ;
 wire \genblk1.genblk1.pcpi_mul.rd[58] ;
 wire \genblk1.genblk1.pcpi_mul.rd[59] ;
 wire \genblk1.genblk1.pcpi_mul.rd[5] ;
 wire \genblk1.genblk1.pcpi_mul.rd[60] ;
 wire \genblk1.genblk1.pcpi_mul.rd[61] ;
 wire \genblk1.genblk1.pcpi_mul.rd[62] ;
 wire \genblk1.genblk1.pcpi_mul.rd[63] ;
 wire \genblk1.genblk1.pcpi_mul.rd[6] ;
 wire \genblk1.genblk1.pcpi_mul.rd[7] ;
 wire \genblk1.genblk1.pcpi_mul.rd[8] ;
 wire \genblk1.genblk1.pcpi_mul.rd[9] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[12] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[16] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[20] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[24] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[28] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[32] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[36] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[40] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[44] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[48] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[4] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[52] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[56] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[60] ;
 wire \genblk1.genblk1.pcpi_mul.rdx[8] ;
 wire \genblk1.genblk1.pcpi_mul.rs1[0] ;
 wire \genblk1.genblk1.pcpi_mul.rs2[63] ;
 wire \genblk2.pcpi_div.dividend[0] ;
 wire \genblk2.pcpi_div.dividend[10] ;
 wire \genblk2.pcpi_div.dividend[11] ;
 wire \genblk2.pcpi_div.dividend[12] ;
 wire \genblk2.pcpi_div.dividend[13] ;
 wire \genblk2.pcpi_div.dividend[14] ;
 wire \genblk2.pcpi_div.dividend[15] ;
 wire \genblk2.pcpi_div.dividend[16] ;
 wire \genblk2.pcpi_div.dividend[17] ;
 wire \genblk2.pcpi_div.dividend[18] ;
 wire \genblk2.pcpi_div.dividend[19] ;
 wire \genblk2.pcpi_div.dividend[1] ;
 wire \genblk2.pcpi_div.dividend[20] ;
 wire \genblk2.pcpi_div.dividend[21] ;
 wire \genblk2.pcpi_div.dividend[22] ;
 wire \genblk2.pcpi_div.dividend[23] ;
 wire \genblk2.pcpi_div.dividend[24] ;
 wire \genblk2.pcpi_div.dividend[25] ;
 wire \genblk2.pcpi_div.dividend[26] ;
 wire \genblk2.pcpi_div.dividend[27] ;
 wire \genblk2.pcpi_div.dividend[28] ;
 wire \genblk2.pcpi_div.dividend[29] ;
 wire \genblk2.pcpi_div.dividend[2] ;
 wire \genblk2.pcpi_div.dividend[30] ;
 wire \genblk2.pcpi_div.dividend[31] ;
 wire \genblk2.pcpi_div.dividend[3] ;
 wire \genblk2.pcpi_div.dividend[4] ;
 wire \genblk2.pcpi_div.dividend[5] ;
 wire \genblk2.pcpi_div.dividend[6] ;
 wire \genblk2.pcpi_div.dividend[7] ;
 wire \genblk2.pcpi_div.dividend[8] ;
 wire \genblk2.pcpi_div.dividend[9] ;
 wire \genblk2.pcpi_div.divisor[0] ;
 wire \genblk2.pcpi_div.divisor[10] ;
 wire \genblk2.pcpi_div.divisor[11] ;
 wire \genblk2.pcpi_div.divisor[12] ;
 wire \genblk2.pcpi_div.divisor[13] ;
 wire \genblk2.pcpi_div.divisor[14] ;
 wire \genblk2.pcpi_div.divisor[15] ;
 wire \genblk2.pcpi_div.divisor[16] ;
 wire \genblk2.pcpi_div.divisor[17] ;
 wire \genblk2.pcpi_div.divisor[18] ;
 wire \genblk2.pcpi_div.divisor[19] ;
 wire \genblk2.pcpi_div.divisor[1] ;
 wire \genblk2.pcpi_div.divisor[20] ;
 wire \genblk2.pcpi_div.divisor[21] ;
 wire \genblk2.pcpi_div.divisor[22] ;
 wire \genblk2.pcpi_div.divisor[23] ;
 wire \genblk2.pcpi_div.divisor[24] ;
 wire \genblk2.pcpi_div.divisor[25] ;
 wire \genblk2.pcpi_div.divisor[26] ;
 wire \genblk2.pcpi_div.divisor[27] ;
 wire \genblk2.pcpi_div.divisor[28] ;
 wire \genblk2.pcpi_div.divisor[29] ;
 wire \genblk2.pcpi_div.divisor[2] ;
 wire \genblk2.pcpi_div.divisor[30] ;
 wire \genblk2.pcpi_div.divisor[31] ;
 wire \genblk2.pcpi_div.divisor[32] ;
 wire \genblk2.pcpi_div.divisor[33] ;
 wire \genblk2.pcpi_div.divisor[34] ;
 wire \genblk2.pcpi_div.divisor[35] ;
 wire \genblk2.pcpi_div.divisor[36] ;
 wire \genblk2.pcpi_div.divisor[37] ;
 wire \genblk2.pcpi_div.divisor[38] ;
 wire \genblk2.pcpi_div.divisor[39] ;
 wire \genblk2.pcpi_div.divisor[3] ;
 wire \genblk2.pcpi_div.divisor[40] ;
 wire \genblk2.pcpi_div.divisor[41] ;
 wire \genblk2.pcpi_div.divisor[42] ;
 wire \genblk2.pcpi_div.divisor[43] ;
 wire \genblk2.pcpi_div.divisor[44] ;
 wire \genblk2.pcpi_div.divisor[45] ;
 wire \genblk2.pcpi_div.divisor[46] ;
 wire \genblk2.pcpi_div.divisor[47] ;
 wire \genblk2.pcpi_div.divisor[48] ;
 wire \genblk2.pcpi_div.divisor[49] ;
 wire \genblk2.pcpi_div.divisor[4] ;
 wire \genblk2.pcpi_div.divisor[50] ;
 wire \genblk2.pcpi_div.divisor[51] ;
 wire \genblk2.pcpi_div.divisor[52] ;
 wire \genblk2.pcpi_div.divisor[53] ;
 wire \genblk2.pcpi_div.divisor[54] ;
 wire \genblk2.pcpi_div.divisor[55] ;
 wire \genblk2.pcpi_div.divisor[56] ;
 wire \genblk2.pcpi_div.divisor[57] ;
 wire \genblk2.pcpi_div.divisor[58] ;
 wire \genblk2.pcpi_div.divisor[59] ;
 wire \genblk2.pcpi_div.divisor[5] ;
 wire \genblk2.pcpi_div.divisor[60] ;
 wire \genblk2.pcpi_div.divisor[61] ;
 wire \genblk2.pcpi_div.divisor[62] ;
 wire \genblk2.pcpi_div.divisor[6] ;
 wire \genblk2.pcpi_div.divisor[7] ;
 wire \genblk2.pcpi_div.divisor[8] ;
 wire \genblk2.pcpi_div.divisor[9] ;
 wire \genblk2.pcpi_div.instr_div ;
 wire \genblk2.pcpi_div.instr_divu ;
 wire \genblk2.pcpi_div.instr_rem ;
 wire \genblk2.pcpi_div.instr_remu ;
 wire \genblk2.pcpi_div.outsign ;
 wire \genblk2.pcpi_div.pcpi_rd[0] ;
 wire \genblk2.pcpi_div.pcpi_rd[10] ;
 wire \genblk2.pcpi_div.pcpi_rd[11] ;
 wire \genblk2.pcpi_div.pcpi_rd[12] ;
 wire \genblk2.pcpi_div.pcpi_rd[13] ;
 wire \genblk2.pcpi_div.pcpi_rd[14] ;
 wire \genblk2.pcpi_div.pcpi_rd[15] ;
 wire \genblk2.pcpi_div.pcpi_rd[16] ;
 wire \genblk2.pcpi_div.pcpi_rd[17] ;
 wire \genblk2.pcpi_div.pcpi_rd[18] ;
 wire \genblk2.pcpi_div.pcpi_rd[19] ;
 wire \genblk2.pcpi_div.pcpi_rd[1] ;
 wire \genblk2.pcpi_div.pcpi_rd[20] ;
 wire \genblk2.pcpi_div.pcpi_rd[21] ;
 wire \genblk2.pcpi_div.pcpi_rd[22] ;
 wire \genblk2.pcpi_div.pcpi_rd[23] ;
 wire \genblk2.pcpi_div.pcpi_rd[24] ;
 wire \genblk2.pcpi_div.pcpi_rd[25] ;
 wire \genblk2.pcpi_div.pcpi_rd[26] ;
 wire \genblk2.pcpi_div.pcpi_rd[27] ;
 wire \genblk2.pcpi_div.pcpi_rd[28] ;
 wire \genblk2.pcpi_div.pcpi_rd[29] ;
 wire \genblk2.pcpi_div.pcpi_rd[2] ;
 wire \genblk2.pcpi_div.pcpi_rd[30] ;
 wire \genblk2.pcpi_div.pcpi_rd[31] ;
 wire \genblk2.pcpi_div.pcpi_rd[3] ;
 wire \genblk2.pcpi_div.pcpi_rd[4] ;
 wire \genblk2.pcpi_div.pcpi_rd[5] ;
 wire \genblk2.pcpi_div.pcpi_rd[6] ;
 wire \genblk2.pcpi_div.pcpi_rd[7] ;
 wire \genblk2.pcpi_div.pcpi_rd[8] ;
 wire \genblk2.pcpi_div.pcpi_rd[9] ;
 wire \genblk2.pcpi_div.pcpi_ready ;
 wire \genblk2.pcpi_div.pcpi_wait ;
 wire \genblk2.pcpi_div.pcpi_wait_q ;
 wire \genblk2.pcpi_div.quotient[0] ;
 wire \genblk2.pcpi_div.quotient[10] ;
 wire \genblk2.pcpi_div.quotient[11] ;
 wire \genblk2.pcpi_div.quotient[12] ;
 wire \genblk2.pcpi_div.quotient[13] ;
 wire \genblk2.pcpi_div.quotient[14] ;
 wire \genblk2.pcpi_div.quotient[15] ;
 wire \genblk2.pcpi_div.quotient[16] ;
 wire \genblk2.pcpi_div.quotient[17] ;
 wire \genblk2.pcpi_div.quotient[18] ;
 wire \genblk2.pcpi_div.quotient[19] ;
 wire \genblk2.pcpi_div.quotient[1] ;
 wire \genblk2.pcpi_div.quotient[20] ;
 wire \genblk2.pcpi_div.quotient[21] ;
 wire \genblk2.pcpi_div.quotient[22] ;
 wire \genblk2.pcpi_div.quotient[23] ;
 wire \genblk2.pcpi_div.quotient[24] ;
 wire \genblk2.pcpi_div.quotient[25] ;
 wire \genblk2.pcpi_div.quotient[26] ;
 wire \genblk2.pcpi_div.quotient[27] ;
 wire \genblk2.pcpi_div.quotient[28] ;
 wire \genblk2.pcpi_div.quotient[29] ;
 wire \genblk2.pcpi_div.quotient[2] ;
 wire \genblk2.pcpi_div.quotient[30] ;
 wire \genblk2.pcpi_div.quotient[31] ;
 wire \genblk2.pcpi_div.quotient[3] ;
 wire \genblk2.pcpi_div.quotient[4] ;
 wire \genblk2.pcpi_div.quotient[5] ;
 wire \genblk2.pcpi_div.quotient[6] ;
 wire \genblk2.pcpi_div.quotient[7] ;
 wire \genblk2.pcpi_div.quotient[8] ;
 wire \genblk2.pcpi_div.quotient[9] ;
 wire \genblk2.pcpi_div.quotient_msk[0] ;
 wire \genblk2.pcpi_div.quotient_msk[10] ;
 wire \genblk2.pcpi_div.quotient_msk[11] ;
 wire \genblk2.pcpi_div.quotient_msk[12] ;
 wire \genblk2.pcpi_div.quotient_msk[13] ;
 wire \genblk2.pcpi_div.quotient_msk[14] ;
 wire \genblk2.pcpi_div.quotient_msk[15] ;
 wire \genblk2.pcpi_div.quotient_msk[16] ;
 wire \genblk2.pcpi_div.quotient_msk[17] ;
 wire \genblk2.pcpi_div.quotient_msk[18] ;
 wire \genblk2.pcpi_div.quotient_msk[19] ;
 wire \genblk2.pcpi_div.quotient_msk[1] ;
 wire \genblk2.pcpi_div.quotient_msk[20] ;
 wire \genblk2.pcpi_div.quotient_msk[21] ;
 wire \genblk2.pcpi_div.quotient_msk[22] ;
 wire \genblk2.pcpi_div.quotient_msk[23] ;
 wire \genblk2.pcpi_div.quotient_msk[24] ;
 wire \genblk2.pcpi_div.quotient_msk[25] ;
 wire \genblk2.pcpi_div.quotient_msk[26] ;
 wire \genblk2.pcpi_div.quotient_msk[27] ;
 wire \genblk2.pcpi_div.quotient_msk[28] ;
 wire \genblk2.pcpi_div.quotient_msk[29] ;
 wire \genblk2.pcpi_div.quotient_msk[2] ;
 wire \genblk2.pcpi_div.quotient_msk[30] ;
 wire \genblk2.pcpi_div.quotient_msk[31] ;
 wire \genblk2.pcpi_div.quotient_msk[3] ;
 wire \genblk2.pcpi_div.quotient_msk[4] ;
 wire \genblk2.pcpi_div.quotient_msk[5] ;
 wire \genblk2.pcpi_div.quotient_msk[6] ;
 wire \genblk2.pcpi_div.quotient_msk[7] ;
 wire \genblk2.pcpi_div.quotient_msk[8] ;
 wire \genblk2.pcpi_div.quotient_msk[9] ;
 wire \genblk2.pcpi_div.running ;
 wire instr_add;
 wire instr_addi;
 wire instr_and;
 wire instr_andi;
 wire instr_auipc;
 wire instr_beq;
 wire instr_bge;
 wire instr_bgeu;
 wire instr_blt;
 wire instr_bltu;
 wire instr_bne;
 wire instr_ecall_ebreak;
 wire instr_fence;
 wire instr_jal;
 wire instr_jalr;
 wire instr_lb;
 wire instr_lbu;
 wire instr_lh;
 wire instr_lhu;
 wire instr_lui;
 wire instr_lw;
 wire instr_or;
 wire instr_ori;
 wire instr_rdcycle;
 wire instr_rdcycleh;
 wire instr_rdinstr;
 wire instr_rdinstrh;
 wire instr_sb;
 wire instr_sh;
 wire instr_sll;
 wire instr_slli;
 wire instr_slt;
 wire instr_slti;
 wire instr_sltiu;
 wire instr_sltu;
 wire instr_sra;
 wire instr_srai;
 wire instr_srl;
 wire instr_srli;
 wire instr_sub;
 wire instr_sw;
 wire instr_xor;
 wire instr_xori;
 wire is_alu_reg_imm;
 wire is_alu_reg_reg;
 wire is_beq_bne_blt_bge_bltu_bgeu;
 wire is_compare;
 wire is_jalr_addi_slti_sltiu_xori_ori_andi;
 wire is_lb_lh_lw_lbu_lhu;
 wire is_lui_auipc_jal;
 wire is_sb_sh_sw;
 wire is_sll_srl_sra;
 wire is_slli_srli_srai;
 wire is_slti_blt_slt;
 wire is_sltiu_bltu_sltu;
 wire latched_branch;
 wire latched_is_lb;
 wire latched_is_lh;
 wire \latched_rd[0] ;
 wire \latched_rd[1] ;
 wire \latched_rd[2] ;
 wire \latched_rd[3] ;
 wire \latched_rd[4] ;
 wire latched_stalu;
 wire latched_store;
 wire net1275;
 wire net1276;
 wire mem_do_prefetch;
 wire mem_do_rdata;
 wire mem_do_rinst;
 wire mem_do_wdata;
 wire net1277;
 wire net1278;
 wire \mem_rdata_q[0] ;
 wire \mem_rdata_q[10] ;
 wire \mem_rdata_q[11] ;
 wire \mem_rdata_q[12] ;
 wire \mem_rdata_q[13] ;
 wire \mem_rdata_q[14] ;
 wire \mem_rdata_q[15] ;
 wire \mem_rdata_q[16] ;
 wire \mem_rdata_q[17] ;
 wire \mem_rdata_q[18] ;
 wire \mem_rdata_q[19] ;
 wire \mem_rdata_q[1] ;
 wire \mem_rdata_q[20] ;
 wire \mem_rdata_q[21] ;
 wire \mem_rdata_q[22] ;
 wire \mem_rdata_q[23] ;
 wire \mem_rdata_q[24] ;
 wire \mem_rdata_q[25] ;
 wire \mem_rdata_q[26] ;
 wire \mem_rdata_q[27] ;
 wire \mem_rdata_q[28] ;
 wire \mem_rdata_q[29] ;
 wire \mem_rdata_q[2] ;
 wire \mem_rdata_q[30] ;
 wire \mem_rdata_q[31] ;
 wire \mem_rdata_q[3] ;
 wire \mem_rdata_q[4] ;
 wire \mem_rdata_q[5] ;
 wire \mem_rdata_q[6] ;
 wire \mem_rdata_q[7] ;
 wire \mem_rdata_q[8] ;
 wire \mem_rdata_q[9] ;
 wire \mem_state[0] ;
 wire \mem_state[1] ;
 wire \mem_wordsize[0] ;
 wire \mem_wordsize[1] ;
 wire \mem_wordsize[2] ;
 wire pcpi_timeout;
 wire \pcpi_timeout_counter[0] ;
 wire \pcpi_timeout_counter[1] ;
 wire \pcpi_timeout_counter[2] ;
 wire \pcpi_timeout_counter[3] ;
 wire \reg_next_pc[10] ;
 wire \reg_next_pc[11] ;
 wire \reg_next_pc[12] ;
 wire \reg_next_pc[13] ;
 wire \reg_next_pc[14] ;
 wire \reg_next_pc[15] ;
 wire \reg_next_pc[16] ;
 wire \reg_next_pc[17] ;
 wire \reg_next_pc[18] ;
 wire \reg_next_pc[19] ;
 wire \reg_next_pc[1] ;
 wire \reg_next_pc[20] ;
 wire \reg_next_pc[21] ;
 wire \reg_next_pc[22] ;
 wire \reg_next_pc[23] ;
 wire \reg_next_pc[24] ;
 wire \reg_next_pc[25] ;
 wire \reg_next_pc[26] ;
 wire \reg_next_pc[27] ;
 wire \reg_next_pc[28] ;
 wire \reg_next_pc[29] ;
 wire \reg_next_pc[2] ;
 wire \reg_next_pc[30] ;
 wire \reg_next_pc[31] ;
 wire \reg_next_pc[3] ;
 wire \reg_next_pc[4] ;
 wire \reg_next_pc[5] ;
 wire \reg_next_pc[6] ;
 wire \reg_next_pc[7] ;
 wire \reg_next_pc[8] ;
 wire \reg_next_pc[9] ;
 wire \reg_out[0] ;
 wire \reg_out[10] ;
 wire \reg_out[11] ;
 wire \reg_out[12] ;
 wire \reg_out[13] ;
 wire \reg_out[14] ;
 wire \reg_out[15] ;
 wire \reg_out[16] ;
 wire \reg_out[17] ;
 wire \reg_out[18] ;
 wire \reg_out[19] ;
 wire \reg_out[1] ;
 wire \reg_out[20] ;
 wire \reg_out[21] ;
 wire \reg_out[22] ;
 wire \reg_out[23] ;
 wire \reg_out[24] ;
 wire \reg_out[25] ;
 wire \reg_out[26] ;
 wire \reg_out[27] ;
 wire \reg_out[28] ;
 wire \reg_out[29] ;
 wire \reg_out[2] ;
 wire \reg_out[30] ;
 wire \reg_out[31] ;
 wire \reg_out[3] ;
 wire \reg_out[4] ;
 wire \reg_out[5] ;
 wire \reg_out[6] ;
 wire \reg_out[7] ;
 wire \reg_out[8] ;
 wire \reg_out[9] ;
 wire \reg_pc[10] ;
 wire \reg_pc[11] ;
 wire \reg_pc[12] ;
 wire \reg_pc[13] ;
 wire \reg_pc[14] ;
 wire \reg_pc[15] ;
 wire \reg_pc[16] ;
 wire \reg_pc[17] ;
 wire \reg_pc[18] ;
 wire \reg_pc[19] ;
 wire \reg_pc[1] ;
 wire \reg_pc[20] ;
 wire \reg_pc[21] ;
 wire \reg_pc[22] ;
 wire \reg_pc[23] ;
 wire \reg_pc[24] ;
 wire \reg_pc[25] ;
 wire \reg_pc[26] ;
 wire \reg_pc[27] ;
 wire \reg_pc[28] ;
 wire \reg_pc[29] ;
 wire \reg_pc[2] ;
 wire \reg_pc[30] ;
 wire \reg_pc[31] ;
 wire \reg_pc[3] ;
 wire \reg_pc[4] ;
 wire \reg_pc[5] ;
 wire \reg_pc[6] ;
 wire \reg_pc[7] ;
 wire \reg_pc[8] ;
 wire \reg_pc[9] ;
 wire \reg_sh[0] ;
 wire \reg_sh[1] ;
 wire \reg_sh[2] ;
 wire \reg_sh[3] ;
 wire \reg_sh[4] ;
 wire net1279;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1280;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1281;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire clknet_leaf_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;

 sky130_fd_sc_hd__inv_2 _06751_ (.A(\genblk2.pcpi_div.divisor[20] ),
    .Y(_02359_));
 sky130_fd_sc_hd__inv_2 _06752_ (.A(\genblk2.pcpi_div.divisor[16] ),
    .Y(_02360_));
 sky130_fd_sc_hd__inv_2 _06753_ (.A(\genblk2.pcpi_div.divisor[8] ),
    .Y(_02361_));
 sky130_fd_sc_hd__inv_2 _06754_ (.A(\genblk2.pcpi_div.running ),
    .Y(_02362_));
 sky130_fd_sc_hd__inv_2 _06755_ (.A(net1072),
    .Y(_02363_));
 sky130_fd_sc_hd__inv_2 _06756_ (.A(net1145),
    .Y(_02364_));
 sky130_fd_sc_hd__inv_2 _06757_ (.A(instr_bgeu),
    .Y(_02365_));
 sky130_fd_sc_hd__inv_2 _06758_ (.A(instr_bge),
    .Y(_02366_));
 sky130_fd_sc_hd__inv_2 _06759_ (.A(latched_is_lb),
    .Y(_02367_));
 sky130_fd_sc_hd__inv_2 _06760_ (.A(latched_store),
    .Y(_02368_));
 sky130_fd_sc_hd__inv_2 _06761_ (.A(mem_do_rinst),
    .Y(_02369_));
 sky130_fd_sc_hd__inv_2 _06762_ (.A(net1089),
    .Y(_02370_));
 sky130_fd_sc_hd__inv_2 _06763_ (.A(\reg_pc[2] ),
    .Y(_02371_));
 sky130_fd_sc_hd__inv_2 _06764_ (.A(net2590),
    .Y(_02372_));
 sky130_fd_sc_hd__inv_2 _06765_ (.A(net2584),
    .Y(_02373_));
 sky130_fd_sc_hd__inv_2 _06766_ (.A(net2582),
    .Y(_02374_));
 sky130_fd_sc_hd__inv_2 _06767_ (.A(net2615),
    .Y(_02375_));
 sky130_fd_sc_hd__inv_2 _06768_ (.A(net2561),
    .Y(_02376_));
 sky130_fd_sc_hd__inv_2 _06769_ (.A(net1181),
    .Y(_02377_));
 sky130_fd_sc_hd__inv_2 _06770_ (.A(net1227),
    .Y(_02378_));
 sky130_fd_sc_hd__inv_2 _06771_ (.A(net1087),
    .Y(_02379_));
 sky130_fd_sc_hd__clkinv_4 _06772_ (.A(net1185),
    .Y(_02380_));
 sky130_fd_sc_hd__inv_2 _06773_ (.A(net1150),
    .Y(_02381_));
 sky130_fd_sc_hd__inv_2 _06774_ (.A(net2852),
    .Y(_02382_));
 sky130_fd_sc_hd__inv_2 _06775_ (.A(net1047),
    .Y(_02383_));
 sky130_fd_sc_hd__inv_2 _06776_ (.A(net1053),
    .Y(_02384_));
 sky130_fd_sc_hd__inv_2 _06777_ (.A(\reg_sh[0] ),
    .Y(_02385_));
 sky130_fd_sc_hd__inv_2 _06778_ (.A(net2768),
    .Y(_02386_));
 sky130_fd_sc_hd__inv_2 _06779_ (.A(net1061),
    .Y(_02387_));
 sky130_fd_sc_hd__inv_2 _06780_ (.A(\mem_rdata_q[14] ),
    .Y(_02388_));
 sky130_fd_sc_hd__inv_2 _06781_ (.A(\genblk2.pcpi_div.dividend[30] ),
    .Y(_02389_));
 sky130_fd_sc_hd__inv_2 _06782_ (.A(\genblk2.pcpi_div.dividend[14] ),
    .Y(_02390_));
 sky130_fd_sc_hd__inv_2 _06783_ (.A(\genblk2.pcpi_div.dividend[6] ),
    .Y(_02391_));
 sky130_fd_sc_hd__inv_2 _06784_ (.A(net1176),
    .Y(_02392_));
 sky130_fd_sc_hd__inv_2 _06785_ (.A(net1174),
    .Y(_02393_));
 sky130_fd_sc_hd__inv_2 _06786_ (.A(net240),
    .Y(_02394_));
 sky130_fd_sc_hd__inv_2 _06787_ (.A(net1161),
    .Y(_02395_));
 sky130_fd_sc_hd__inv_2 _06788_ (.A(net251),
    .Y(_02396_));
 sky130_fd_sc_hd__inv_2 _06789_ (.A(net254),
    .Y(_02397_));
 sky130_fd_sc_hd__inv_2 _06790_ (.A(net256),
    .Y(_02398_));
 sky130_fd_sc_hd__inv_2 _06791_ (.A(net255),
    .Y(_02399_));
 sky130_fd_sc_hd__inv_2 _06792_ (.A(\mem_rdata_q[2] ),
    .Y(_02400_));
 sky130_fd_sc_hd__inv_2 _06793_ (.A(\mem_rdata_q[5] ),
    .Y(_02401_));
 sky130_fd_sc_hd__inv_2 _06794_ (.A(net1044),
    .Y(_02402_));
 sky130_fd_sc_hd__inv_2 _06795_ (.A(net1031),
    .Y(_02403_));
 sky130_fd_sc_hd__inv_2 _06796_ (.A(net1028),
    .Y(_02404_));
 sky130_fd_sc_hd__inv_2 _06797_ (.A(net1026),
    .Y(_02405_));
 sky130_fd_sc_hd__inv_2 _06798_ (.A(net1024),
    .Y(_02406_));
 sky130_fd_sc_hd__inv_2 _06799_ (.A(net1018),
    .Y(_02407_));
 sky130_fd_sc_hd__inv_2 _06800_ (.A(net1016),
    .Y(_02408_));
 sky130_fd_sc_hd__inv_2 _06801_ (.A(net1012),
    .Y(_02409_));
 sky130_fd_sc_hd__inv_2 _06802_ (.A(net1009),
    .Y(_02410_));
 sky130_fd_sc_hd__inv_2 _06803_ (.A(net1006),
    .Y(_02411_));
 sky130_fd_sc_hd__inv_2 _06804_ (.A(net996),
    .Y(_02412_));
 sky130_fd_sc_hd__inv_2 _06805_ (.A(is_sltiu_bltu_sltu),
    .Y(_02413_));
 sky130_fd_sc_hd__inv_2 _06806_ (.A(net2515),
    .Y(_02414_));
 sky130_fd_sc_hd__inv_2 _06807_ (.A(\genblk1.genblk1.pcpi_mul.mul_counter[5] ),
    .Y(_02415_));
 sky130_fd_sc_hd__or2_1 _06808_ (.A(mem_do_rinst),
    .B(mem_do_prefetch),
    .X(_02416_));
 sky130_fd_sc_hd__or2_1 _06809_ (.A(mem_do_rdata),
    .B(net983),
    .X(_02417_));
 sky130_fd_sc_hd__nor2_1 _06810_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .Y(_02418_));
 sky130_fd_sc_hd__or2_1 _06811_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .X(_02419_));
 sky130_fd_sc_hd__and3_1 _06812_ (.A(net1234),
    .B(_02417_),
    .C(_02418_),
    .X(net96));
 sky130_fd_sc_hd__and3_1 _06813_ (.A(mem_do_wdata),
    .B(net1234),
    .C(_02418_),
    .X(net129));
 sky130_fd_sc_hd__or3_1 _06814_ (.A(net2572),
    .B(net2550),
    .C(net1649),
    .X(_00003_));
 sky130_fd_sc_hd__nor3_1 _06815_ (.A(net1133),
    .B(net1141),
    .C(net1137),
    .Y(_02420_));
 sky130_fd_sc_hd__or3_1 _06816_ (.A(net1134),
    .B(instr_rdcycleh),
    .C(instr_rdinstr),
    .X(_02421_));
 sky130_fd_sc_hd__or4_1 _06817_ (.A(instr_slli),
    .B(instr_sb),
    .C(instr_lw),
    .D(instr_jalr),
    .X(_02422_));
 sky130_fd_sc_hd__or4_1 _06818_ (.A(instr_beq),
    .B(instr_jal),
    .C(instr_rdcycle),
    .D(instr_srai),
    .X(_02423_));
 sky130_fd_sc_hd__or4_1 _06819_ (.A(instr_xori),
    .B(instr_addi),
    .C(instr_blt),
    .D(instr_bne),
    .X(_02424_));
 sky130_fd_sc_hd__or4_1 _06820_ (.A(instr_sll),
    .B(net1145),
    .C(instr_add),
    .D(instr_andi),
    .X(_02425_));
 sky130_fd_sc_hd__or4_1 _06821_ (.A(instr_fence),
    .B(instr_and),
    .C(instr_sra),
    .D(instr_xor),
    .X(_02426_));
 sky130_fd_sc_hd__or4_1 _06822_ (.A(_02423_),
    .B(_02424_),
    .C(_02425_),
    .D(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__or2_1 _06823_ (.A(instr_auipc),
    .B(instr_lui),
    .X(_02428_));
 sky130_fd_sc_hd__or4_1 _06824_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_bgeu),
    .D(instr_bge),
    .X(_02429_));
 sky130_fd_sc_hd__or4_1 _06825_ (.A(instr_sw),
    .B(instr_sh),
    .C(net970),
    .D(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__or4_1 _06826_ (.A(instr_srl),
    .B(instr_srli),
    .C(instr_lbu),
    .D(instr_lb),
    .X(_02431_));
 sky130_fd_sc_hd__nor2_2 _06827_ (.A(instr_or),
    .B(instr_ori),
    .Y(_02432_));
 sky130_fd_sc_hd__or2_1 _06828_ (.A(instr_or),
    .B(instr_ori),
    .X(_02433_));
 sky130_fd_sc_hd__or4_1 _06829_ (.A(instr_lhu),
    .B(instr_lh),
    .C(_02431_),
    .D(net966),
    .X(_02434_));
 sky130_fd_sc_hd__or3_1 _06830_ (.A(_02427_),
    .B(_02430_),
    .C(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__or4_2 _06831_ (.A(_00003_),
    .B(net975),
    .C(_02422_),
    .D(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__or2_1 _06832_ (.A(_02379_),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__nor2_1 _06833_ (.A(\genblk1.genblk1.pcpi_mul.pcpi_ready ),
    .B(net1113),
    .Y(_02438_));
 sky130_fd_sc_hd__and2b_1 _06834_ (.A_N(_02437_),
    .B(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__nor2_1 _06835_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_02440_));
 sky130_fd_sc_hd__and3b_1 _06836_ (.A_N(_02440_),
    .B(_02439_),
    .C(net1232),
    .X(_02441_));
 sky130_fd_sc_hd__and2_1 _06837_ (.A(net1232),
    .B(net2673),
    .X(_00582_));
 sky130_fd_sc_hd__a21o_1 _06838_ (.A1(net203),
    .A2(net1054),
    .B1(\mem_wordsize[0] ),
    .X(_02442_));
 sky130_fd_sc_hd__or2_4 _06839_ (.A(net1048),
    .B(net1051),
    .X(_02443_));
 sky130_fd_sc_hd__o211a_1 _06840_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .B1(_02442_),
    .C1(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__a21oi_2 _06841_ (.A1(mem_do_rinst),
    .A2(\reg_pc[1] ),
    .B1(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__or2_1 _06842_ (.A(net1208),
    .B(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__or3b_1 _06843_ (.A(_02441_),
    .B(_00582_),
    .C_N(_02446_),
    .X(_00004_));
 sky130_fd_sc_hd__or3_1 _06844_ (.A(mem_do_wdata),
    .B(mem_do_rdata),
    .C(mem_do_rinst),
    .X(_02447_));
 sky130_fd_sc_hd__and2_1 _06845_ (.A(\mem_state[0] ),
    .B(\mem_state[1] ),
    .X(_02448_));
 sky130_fd_sc_hd__and2_1 _06846_ (.A(net33),
    .B(net134),
    .X(_02449_));
 sky130_fd_sc_hd__nand2_2 _06847_ (.A(net33),
    .B(net134),
    .Y(_02450_));
 sky130_fd_sc_hd__a32o_2 _06848_ (.A1(_02419_),
    .A2(_02447_),
    .A3(net965),
    .B1(_02448_),
    .B2(mem_do_rinst),
    .X(_02451_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(net1232),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__nand2_1 _06850_ (.A(mem_do_prefetch),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_1 _06851_ (.A(net1061),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__nor3_1 _06852_ (.A(mem_do_rdata),
    .B(net1208),
    .C(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__or3_1 _06853_ (.A(instr_lhu),
    .B(instr_lw),
    .C(instr_lh),
    .X(_02456_));
 sky130_fd_sc_hd__or4b_1 _06854_ (.A(instr_lbu),
    .B(_02456_),
    .C(instr_lb),
    .D_N(net410),
    .X(_02457_));
 sky130_fd_sc_hd__a22o_1 _06855_ (.A1(mem_do_rdata),
    .A2(net1061),
    .B1(\cpu_state[6] ),
    .B2(mem_do_wdata),
    .X(_02458_));
 sky130_fd_sc_hd__nand2_1 _06856_ (.A(_02453_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__and4b_1 _06857_ (.A_N(mem_do_wdata),
    .B(net1232),
    .C(\cpu_state[6] ),
    .D(_02453_),
    .X(_02460_));
 sky130_fd_sc_hd__or4b_1 _06858_ (.A(instr_sw),
    .B(instr_sh),
    .C(instr_sb),
    .D_N(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__nor2_2 _06859_ (.A(net1060),
    .B(\cpu_state[6] ),
    .Y(_02462_));
 sky130_fd_sc_hd__or2_1 _06860_ (.A(net1060),
    .B(\cpu_state[6] ),
    .X(_02463_));
 sky130_fd_sc_hd__and3b_1 _06861_ (.A_N(_02451_),
    .B(net958),
    .C(mem_do_prefetch),
    .X(_02464_));
 sky130_fd_sc_hd__o21ai_1 _06862_ (.A1(net1089),
    .A2(net958),
    .B1(_02459_),
    .Y(_02465_));
 sky130_fd_sc_hd__nand2_1 _06863_ (.A(_02457_),
    .B(_02461_),
    .Y(_02466_));
 sky130_fd_sc_hd__or4_1 _06864_ (.A(net1208),
    .B(_02464_),
    .C(_02465_),
    .D(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__nor2_1 _06865_ (.A(_02370_),
    .B(net1208),
    .Y(_02468_));
 sky130_fd_sc_hd__a221o_1 _06866_ (.A1(instr_lw),
    .A2(net410),
    .B1(_02460_),
    .B2(instr_sw),
    .C1(net850),
    .X(_02469_));
 sky130_fd_sc_hd__a21o_1 _06867_ (.A1(net2132),
    .A2(_02467_),
    .B1(_02469_),
    .X(_00012_));
 sky130_fd_sc_hd__o21a_1 _06868_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(net410),
    .X(_02470_));
 sky130_fd_sc_hd__a221o_1 _06869_ (.A1(net2912),
    .A2(_02460_),
    .B1(_02467_),
    .B2(net1057),
    .C1(_02470_),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _06870_ (.A(net1152),
    .B(net970),
    .X(_00001_));
 sky130_fd_sc_hd__or3_1 _06871_ (.A(net2654),
    .B(instr_slti),
    .C(net2609),
    .X(_00002_));
 sky130_fd_sc_hd__nor2_1 _06872_ (.A(instr_rdcycle),
    .B(net975),
    .Y(_02471_));
 sky130_fd_sc_hd__o21a_1 _06873_ (.A1(instr_rdcycle),
    .A2(net975),
    .B1(net1088),
    .X(_02472_));
 sky130_fd_sc_hd__or2_1 _06874_ (.A(\reg_sh[3] ),
    .B(\reg_sh[2] ),
    .X(_02473_));
 sky130_fd_sc_hd__nor2_2 _06875_ (.A(\reg_sh[4] ),
    .B(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__or2_2 _06876_ (.A(\reg_sh[4] ),
    .B(_02473_),
    .X(_02475_));
 sky130_fd_sc_hd__nor2_1 _06877_ (.A(\reg_sh[1] ),
    .B(\reg_sh[0] ),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_1 _06878_ (.A(_02474_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__and3_1 _06879_ (.A(net1066),
    .B(_02474_),
    .C(_02476_),
    .X(_02478_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(net1185),
    .B(net850),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_4 _06881_ (.A(_02380_),
    .B(net985),
    .Y(_02480_));
 sky130_fd_sc_hd__nand2_1 _06882_ (.A(net1182),
    .B(net1149),
    .Y(_02481_));
 sky130_fd_sc_hd__a211o_1 _06883_ (.A1(net850),
    .A2(_02480_),
    .B1(_02478_),
    .C1(_02472_),
    .X(_02482_));
 sky130_fd_sc_hd__or2_1 _06884_ (.A(mem_do_prefetch),
    .B(_02452_),
    .X(_02483_));
 sky130_fd_sc_hd__nor2_1 _06885_ (.A(net961),
    .B(_02483_),
    .Y(_00814_));
 sky130_fd_sc_hd__nor2_1 _06886_ (.A(_02437_),
    .B(_02438_),
    .Y(_02484_));
 sky130_fd_sc_hd__o31a_1 _06887_ (.A1(_02482_),
    .A2(_00814_),
    .A3(_02484_),
    .B1(_02445_),
    .X(_02485_));
 sky130_fd_sc_hd__nand2_1 _06888_ (.A(net1072),
    .B(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_02486_));
 sky130_fd_sc_hd__nor2_1 _06889_ (.A(net991),
    .B(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_02487_));
 sky130_fd_sc_hd__a32o_1 _06890_ (.A1(net1072),
    .A2(is_beq_bne_blt_bge_bltu_bgeu),
    .A3(_02451_),
    .B1(_02380_),
    .B2(net1089),
    .X(_02488_));
 sky130_fd_sc_hd__o41a_1 _06891_ (.A1(net1208),
    .A2(_02485_),
    .A3(_02487_),
    .A4(_02488_),
    .B1(_02446_),
    .X(_00005_));
 sky130_fd_sc_hd__nand2_8 _06892_ (.A(net1184),
    .B(net985),
    .Y(_02489_));
 sky130_fd_sc_hd__nor2_1 _06893_ (.A(instr_jal),
    .B(_02479_),
    .Y(_02490_));
 sky130_fd_sc_hd__and2_1 _06894_ (.A(_02445_),
    .B(_02490_),
    .X(_00006_));
 sky130_fd_sc_hd__or3b_1 _06895_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_lui_auipc_jal),
    .C_N(net1088),
    .X(_02491_));
 sky130_fd_sc_hd__and2_1 _06896_ (.A(is_lb_lh_lw_lbu_lhu),
    .B(_02436_),
    .X(_02492_));
 sky130_fd_sc_hd__nor2_1 _06897_ (.A(_02491_),
    .B(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__and2_1 _06898_ (.A(net1232),
    .B(_02445_),
    .X(_02494_));
 sky130_fd_sc_hd__and4b_1 _06899_ (.A_N(is_slli_srli_srai),
    .B(_02471_),
    .C(_02493_),
    .D(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__a41o_1 _06900_ (.A1(net1232),
    .A2(_02439_),
    .A3(_02440_),
    .A4(_02445_),
    .B1(_02495_),
    .X(_00007_));
 sky130_fd_sc_hd__and4bb_1 _06901_ (.A_N(is_sll_srl_sra),
    .B_N(is_sb_sh_sw),
    .C(_02436_),
    .D(net1087),
    .X(_02496_));
 sky130_fd_sc_hd__o21a_1 _06902_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(is_lui_auipc_jal),
    .B1(net1088),
    .X(_02497_));
 sky130_fd_sc_hd__nor2_1 _06903_ (.A(_02451_),
    .B(_02486_),
    .Y(_02498_));
 sky130_fd_sc_hd__o31a_1 _06904_ (.A1(_02496_),
    .A2(_02497_),
    .A3(_02498_),
    .B1(_02494_),
    .X(_00008_));
 sky130_fd_sc_hd__o21a_1 _06905_ (.A1(instr_lhu),
    .A2(instr_lh),
    .B1(net410),
    .X(_02499_));
 sky130_fd_sc_hd__a221o_1 _06906_ (.A1(net2932),
    .A2(_02460_),
    .B1(_02467_),
    .B2(net1054),
    .C1(_02499_),
    .X(_00014_));
 sky130_fd_sc_hd__or3_1 _06907_ (.A(\genblk1.genblk1.pcpi_mul.instr_mulhsu ),
    .B(\genblk1.genblk1.pcpi_mul.instr_mulh ),
    .C(\genblk1.genblk1.pcpi_mul.instr_mulhu ),
    .X(_02500_));
 sky130_fd_sc_hd__or2_1 _06908_ (.A(net1316),
    .B(net956),
    .X(\genblk1.genblk1.pcpi_mul.instr_any_mul ));
 sky130_fd_sc_hd__and2_2 _06909_ (.A(net1066),
    .B(_02475_),
    .X(_02501_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(net1066),
    .B(_02475_),
    .Y(_02502_));
 sky130_fd_sc_hd__a22oi_1 _06911_ (.A1(net1084),
    .A2(is_sll_srl_sra),
    .B1(_02477_),
    .B2(net1068),
    .Y(_02503_));
 sky130_fd_sc_hd__nand2_1 _06912_ (.A(net1088),
    .B(net2671),
    .Y(_02504_));
 sky130_fd_sc_hd__a21boi_1 _06913_ (.A1(_02503_),
    .A2(_02504_),
    .B1_N(_02494_),
    .Y(_00009_));
 sky130_fd_sc_hd__a22o_1 _06914_ (.A1(net1084),
    .A2(is_sb_sh_sw),
    .B1(_02483_),
    .B2(\cpu_state[6] ),
    .X(_02505_));
 sky130_fd_sc_hd__and2_1 _06915_ (.A(_02494_),
    .B(_02505_),
    .X(_00010_));
 sky130_fd_sc_hd__and3_1 _06916_ (.A(net1088),
    .B(_02492_),
    .C(_02494_),
    .X(_02506_));
 sky130_fd_sc_hd__a31o_1 _06917_ (.A1(net1061),
    .A2(_02483_),
    .A3(_02494_),
    .B1(_02506_),
    .X(_00011_));
 sky130_fd_sc_hd__and2_1 _06918_ (.A(net1237),
    .B(net3031),
    .X(_00049_));
 sky130_fd_sc_hd__or2_2 _06919_ (.A(\genblk2.pcpi_div.instr_div ),
    .B(\genblk2.pcpi_div.instr_rem ),
    .X(_02507_));
 sky130_fd_sc_hd__nor2_1 _06920_ (.A(\genblk2.pcpi_div.instr_div ),
    .B(\genblk2.pcpi_div.instr_divu ),
    .Y(_02508_));
 sky130_fd_sc_hd__or2_2 _06921_ (.A(\genblk2.pcpi_div.instr_div ),
    .B(\genblk2.pcpi_div.instr_divu ),
    .X(_02509_));
 sky130_fd_sc_hd__o31a_1 _06922_ (.A1(\genblk2.pcpi_div.instr_rem ),
    .A2(net1370),
    .A3(_02509_),
    .B1(net1237),
    .X(_00048_));
 sky130_fd_sc_hd__and2_2 _06923_ (.A(net1237),
    .B(\genblk1.genblk1.pcpi_mul.mul_finish ),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _06924_ (.A0(\genblk2.pcpi_div.dividend[0] ),
    .A1(\genblk2.pcpi_div.quotient[0] ),
    .S(_02509_),
    .X(_00016_));
 sky130_fd_sc_hd__and3_1 _06925_ (.A(\genblk2.pcpi_div.quotient[0] ),
    .B(net1126),
    .C(\genblk2.pcpi_div.quotient[1] ),
    .X(_02510_));
 sky130_fd_sc_hd__a21oi_1 _06926_ (.A1(\genblk2.pcpi_div.quotient[0] ),
    .A2(net1126),
    .B1(net2999),
    .Y(_02511_));
 sky130_fd_sc_hd__and3_1 _06927_ (.A(\genblk2.pcpi_div.dividend[1] ),
    .B(\genblk2.pcpi_div.dividend[0] ),
    .C(net1126),
    .X(_02512_));
 sky130_fd_sc_hd__a21oi_1 _06928_ (.A1(\genblk2.pcpi_div.dividend[0] ),
    .A2(net1126),
    .B1(\genblk2.pcpi_div.dividend[1] ),
    .Y(_02513_));
 sky130_fd_sc_hd__or3_1 _06929_ (.A(_02509_),
    .B(_02512_),
    .C(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__o31ai_1 _06930_ (.A1(net953),
    .A2(_02510_),
    .A3(_02511_),
    .B1(_02514_),
    .Y(_00027_));
 sky130_fd_sc_hd__or2_1 _06931_ (.A(\genblk2.pcpi_div.quotient[0] ),
    .B(\genblk2.pcpi_div.quotient[1] ),
    .X(_02515_));
 sky130_fd_sc_hd__a21oi_1 _06932_ (.A1(net1126),
    .A2(_02515_),
    .B1(\genblk2.pcpi_div.quotient[2] ),
    .Y(_02516_));
 sky130_fd_sc_hd__a31o_1 _06933_ (.A1(net1126),
    .A2(\genblk2.pcpi_div.quotient[2] ),
    .A3(_02515_),
    .B1(net953),
    .X(_02517_));
 sky130_fd_sc_hd__o21ai_1 _06934_ (.A1(\genblk2.pcpi_div.dividend[1] ),
    .A2(\genblk2.pcpi_div.dividend[0] ),
    .B1(net1126),
    .Y(_02518_));
 sky130_fd_sc_hd__xnor2_1 _06935_ (.A(\genblk2.pcpi_div.dividend[2] ),
    .B(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__a2bb2o_1 _06936_ (.A1_N(_02516_),
    .A2_N(_02517_),
    .B1(_02519_),
    .B2(net953),
    .X(_00038_));
 sky130_fd_sc_hd__or3_1 _06937_ (.A(\genblk2.pcpi_div.dividend[2] ),
    .B(\genblk2.pcpi_div.dividend[1] ),
    .C(\genblk2.pcpi_div.dividend[0] ),
    .X(_02520_));
 sky130_fd_sc_hd__a21oi_1 _06938_ (.A1(\genblk2.pcpi_div.outsign ),
    .A2(_02520_),
    .B1(\genblk2.pcpi_div.dividend[3] ),
    .Y(_02521_));
 sky130_fd_sc_hd__a31o_1 _06939_ (.A1(\genblk2.pcpi_div.dividend[3] ),
    .A2(net1126),
    .A3(_02520_),
    .B1(net949),
    .X(_02522_));
 sky130_fd_sc_hd__o31a_1 _06940_ (.A1(\genblk2.pcpi_div.quotient[0] ),
    .A2(\genblk2.pcpi_div.quotient[1] ),
    .A3(\genblk2.pcpi_div.quotient[2] ),
    .B1(net1125),
    .X(_02523_));
 sky130_fd_sc_hd__xor2_1 _06941_ (.A(\genblk2.pcpi_div.quotient[3] ),
    .B(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__a2bb2o_1 _06942_ (.A1_N(_02521_),
    .A2_N(_02522_),
    .B1(_02524_),
    .B2(net949),
    .X(_00041_));
 sky130_fd_sc_hd__or4_2 _06943_ (.A(\genblk2.pcpi_div.quotient[0] ),
    .B(\genblk2.pcpi_div.quotient[1] ),
    .C(\genblk2.pcpi_div.quotient[2] ),
    .D(\genblk2.pcpi_div.quotient[3] ),
    .X(_02525_));
 sky130_fd_sc_hd__a21oi_1 _06944_ (.A1(net1125),
    .A2(_02525_),
    .B1(\genblk2.pcpi_div.quotient[4] ),
    .Y(_02526_));
 sky130_fd_sc_hd__a31o_1 _06945_ (.A1(net1125),
    .A2(\genblk2.pcpi_div.quotient[4] ),
    .A3(_02525_),
    .B1(net953),
    .X(_02527_));
 sky130_fd_sc_hd__or4_2 _06946_ (.A(\genblk2.pcpi_div.dividend[3] ),
    .B(\genblk2.pcpi_div.dividend[2] ),
    .C(\genblk2.pcpi_div.dividend[1] ),
    .D(\genblk2.pcpi_div.dividend[0] ),
    .X(_02528_));
 sky130_fd_sc_hd__a21oi_1 _06947_ (.A1(net1125),
    .A2(_02528_),
    .B1(net3058),
    .Y(_02529_));
 sky130_fd_sc_hd__a31o_1 _06948_ (.A1(\genblk2.pcpi_div.dividend[4] ),
    .A2(net1125),
    .A3(_02528_),
    .B1(net949),
    .X(_02530_));
 sky130_fd_sc_hd__o22ai_1 _06949_ (.A1(_02526_),
    .A2(_02527_),
    .B1(_02529_),
    .B2(_02530_),
    .Y(_00042_));
 sky130_fd_sc_hd__o21ai_1 _06950_ (.A1(\genblk2.pcpi_div.dividend[4] ),
    .A2(_02528_),
    .B1(net1125),
    .Y(_02531_));
 sky130_fd_sc_hd__xnor2_1 _06951_ (.A(\genblk2.pcpi_div.dividend[5] ),
    .B(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__o21ai_1 _06952_ (.A1(\genblk2.pcpi_div.quotient[4] ),
    .A2(_02525_),
    .B1(net1125),
    .Y(_02533_));
 sky130_fd_sc_hd__xnor2_1 _06953_ (.A(\genblk2.pcpi_div.quotient[5] ),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__mux2_1 _06954_ (.A0(_02532_),
    .A1(_02534_),
    .S(net949),
    .X(_00043_));
 sky130_fd_sc_hd__o31a_1 _06955_ (.A1(\genblk2.pcpi_div.quotient[4] ),
    .A2(\genblk2.pcpi_div.quotient[5] ),
    .A3(_02525_),
    .B1(net1125),
    .X(_02535_));
 sky130_fd_sc_hd__or2_1 _06956_ (.A(\genblk2.pcpi_div.quotient[6] ),
    .B(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__a21oi_1 _06957_ (.A1(\genblk2.pcpi_div.quotient[6] ),
    .A2(_02535_),
    .B1(net953),
    .Y(_02537_));
 sky130_fd_sc_hd__or3_1 _06958_ (.A(\genblk2.pcpi_div.dividend[5] ),
    .B(\genblk2.pcpi_div.dividend[4] ),
    .C(_02528_),
    .X(_02538_));
 sky130_fd_sc_hd__a21oi_1 _06959_ (.A1(net1126),
    .A2(_02538_),
    .B1(\genblk2.pcpi_div.dividend[6] ),
    .Y(_02539_));
 sky130_fd_sc_hd__a31o_1 _06960_ (.A1(\genblk2.pcpi_div.dividend[6] ),
    .A2(net1125),
    .A3(_02538_),
    .B1(net949),
    .X(_02540_));
 sky130_fd_sc_hd__a2bb2o_1 _06961_ (.A1_N(_02540_),
    .A2_N(_02539_),
    .B1(_02537_),
    .B2(_02536_),
    .X(_00044_));
 sky130_fd_sc_hd__or2_1 _06962_ (.A(\genblk2.pcpi_div.dividend[6] ),
    .B(_02538_),
    .X(_02541_));
 sky130_fd_sc_hd__a21oi_1 _06963_ (.A1(net1119),
    .A2(_02541_),
    .B1(\genblk2.pcpi_div.dividend[7] ),
    .Y(_02542_));
 sky130_fd_sc_hd__a31o_1 _06964_ (.A1(\genblk2.pcpi_div.dividend[7] ),
    .A2(net1119),
    .A3(_02541_),
    .B1(net948),
    .X(_02543_));
 sky130_fd_sc_hd__or4_1 _06965_ (.A(\genblk2.pcpi_div.quotient[4] ),
    .B(\genblk2.pcpi_div.quotient[5] ),
    .C(\genblk2.pcpi_div.quotient[6] ),
    .D(_02525_),
    .X(_02544_));
 sky130_fd_sc_hd__and3_1 _06966_ (.A(net1120),
    .B(\genblk2.pcpi_div.quotient[7] ),
    .C(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__a21oi_1 _06967_ (.A1(net1120),
    .A2(_02544_),
    .B1(\genblk2.pcpi_div.quotient[7] ),
    .Y(_02546_));
 sky130_fd_sc_hd__or3_1 _06968_ (.A(net951),
    .B(_02545_),
    .C(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__o21ai_1 _06969_ (.A1(_02542_),
    .A2(_02543_),
    .B1(_02547_),
    .Y(_00045_));
 sky130_fd_sc_hd__o21ai_1 _06970_ (.A1(\genblk2.pcpi_div.dividend[7] ),
    .A2(_02541_),
    .B1(net1118),
    .Y(_02548_));
 sky130_fd_sc_hd__xnor2_1 _06971_ (.A(\genblk2.pcpi_div.dividend[8] ),
    .B(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__or2_1 _06972_ (.A(\genblk2.pcpi_div.quotient[7] ),
    .B(_02544_),
    .X(_02550_));
 sky130_fd_sc_hd__a21oi_1 _06973_ (.A1(net1120),
    .A2(_02550_),
    .B1(\genblk2.pcpi_div.quotient[8] ),
    .Y(_02551_));
 sky130_fd_sc_hd__a31o_1 _06974_ (.A1(net1120),
    .A2(\genblk2.pcpi_div.quotient[8] ),
    .A3(_02550_),
    .B1(net951),
    .X(_02552_));
 sky130_fd_sc_hd__a2bb2o_1 _06975_ (.A1_N(_02551_),
    .A2_N(_02552_),
    .B1(net951),
    .B2(_02549_),
    .X(_00046_));
 sky130_fd_sc_hd__or3_1 _06976_ (.A(\genblk2.pcpi_div.dividend[8] ),
    .B(\genblk2.pcpi_div.dividend[7] ),
    .C(_02541_),
    .X(_02553_));
 sky130_fd_sc_hd__and3_1 _06977_ (.A(\genblk2.pcpi_div.dividend[9] ),
    .B(net1119),
    .C(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__a21oi_1 _06978_ (.A1(net1119),
    .A2(_02553_),
    .B1(\genblk2.pcpi_div.dividend[9] ),
    .Y(_02555_));
 sky130_fd_sc_hd__or3_1 _06979_ (.A(\genblk2.pcpi_div.quotient[7] ),
    .B(\genblk2.pcpi_div.quotient[8] ),
    .C(_02544_),
    .X(_02556_));
 sky130_fd_sc_hd__and3_1 _06980_ (.A(net1119),
    .B(\genblk2.pcpi_div.quotient[9] ),
    .C(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__a21oi_1 _06981_ (.A1(net1119),
    .A2(_02556_),
    .B1(\genblk2.pcpi_div.quotient[9] ),
    .Y(_02558_));
 sky130_fd_sc_hd__or3_1 _06982_ (.A(net951),
    .B(_02557_),
    .C(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__o31ai_1 _06983_ (.A1(net948),
    .A2(_02554_),
    .A3(_02555_),
    .B1(_02559_),
    .Y(_00047_));
 sky130_fd_sc_hd__o21ai_1 _06984_ (.A1(\genblk2.pcpi_div.dividend[9] ),
    .A2(_02553_),
    .B1(net1119),
    .Y(_02560_));
 sky130_fd_sc_hd__xnor2_1 _06985_ (.A(\genblk2.pcpi_div.dividend[10] ),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__or2_1 _06986_ (.A(\genblk2.pcpi_div.quotient[9] ),
    .B(_02556_),
    .X(_02562_));
 sky130_fd_sc_hd__a21oi_1 _06987_ (.A1(net1119),
    .A2(_02562_),
    .B1(\genblk2.pcpi_div.quotient[10] ),
    .Y(_02563_));
 sky130_fd_sc_hd__a31o_1 _06988_ (.A1(net1120),
    .A2(\genblk2.pcpi_div.quotient[10] ),
    .A3(_02562_),
    .B1(net951),
    .X(_02564_));
 sky130_fd_sc_hd__a2bb2o_1 _06989_ (.A1_N(_02563_),
    .A2_N(_02564_),
    .B1(net951),
    .B2(_02561_),
    .X(_00017_));
 sky130_fd_sc_hd__or3_1 _06990_ (.A(\genblk2.pcpi_div.quotient[9] ),
    .B(\genblk2.pcpi_div.quotient[10] ),
    .C(_02556_),
    .X(_02565_));
 sky130_fd_sc_hd__and3_1 _06991_ (.A(net1118),
    .B(\genblk2.pcpi_div.quotient[11] ),
    .C(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__a21oi_1 _06992_ (.A1(net1118),
    .A2(_02565_),
    .B1(\genblk2.pcpi_div.quotient[11] ),
    .Y(_02567_));
 sky130_fd_sc_hd__or3_1 _06993_ (.A(net951),
    .B(_02566_),
    .C(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__or3_1 _06994_ (.A(\genblk2.pcpi_div.dividend[10] ),
    .B(\genblk2.pcpi_div.dividend[9] ),
    .C(_02553_),
    .X(_02569_));
 sky130_fd_sc_hd__and3_1 _06995_ (.A(\genblk2.pcpi_div.dividend[11] ),
    .B(net1118),
    .C(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__a21oi_1 _06996_ (.A1(net1118),
    .A2(_02569_),
    .B1(\genblk2.pcpi_div.dividend[11] ),
    .Y(_02571_));
 sky130_fd_sc_hd__o31ai_1 _06997_ (.A1(net948),
    .A2(_02570_),
    .A3(_02571_),
    .B1(_02568_),
    .Y(_00018_));
 sky130_fd_sc_hd__or2_1 _06998_ (.A(\genblk2.pcpi_div.dividend[11] ),
    .B(_02569_),
    .X(_02572_));
 sky130_fd_sc_hd__a21oi_1 _06999_ (.A1(net1118),
    .A2(_02572_),
    .B1(net3025),
    .Y(_02573_));
 sky130_fd_sc_hd__a31o_1 _07000_ (.A1(\genblk2.pcpi_div.dividend[12] ),
    .A2(net1118),
    .A3(_02572_),
    .B1(net947),
    .X(_02574_));
 sky130_fd_sc_hd__or2_1 _07001_ (.A(\genblk2.pcpi_div.quotient[11] ),
    .B(_02565_),
    .X(_02575_));
 sky130_fd_sc_hd__a21oi_1 _07002_ (.A1(net1118),
    .A2(_02575_),
    .B1(net2961),
    .Y(_02576_));
 sky130_fd_sc_hd__a31o_1 _07003_ (.A1(net1118),
    .A2(\genblk2.pcpi_div.quotient[12] ),
    .A3(_02575_),
    .B1(net950),
    .X(_02577_));
 sky130_fd_sc_hd__o22ai_1 _07004_ (.A1(_02573_),
    .A2(_02574_),
    .B1(_02576_),
    .B2(_02577_),
    .Y(_00019_));
 sky130_fd_sc_hd__or2_1 _07005_ (.A(\genblk2.pcpi_div.dividend[12] ),
    .B(_02572_),
    .X(_02578_));
 sky130_fd_sc_hd__and3_1 _07006_ (.A(\genblk2.pcpi_div.dividend[13] ),
    .B(net1115),
    .C(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__a21oi_1 _07007_ (.A1(net1115),
    .A2(_02578_),
    .B1(\genblk2.pcpi_div.dividend[13] ),
    .Y(_02580_));
 sky130_fd_sc_hd__or3_1 _07008_ (.A(net947),
    .B(_02579_),
    .C(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__o21a_1 _07009_ (.A1(\genblk2.pcpi_div.quotient[12] ),
    .A2(_02575_),
    .B1(net1118),
    .X(_02582_));
 sky130_fd_sc_hd__xnor2_1 _07010_ (.A(\genblk2.pcpi_div.quotient[13] ),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__o21ai_1 _07011_ (.A1(net950),
    .A2(_02583_),
    .B1(_02581_),
    .Y(_00020_));
 sky130_fd_sc_hd__or2_1 _07012_ (.A(\genblk2.pcpi_div.dividend[13] ),
    .B(_02578_),
    .X(_02584_));
 sky130_fd_sc_hd__a21oi_1 _07013_ (.A1(net1115),
    .A2(_02584_),
    .B1(net3043),
    .Y(_02585_));
 sky130_fd_sc_hd__a31o_1 _07014_ (.A1(\genblk2.pcpi_div.dividend[14] ),
    .A2(net1115),
    .A3(_02584_),
    .B1(net947),
    .X(_02586_));
 sky130_fd_sc_hd__or3_1 _07015_ (.A(\genblk2.pcpi_div.quotient[12] ),
    .B(\genblk2.pcpi_div.quotient[13] ),
    .C(_02575_),
    .X(_02587_));
 sky130_fd_sc_hd__a21oi_1 _07016_ (.A1(net1115),
    .A2(_02587_),
    .B1(\genblk2.pcpi_div.quotient[14] ),
    .Y(_02588_));
 sky130_fd_sc_hd__a31o_1 _07017_ (.A1(net1115),
    .A2(\genblk2.pcpi_div.quotient[14] ),
    .A3(_02587_),
    .B1(net950),
    .X(_02589_));
 sky130_fd_sc_hd__or2_1 _07018_ (.A(_02588_),
    .B(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__o21ai_1 _07019_ (.A1(_02585_),
    .A2(_02586_),
    .B1(_02590_),
    .Y(_00021_));
 sky130_fd_sc_hd__o21ai_1 _07020_ (.A1(\genblk2.pcpi_div.dividend[14] ),
    .A2(_02584_),
    .B1(net1115),
    .Y(_02591_));
 sky130_fd_sc_hd__xnor2_1 _07021_ (.A(\genblk2.pcpi_div.dividend[15] ),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__or2_1 _07022_ (.A(\genblk2.pcpi_div.quotient[14] ),
    .B(_02587_),
    .X(_02593_));
 sky130_fd_sc_hd__a21oi_1 _07023_ (.A1(net1115),
    .A2(_02593_),
    .B1(\genblk2.pcpi_div.quotient[15] ),
    .Y(_02594_));
 sky130_fd_sc_hd__a31o_1 _07024_ (.A1(net1116),
    .A2(\genblk2.pcpi_div.quotient[15] ),
    .A3(_02593_),
    .B1(net950),
    .X(_02595_));
 sky130_fd_sc_hd__a2bb2o_1 _07025_ (.A1_N(_02594_),
    .A2_N(_02595_),
    .B1(net950),
    .B2(_02592_),
    .X(_00022_));
 sky130_fd_sc_hd__or3_1 _07026_ (.A(\genblk2.pcpi_div.dividend[15] ),
    .B(\genblk2.pcpi_div.dividend[14] ),
    .C(_02584_),
    .X(_02596_));
 sky130_fd_sc_hd__a21oi_1 _07027_ (.A1(net1114),
    .A2(_02596_),
    .B1(\genblk2.pcpi_div.dividend[16] ),
    .Y(_02597_));
 sky130_fd_sc_hd__a31o_1 _07028_ (.A1(\genblk2.pcpi_div.dividend[16] ),
    .A2(net1114),
    .A3(_02596_),
    .B1(net947),
    .X(_02598_));
 sky130_fd_sc_hd__or3_1 _07029_ (.A(\genblk2.pcpi_div.quotient[14] ),
    .B(\genblk2.pcpi_div.quotient[15] ),
    .C(_02587_),
    .X(_02599_));
 sky130_fd_sc_hd__a21oi_1 _07030_ (.A1(net1115),
    .A2(_02599_),
    .B1(\genblk2.pcpi_div.quotient[16] ),
    .Y(_02600_));
 sky130_fd_sc_hd__a31o_1 _07031_ (.A1(net1115),
    .A2(\genblk2.pcpi_div.quotient[16] ),
    .A3(_02599_),
    .B1(net950),
    .X(_02601_));
 sky130_fd_sc_hd__or2_1 _07032_ (.A(_02600_),
    .B(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__o21ai_1 _07033_ (.A1(_02597_),
    .A2(_02598_),
    .B1(_02602_),
    .Y(_00023_));
 sky130_fd_sc_hd__or2_1 _07034_ (.A(\genblk2.pcpi_div.dividend[16] ),
    .B(_02596_),
    .X(_02603_));
 sky130_fd_sc_hd__and3_1 _07035_ (.A(\genblk2.pcpi_div.dividend[17] ),
    .B(net1114),
    .C(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__a21oi_1 _07036_ (.A1(net1114),
    .A2(_02603_),
    .B1(\genblk2.pcpi_div.dividend[17] ),
    .Y(_02605_));
 sky130_fd_sc_hd__or3_1 _07037_ (.A(net947),
    .B(_02604_),
    .C(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__or2_1 _07038_ (.A(\genblk2.pcpi_div.quotient[16] ),
    .B(_02599_),
    .X(_02607_));
 sky130_fd_sc_hd__a21oi_1 _07039_ (.A1(net1114),
    .A2(_02607_),
    .B1(\genblk2.pcpi_div.quotient[17] ),
    .Y(_02608_));
 sky130_fd_sc_hd__a31o_1 _07040_ (.A1(net1114),
    .A2(\genblk2.pcpi_div.quotient[17] ),
    .A3(_02607_),
    .B1(net950),
    .X(_02609_));
 sky130_fd_sc_hd__o21ai_1 _07041_ (.A1(_02608_),
    .A2(_02609_),
    .B1(_02606_),
    .Y(_00024_));
 sky130_fd_sc_hd__or2_1 _07042_ (.A(\genblk2.pcpi_div.quotient[17] ),
    .B(_02607_),
    .X(_02610_));
 sky130_fd_sc_hd__and3_1 _07043_ (.A(net1116),
    .B(\genblk2.pcpi_div.quotient[18] ),
    .C(_02610_),
    .X(_02611_));
 sky130_fd_sc_hd__a21oi_1 _07044_ (.A1(net1116),
    .A2(_02610_),
    .B1(\genblk2.pcpi_div.quotient[18] ),
    .Y(_02612_));
 sky130_fd_sc_hd__or3_1 _07045_ (.A(net950),
    .B(_02611_),
    .C(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__or2_1 _07046_ (.A(\genblk2.pcpi_div.dividend[17] ),
    .B(_02603_),
    .X(_02614_));
 sky130_fd_sc_hd__a21oi_1 _07047_ (.A1(net1114),
    .A2(_02614_),
    .B1(net3021),
    .Y(_02615_));
 sky130_fd_sc_hd__a31o_1 _07048_ (.A1(\genblk2.pcpi_div.dividend[18] ),
    .A2(net1114),
    .A3(_02614_),
    .B1(net947),
    .X(_02616_));
 sky130_fd_sc_hd__o21ai_1 _07049_ (.A1(_02615_),
    .A2(_02616_),
    .B1(_02613_),
    .Y(_00025_));
 sky130_fd_sc_hd__o21ai_1 _07050_ (.A1(\genblk2.pcpi_div.quotient[18] ),
    .A2(_02610_),
    .B1(net1116),
    .Y(_02617_));
 sky130_fd_sc_hd__xnor2_1 _07051_ (.A(\genblk2.pcpi_div.quotient[19] ),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__or3_1 _07052_ (.A(\genblk2.pcpi_div.dividend[18] ),
    .B(\genblk2.pcpi_div.dividend[17] ),
    .C(_02603_),
    .X(_02619_));
 sky130_fd_sc_hd__a21oi_1 _07053_ (.A1(net1114),
    .A2(_02619_),
    .B1(\genblk2.pcpi_div.dividend[19] ),
    .Y(_02620_));
 sky130_fd_sc_hd__a31o_1 _07054_ (.A1(\genblk2.pcpi_div.dividend[19] ),
    .A2(net1114),
    .A3(_02619_),
    .B1(net947),
    .X(_02621_));
 sky130_fd_sc_hd__a2bb2o_1 _07055_ (.A1_N(_02621_),
    .A2_N(_02620_),
    .B1(_02618_),
    .B2(net947),
    .X(_00026_));
 sky130_fd_sc_hd__or2_1 _07056_ (.A(\genblk2.pcpi_div.dividend[19] ),
    .B(_02619_),
    .X(_02622_));
 sky130_fd_sc_hd__a21oi_1 _07057_ (.A1(net1117),
    .A2(_02622_),
    .B1(\genblk2.pcpi_div.dividend[20] ),
    .Y(_02623_));
 sky130_fd_sc_hd__a31o_1 _07058_ (.A1(\genblk2.pcpi_div.dividend[20] ),
    .A2(net1117),
    .A3(_02622_),
    .B1(net947),
    .X(_02624_));
 sky130_fd_sc_hd__or3_1 _07059_ (.A(\genblk2.pcpi_div.quotient[18] ),
    .B(\genblk2.pcpi_div.quotient[19] ),
    .C(_02610_),
    .X(_02625_));
 sky130_fd_sc_hd__a21oi_1 _07060_ (.A1(net1117),
    .A2(_02625_),
    .B1(net2761),
    .Y(_02626_));
 sky130_fd_sc_hd__a31o_1 _07061_ (.A1(net1117),
    .A2(\genblk2.pcpi_div.quotient[20] ),
    .A3(_02625_),
    .B1(net950),
    .X(_02627_));
 sky130_fd_sc_hd__o22ai_1 _07062_ (.A1(_02623_),
    .A2(_02624_),
    .B1(_02626_),
    .B2(_02627_),
    .Y(_00028_));
 sky130_fd_sc_hd__or2_1 _07063_ (.A(\genblk2.pcpi_div.quotient[20] ),
    .B(_02625_),
    .X(_02628_));
 sky130_fd_sc_hd__and3_1 _07064_ (.A(net1124),
    .B(\genblk2.pcpi_div.quotient[21] ),
    .C(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__a21oi_1 _07065_ (.A1(net1117),
    .A2(_02628_),
    .B1(\genblk2.pcpi_div.quotient[21] ),
    .Y(_02630_));
 sky130_fd_sc_hd__or2_1 _07066_ (.A(\genblk2.pcpi_div.dividend[20] ),
    .B(_02622_),
    .X(_02631_));
 sky130_fd_sc_hd__a21oi_1 _07067_ (.A1(net1117),
    .A2(_02631_),
    .B1(\genblk2.pcpi_div.dividend[21] ),
    .Y(_02632_));
 sky130_fd_sc_hd__a31o_1 _07068_ (.A1(\genblk2.pcpi_div.dividend[21] ),
    .A2(net1117),
    .A3(_02631_),
    .B1(net947),
    .X(_02633_));
 sky130_fd_sc_hd__o32a_1 _07069_ (.A1(net950),
    .A2(_02629_),
    .A3(_02630_),
    .B1(_02632_),
    .B2(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__inv_2 _07070_ (.A(_02634_),
    .Y(_00029_));
 sky130_fd_sc_hd__or2_1 _07071_ (.A(\genblk2.pcpi_div.dividend[21] ),
    .B(_02631_),
    .X(_02635_));
 sky130_fd_sc_hd__a21oi_1 _07072_ (.A1(net1117),
    .A2(_02635_),
    .B1(\genblk2.pcpi_div.dividend[22] ),
    .Y(_02636_));
 sky130_fd_sc_hd__a31o_1 _07073_ (.A1(\genblk2.pcpi_div.dividend[22] ),
    .A2(net1121),
    .A3(_02635_),
    .B1(net949),
    .X(_02637_));
 sky130_fd_sc_hd__o21ai_1 _07074_ (.A1(\genblk2.pcpi_div.quotient[21] ),
    .A2(_02628_),
    .B1(net1117),
    .Y(_02638_));
 sky130_fd_sc_hd__xnor2_1 _07075_ (.A(\genblk2.pcpi_div.quotient[22] ),
    .B(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hd__a2bb2o_1 _07076_ (.A1_N(_02636_),
    .A2_N(_02637_),
    .B1(_02639_),
    .B2(net949),
    .X(_00030_));
 sky130_fd_sc_hd__or3_1 _07077_ (.A(\genblk2.pcpi_div.dividend[22] ),
    .B(\genblk2.pcpi_div.dividend[21] ),
    .C(_02631_),
    .X(_02640_));
 sky130_fd_sc_hd__and3_1 _07078_ (.A(\genblk2.pcpi_div.dividend[23] ),
    .B(net1121),
    .C(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__a21oi_1 _07079_ (.A1(net1121),
    .A2(_02640_),
    .B1(\genblk2.pcpi_div.dividend[23] ),
    .Y(_02642_));
 sky130_fd_sc_hd__or3_1 _07080_ (.A(net948),
    .B(_02641_),
    .C(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__or3_1 _07081_ (.A(\genblk2.pcpi_div.quotient[21] ),
    .B(\genblk2.pcpi_div.quotient[22] ),
    .C(_02628_),
    .X(_02644_));
 sky130_fd_sc_hd__a21oi_1 _07082_ (.A1(net1121),
    .A2(_02644_),
    .B1(net2766),
    .Y(_02645_));
 sky130_fd_sc_hd__a31o_1 _07083_ (.A1(net1121),
    .A2(\genblk2.pcpi_div.quotient[23] ),
    .A3(_02644_),
    .B1(net953),
    .X(_02646_));
 sky130_fd_sc_hd__o21ai_1 _07084_ (.A1(_02645_),
    .A2(_02646_),
    .B1(_02643_),
    .Y(_00031_));
 sky130_fd_sc_hd__or2_1 _07085_ (.A(\genblk2.pcpi_div.dividend[23] ),
    .B(_02640_),
    .X(_02647_));
 sky130_fd_sc_hd__a21oi_1 _07086_ (.A1(net1121),
    .A2(_02647_),
    .B1(\genblk2.pcpi_div.dividend[24] ),
    .Y(_02648_));
 sky130_fd_sc_hd__a31o_1 _07087_ (.A1(\genblk2.pcpi_div.dividend[24] ),
    .A2(net1121),
    .A3(_02647_),
    .B1(net948),
    .X(_02649_));
 sky130_fd_sc_hd__or2_1 _07088_ (.A(\genblk2.pcpi_div.quotient[23] ),
    .B(_02644_),
    .X(_02650_));
 sky130_fd_sc_hd__a21o_1 _07089_ (.A1(net1121),
    .A2(_02650_),
    .B1(\genblk2.pcpi_div.quotient[24] ),
    .X(_02651_));
 sky130_fd_sc_hd__a31oi_1 _07090_ (.A1(net1121),
    .A2(\genblk2.pcpi_div.quotient[24] ),
    .A3(_02650_),
    .B1(net952),
    .Y(_02652_));
 sky130_fd_sc_hd__a2bb2o_1 _07091_ (.A1_N(_02648_),
    .A2_N(_02649_),
    .B1(_02651_),
    .B2(_02652_),
    .X(_00032_));
 sky130_fd_sc_hd__o21ai_1 _07092_ (.A1(\genblk2.pcpi_div.dividend[24] ),
    .A2(_02647_),
    .B1(net1121),
    .Y(_02653_));
 sky130_fd_sc_hd__xnor2_1 _07093_ (.A(\genblk2.pcpi_div.dividend[25] ),
    .B(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__a21oi_1 _07094_ (.A1(net1122),
    .A2(_02651_),
    .B1(\genblk2.pcpi_div.quotient[25] ),
    .Y(_02655_));
 sky130_fd_sc_hd__a31o_1 _07095_ (.A1(net1122),
    .A2(\genblk2.pcpi_div.quotient[25] ),
    .A3(_02651_),
    .B1(net952),
    .X(_02656_));
 sky130_fd_sc_hd__a2bb2o_1 _07096_ (.A1_N(_02655_),
    .A2_N(_02656_),
    .B1(net952),
    .B2(_02654_),
    .X(_00033_));
 sky130_fd_sc_hd__or3_1 _07097_ (.A(\genblk2.pcpi_div.dividend[25] ),
    .B(\genblk2.pcpi_div.dividend[24] ),
    .C(_02647_),
    .X(_02657_));
 sky130_fd_sc_hd__a21o_1 _07098_ (.A1(net1122),
    .A2(_02657_),
    .B1(\genblk2.pcpi_div.dividend[26] ),
    .X(_02658_));
 sky130_fd_sc_hd__a31oi_1 _07099_ (.A1(\genblk2.pcpi_div.dividend[26] ),
    .A2(net1122),
    .A3(_02657_),
    .B1(net948),
    .Y(_02659_));
 sky130_fd_sc_hd__o21a_1 _07100_ (.A1(\genblk2.pcpi_div.quotient[25] ),
    .A2(_02651_),
    .B1(net1122),
    .X(_02660_));
 sky130_fd_sc_hd__or2_1 _07101_ (.A(\genblk2.pcpi_div.quotient[26] ),
    .B(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__a21oi_1 _07102_ (.A1(\genblk2.pcpi_div.quotient[26] ),
    .A2(_02660_),
    .B1(net952),
    .Y(_02662_));
 sky130_fd_sc_hd__a22o_1 _07103_ (.A1(_02658_),
    .A2(_02659_),
    .B1(_02661_),
    .B2(_02662_),
    .X(_00034_));
 sky130_fd_sc_hd__a21oi_1 _07104_ (.A1(net1122),
    .A2(_02661_),
    .B1(net2854),
    .Y(_02663_));
 sky130_fd_sc_hd__a31o_1 _07105_ (.A1(net1123),
    .A2(\genblk2.pcpi_div.quotient[27] ),
    .A3(_02661_),
    .B1(net952),
    .X(_02664_));
 sky130_fd_sc_hd__a21oi_1 _07106_ (.A1(net1122),
    .A2(_02658_),
    .B1(\genblk2.pcpi_div.dividend[27] ),
    .Y(_02665_));
 sky130_fd_sc_hd__a31o_1 _07107_ (.A1(\genblk2.pcpi_div.dividend[27] ),
    .A2(net1122),
    .A3(_02658_),
    .B1(net949),
    .X(_02666_));
 sky130_fd_sc_hd__o22ai_1 _07108_ (.A1(_02663_),
    .A2(_02664_),
    .B1(_02665_),
    .B2(_02666_),
    .Y(_00035_));
 sky130_fd_sc_hd__o31a_1 _07109_ (.A1(\genblk2.pcpi_div.dividend[27] ),
    .A2(\genblk2.pcpi_div.dividend[26] ),
    .A3(_02657_),
    .B1(net1123),
    .X(_02667_));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(\genblk2.pcpi_div.dividend[28] ),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__or2_1 _07111_ (.A(\genblk2.pcpi_div.dividend[28] ),
    .B(_02667_),
    .X(_02669_));
 sky130_fd_sc_hd__o21a_1 _07112_ (.A1(\genblk2.pcpi_div.quotient[27] ),
    .A2(_02661_),
    .B1(net1123),
    .X(_02670_));
 sky130_fd_sc_hd__or2_1 _07113_ (.A(\genblk2.pcpi_div.quotient[28] ),
    .B(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__a21oi_1 _07114_ (.A1(\genblk2.pcpi_div.quotient[28] ),
    .A2(_02670_),
    .B1(net953),
    .Y(_02672_));
 sky130_fd_sc_hd__a32o_1 _07115_ (.A1(net952),
    .A2(_02668_),
    .A3(_02669_),
    .B1(_02671_),
    .B2(_02672_),
    .X(_00036_));
 sky130_fd_sc_hd__a211oi_1 _07116_ (.A1(net1122),
    .A2(\genblk2.pcpi_div.quotient[28] ),
    .B1(\genblk2.pcpi_div.quotient[29] ),
    .C1(_02670_),
    .Y(_02673_));
 sky130_fd_sc_hd__a311o_1 _07117_ (.A1(net1123),
    .A2(\genblk2.pcpi_div.quotient[29] ),
    .A3(_02671_),
    .B1(_02673_),
    .C1(net952),
    .X(_02674_));
 sky130_fd_sc_hd__a21oi_1 _07118_ (.A1(net1123),
    .A2(_02669_),
    .B1(\genblk2.pcpi_div.dividend[29] ),
    .Y(_02675_));
 sky130_fd_sc_hd__a31o_1 _07119_ (.A1(\genblk2.pcpi_div.dividend[29] ),
    .A2(net1123),
    .A3(_02669_),
    .B1(net948),
    .X(_02676_));
 sky130_fd_sc_hd__o21ai_1 _07120_ (.A1(_02675_),
    .A2(_02676_),
    .B1(_02674_),
    .Y(_00037_));
 sky130_fd_sc_hd__or2_1 _07121_ (.A(\genblk2.pcpi_div.dividend[29] ),
    .B(\genblk2.pcpi_div.dividend[28] ),
    .X(_02677_));
 sky130_fd_sc_hd__or4_1 _07122_ (.A(\genblk2.pcpi_div.dividend[27] ),
    .B(\genblk2.pcpi_div.dividend[26] ),
    .C(_02657_),
    .D(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__nand2_1 _07123_ (.A(net1124),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__o21ai_1 _07124_ (.A1(\genblk2.pcpi_div.quotient[29] ),
    .A2(_02671_),
    .B1(net1123),
    .Y(_02680_));
 sky130_fd_sc_hd__or2_1 _07125_ (.A(\genblk2.pcpi_div.quotient[30] ),
    .B(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__a21oi_1 _07126_ (.A1(\genblk2.pcpi_div.quotient[30] ),
    .A2(_02680_),
    .B1(net952),
    .Y(_02682_));
 sky130_fd_sc_hd__xnor2_1 _07127_ (.A(\genblk2.pcpi_div.dividend[30] ),
    .B(_02679_),
    .Y(_02683_));
 sky130_fd_sc_hd__o2bb2a_1 _07128_ (.A1_N(_02681_),
    .A2_N(_02682_),
    .B1(_02683_),
    .B2(net948),
    .X(_00039_));
 sky130_fd_sc_hd__o21ai_1 _07129_ (.A1(\genblk2.pcpi_div.dividend[30] ),
    .A2(_02678_),
    .B1(net1123),
    .Y(_02684_));
 sky130_fd_sc_hd__xnor2_1 _07130_ (.A(\genblk2.pcpi_div.dividend[31] ),
    .B(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__o31a_1 _07131_ (.A1(\genblk2.pcpi_div.quotient[29] ),
    .A2(\genblk2.pcpi_div.quotient[30] ),
    .A3(_02671_),
    .B1(net1123),
    .X(_02686_));
 sky130_fd_sc_hd__xor2_1 _07132_ (.A(\genblk2.pcpi_div.quotient[31] ),
    .B(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__mux2_1 _07133_ (.A0(_02685_),
    .A1(_02687_),
    .S(net948),
    .X(_00040_));
 sky130_fd_sc_hd__and2_1 _07134_ (.A(net1050),
    .B(net1054),
    .X(_02688_));
 sky130_fd_sc_hd__nand2_4 _07135_ (.A(net1048),
    .B(net1054),
    .Y(_02689_));
 sky130_fd_sc_hd__nand2b_2 _07136_ (.A_N(net1054),
    .B(net1057),
    .Y(_02690_));
 sky130_fd_sc_hd__a21bo_4 _07137_ (.A1(_02689_),
    .A2(net942),
    .B1_N(_02443_),
    .X(net130));
 sky130_fd_sc_hd__o211a_1 _07138_ (.A1(net1048),
    .A2(net31),
    .B1(net1057),
    .C1(net1052),
    .X(_02691_));
 sky130_fd_sc_hd__o21a_1 _07139_ (.A1(_02383_),
    .A2(net17),
    .B1(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__nor2_2 _07140_ (.A(net1054),
    .B(net1058),
    .Y(_02693_));
 sky130_fd_sc_hd__nor2_2 _07141_ (.A(_02383_),
    .B(net938),
    .Y(_02694_));
 sky130_fd_sc_hd__a31o_4 _07142_ (.A1(net1050),
    .A2(_02384_),
    .A3(net1056),
    .B1(_02688_),
    .X(_02695_));
 sky130_fd_sc_hd__a221o_1 _07143_ (.A1(net1),
    .A2(net130),
    .B1(_02695_),
    .B2(net8),
    .C1(_02692_),
    .X(_02696_));
 sky130_fd_sc_hd__mux2_1 _07144_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[0] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[0] ),
    .S(net1112),
    .X(_02697_));
 sky130_fd_sc_hd__a22o_1 _07145_ (.A1(net1051),
    .A2(net1066),
    .B1(_02697_),
    .B2(net1086),
    .X(_02698_));
 sky130_fd_sc_hd__a22o_1 _07146_ (.A1(\count_instr[32] ),
    .A2(net1130),
    .B1(net1140),
    .B2(\count_cycle[32] ),
    .X(_02699_));
 sky130_fd_sc_hd__a211o_1 _07147_ (.A1(\count_instr[0] ),
    .A2(net1135),
    .B1(net977),
    .C1(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__nor2_2 _07148_ (.A(net1080),
    .B(net1066),
    .Y(_02701_));
 sky130_fd_sc_hd__and3_2 _07149_ (.A(net991),
    .B(_02387_),
    .C(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__or4_1 _07150_ (.A(net1073),
    .B(net1084),
    .C(net1068),
    .D(net1061),
    .X(_02703_));
 sky130_fd_sc_hd__or2_1 _07151_ (.A(\count_cycle[0] ),
    .B(net975),
    .X(_02704_));
 sky130_fd_sc_hd__a32o_1 _07152_ (.A1(_02700_),
    .A2(net842),
    .A3(_02704_),
    .B1(_02696_),
    .B2(net1060),
    .X(_02705_));
 sky130_fd_sc_hd__a211o_1 _07153_ (.A1(net1073),
    .A2(\decoded_imm[0] ),
    .B1(_02698_),
    .C1(_02705_),
    .X(_06716_));
 sky130_fd_sc_hd__o211a_1 _07154_ (.A1(net1048),
    .A2(net32),
    .B1(net1057),
    .C1(net1052),
    .X(_02706_));
 sky130_fd_sc_hd__o21a_1 _07155_ (.A1(_02383_),
    .A2(net18),
    .B1(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__a221o_1 _07156_ (.A1(net12),
    .A2(net130),
    .B1(_02695_),
    .B2(net9),
    .C1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__or2_1 _07157_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .X(_02709_));
 sky130_fd_sc_hd__nand2_1 _07158_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_02710_));
 sky130_fd_sc_hd__mux2_1 _07159_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[1] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[1] ),
    .S(net1112),
    .X(_02711_));
 sky130_fd_sc_hd__a22o_1 _07160_ (.A1(\count_instr[1] ),
    .A2(net1136),
    .B1(\count_cycle[33] ),
    .B2(net1140),
    .X(_02712_));
 sky130_fd_sc_hd__a211o_1 _07161_ (.A1(\count_instr[33] ),
    .A2(net1130),
    .B1(net977),
    .C1(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__o211a_1 _07162_ (.A1(\count_cycle[1] ),
    .A2(net972),
    .B1(net842),
    .C1(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__a221o_1 _07163_ (.A1(net1049),
    .A2(net1067),
    .B1(_02711_),
    .B2(net1082),
    .C1(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__a21o_1 _07164_ (.A1(net1062),
    .A2(_02708_),
    .B1(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__a31o_1 _07165_ (.A1(net1071),
    .A2(_02709_),
    .A3(_02710_),
    .B1(_02716_),
    .X(_06727_));
 sky130_fd_sc_hd__o211a_1 _07166_ (.A1(net1048),
    .A2(net2),
    .B1(net1057),
    .C1(net1052),
    .X(_02717_));
 sky130_fd_sc_hd__o21a_1 _07167_ (.A1(_02383_),
    .A2(net19),
    .B1(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__a221o_1 _07168_ (.A1(net23),
    .A2(net130),
    .B1(_02695_),
    .B2(net10),
    .C1(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__a22o_1 _07169_ (.A1(\count_instr[34] ),
    .A2(net1130),
    .B1(net1135),
    .B2(\count_instr[2] ),
    .X(_02720_));
 sky130_fd_sc_hd__a211o_1 _07170_ (.A1(net1139),
    .A2(\count_cycle[34] ),
    .B1(net976),
    .C1(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__o211a_1 _07171_ (.A1(\count_cycle[2] ),
    .A2(net971),
    .B1(net842),
    .C1(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__nand2_1 _07172_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .Y(_02723_));
 sky130_fd_sc_hd__nor2_1 _07173_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .Y(_02724_));
 sky130_fd_sc_hd__or2_1 _07174_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .X(_02725_));
 sky130_fd_sc_hd__nand2_1 _07175_ (.A(_02723_),
    .B(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__a21oi_1 _07176_ (.A1(_02710_),
    .A2(_02726_),
    .B1(net991),
    .Y(_02727_));
 sky130_fd_sc_hd__o21a_1 _07177_ (.A1(_02710_),
    .A2(_02726_),
    .B1(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__mux2_1 _07178_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[2] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[2] ),
    .S(net1111),
    .X(_02729_));
 sky130_fd_sc_hd__a221o_1 _07179_ (.A1(net1062),
    .A2(_02719_),
    .B1(_02729_),
    .B2(net1082),
    .C1(_02722_),
    .X(_02730_));
 sky130_fd_sc_hd__a211o_1 _07180_ (.A1(net1065),
    .A2(net1045),
    .B1(_02728_),
    .C1(_02730_),
    .X(_06738_));
 sky130_fd_sc_hd__o21ai_1 _07181_ (.A1(_02710_),
    .A2(_02724_),
    .B1(_02723_),
    .Y(_02731_));
 sky130_fd_sc_hd__nand2_1 _07182_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_02732_));
 sky130_fd_sc_hd__or2_1 _07183_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .X(_02733_));
 sky130_fd_sc_hd__a21o_1 _07184_ (.A1(_02732_),
    .A2(_02733_),
    .B1(_02731_),
    .X(_02734_));
 sky130_fd_sc_hd__and3_1 _07185_ (.A(_02731_),
    .B(_02732_),
    .C(_02733_),
    .X(_02735_));
 sky130_fd_sc_hd__and3b_1 _07186_ (.A_N(_02735_),
    .B(net1074),
    .C(_02734_),
    .X(_02736_));
 sky130_fd_sc_hd__mux2_1 _07187_ (.A0(net3),
    .A1(net20),
    .S(net1048),
    .X(_02737_));
 sky130_fd_sc_hd__and3_1 _07188_ (.A(net1052),
    .B(net1057),
    .C(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__a221o_1 _07189_ (.A1(net26),
    .A2(net130),
    .B1(_02695_),
    .B2(net11),
    .C1(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__a22o_1 _07190_ (.A1(\count_instr[35] ),
    .A2(net1130),
    .B1(net1139),
    .B2(\count_cycle[35] ),
    .X(_02740_));
 sky130_fd_sc_hd__a211o_1 _07191_ (.A1(\count_instr[3] ),
    .A2(net1135),
    .B1(net976),
    .C1(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__o211a_1 _07192_ (.A1(\count_cycle[3] ),
    .A2(net971),
    .B1(net842),
    .C1(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__mux2_1 _07193_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[3] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[3] ),
    .S(net1111),
    .X(_02743_));
 sky130_fd_sc_hd__a221o_1 _07194_ (.A1(net1062),
    .A2(_02739_),
    .B1(_02743_),
    .B2(net1082),
    .C1(_02742_),
    .X(_02744_));
 sky130_fd_sc_hd__a211o_1 _07195_ (.A1(net1065),
    .A2(net1044),
    .B1(_02736_),
    .C1(_02744_),
    .X(_06741_));
 sky130_fd_sc_hd__nand2_1 _07196_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .Y(_02745_));
 sky130_fd_sc_hd__inv_2 _07197_ (.A(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__or2_1 _07198_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .X(_02747_));
 sky130_fd_sc_hd__a21bo_1 _07199_ (.A1(_02731_),
    .A2(_02733_),
    .B1_N(_02732_),
    .X(_02748_));
 sky130_fd_sc_hd__a21o_1 _07200_ (.A1(_02745_),
    .A2(_02747_),
    .B1(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__nand3_1 _07201_ (.A(_02745_),
    .B(_02747_),
    .C(_02748_),
    .Y(_02750_));
 sky130_fd_sc_hd__and3_1 _07202_ (.A(net1074),
    .B(_02749_),
    .C(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__mux2_1 _07203_ (.A0(net4),
    .A1(net21),
    .S(net1048),
    .X(_02752_));
 sky130_fd_sc_hd__and3_1 _07204_ (.A(net203),
    .B(net1057),
    .C(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__a221o_1 _07205_ (.A1(net27),
    .A2(net130),
    .B1(_02695_),
    .B2(net13),
    .C1(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _07206_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[4] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[4] ),
    .S(net1111),
    .X(_02755_));
 sky130_fd_sc_hd__a22o_1 _07207_ (.A1(net1065),
    .A2(net1042),
    .B1(_02755_),
    .B2(net1079),
    .X(_02756_));
 sky130_fd_sc_hd__a211o_1 _07208_ (.A1(net1062),
    .A2(_02754_),
    .B1(_02756_),
    .C1(net842),
    .X(_02757_));
 sky130_fd_sc_hd__a22o_1 _07209_ (.A1(\count_instr[36] ),
    .A2(net1130),
    .B1(net1135),
    .B2(\count_instr[4] ),
    .X(_02758_));
 sky130_fd_sc_hd__a221o_1 _07210_ (.A1(net1139),
    .A2(\count_cycle[36] ),
    .B1(\count_cycle[4] ),
    .B2(net976),
    .C1(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__o22a_1 _07211_ (.A1(_02751_),
    .A2(_02757_),
    .B1(_02759_),
    .B2(_02703_),
    .X(_06742_));
 sky130_fd_sc_hd__nand2_1 _07212_ (.A(_02745_),
    .B(_02750_),
    .Y(_02760_));
 sky130_fd_sc_hd__or2_1 _07213_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .X(_02761_));
 sky130_fd_sc_hd__nand2_1 _07214_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_02762_));
 sky130_fd_sc_hd__nand3_1 _07215_ (.A(_02760_),
    .B(_02761_),
    .C(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__a21o_1 _07216_ (.A1(_02761_),
    .A2(_02762_),
    .B1(_02760_),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _07217_ (.A0(net5),
    .A1(net22),
    .S(net1048),
    .X(_02765_));
 sky130_fd_sc_hd__and3_1 _07218_ (.A(net1052),
    .B(net1057),
    .C(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__a221o_1 _07219_ (.A1(net28),
    .A2(net130),
    .B1(_02695_),
    .B2(net14),
    .C1(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__a22o_1 _07220_ (.A1(\count_instr[37] ),
    .A2(net1130),
    .B1(net1135),
    .B2(\count_instr[5] ),
    .X(_02768_));
 sky130_fd_sc_hd__a211o_1 _07221_ (.A1(net1139),
    .A2(\count_cycle[37] ),
    .B1(net976),
    .C1(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__o211a_1 _07222_ (.A1(\count_cycle[5] ),
    .A2(net971),
    .B1(net841),
    .C1(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__mux2_1 _07223_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[5] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[5] ),
    .S(net1111),
    .X(_02771_));
 sky130_fd_sc_hd__a221o_1 _07224_ (.A1(net1065),
    .A2(net1040),
    .B1(_02771_),
    .B2(net1078),
    .C1(_02770_),
    .X(_02772_));
 sky130_fd_sc_hd__a21o_1 _07225_ (.A1(net1062),
    .A2(_02767_),
    .B1(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__a31o_1 _07226_ (.A1(net1071),
    .A2(_02763_),
    .A3(_02764_),
    .B1(_02773_),
    .X(_06743_));
 sky130_fd_sc_hd__nand2_1 _07227_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .Y(_02774_));
 sky130_fd_sc_hd__inv_2 _07228_ (.A(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__or2_1 _07229_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .X(_02776_));
 sky130_fd_sc_hd__a221o_1 _07230_ (.A1(\reg_pc[5] ),
    .A2(\decoded_imm[5] ),
    .B1(_02747_),
    .B2(_02748_),
    .C1(_02746_),
    .X(_02777_));
 sky130_fd_sc_hd__and2_1 _07231_ (.A(_02761_),
    .B(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__nand3_1 _07232_ (.A(_02774_),
    .B(_02776_),
    .C(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__a21o_1 _07233_ (.A1(_02774_),
    .A2(_02776_),
    .B1(_02778_),
    .X(_02780_));
 sky130_fd_sc_hd__o211a_1 _07234_ (.A1(net1048),
    .A2(net6),
    .B1(net1057),
    .C1(net1052),
    .X(_02781_));
 sky130_fd_sc_hd__o21a_1 _07235_ (.A1(_02383_),
    .A2(net24),
    .B1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__a221o_1 _07236_ (.A1(net29),
    .A2(net130),
    .B1(_02695_),
    .B2(net15),
    .C1(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__a22o_1 _07237_ (.A1(\count_instr[38] ),
    .A2(net1130),
    .B1(net1139),
    .B2(\count_cycle[38] ),
    .X(_02784_));
 sky130_fd_sc_hd__a211o_1 _07238_ (.A1(\count_instr[6] ),
    .A2(net1135),
    .B1(net976),
    .C1(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__o211a_1 _07239_ (.A1(\count_cycle[6] ),
    .A2(net972),
    .B1(net841),
    .C1(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _07240_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[6] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[6] ),
    .S(net1110),
    .X(_02787_));
 sky130_fd_sc_hd__a221o_1 _07241_ (.A1(net1064),
    .A2(net1038),
    .B1(_02787_),
    .B2(net1078),
    .C1(_02786_),
    .X(_02788_));
 sky130_fd_sc_hd__a21o_1 _07242_ (.A1(net1062),
    .A2(_02783_),
    .B1(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__a31o_1 _07243_ (.A1(net1071),
    .A2(_02779_),
    .A3(_02780_),
    .B1(_02789_),
    .X(_06744_));
 sky130_fd_sc_hd__a31oi_1 _07244_ (.A1(_02761_),
    .A2(_02776_),
    .A3(_02777_),
    .B1(_02775_),
    .Y(_02790_));
 sky130_fd_sc_hd__and2_1 _07245_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .X(_02791_));
 sky130_fd_sc_hd__inv_2 _07246_ (.A(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__nor2_1 _07247_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_02793_));
 sky130_fd_sc_hd__or2_1 _07248_ (.A(_02791_),
    .B(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__or2_1 _07249_ (.A(_02790_),
    .B(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__a21oi_1 _07250_ (.A1(_02790_),
    .A2(_02794_),
    .B1(net991),
    .Y(_02796_));
 sky130_fd_sc_hd__or2_1 _07251_ (.A(_02383_),
    .B(net25),
    .X(_02797_));
 sky130_fd_sc_hd__o2111a_1 _07252_ (.A1(net1048),
    .A2(net7),
    .B1(_02797_),
    .C1(net1052),
    .D1(net1057),
    .X(_02798_));
 sky130_fd_sc_hd__a221o_1 _07253_ (.A1(net30),
    .A2(net130),
    .B1(_02695_),
    .B2(net16),
    .C1(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__a22o_1 _07254_ (.A1(\count_instr[39] ),
    .A2(net1130),
    .B1(net1135),
    .B2(\count_instr[7] ),
    .X(_02800_));
 sky130_fd_sc_hd__a211o_1 _07255_ (.A1(net1139),
    .A2(\count_cycle[39] ),
    .B1(net976),
    .C1(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__o211a_1 _07256_ (.A1(\count_cycle[7] ),
    .A2(net971),
    .B1(net841),
    .C1(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _07257_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[7] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[7] ),
    .S(net1110),
    .X(_02803_));
 sky130_fd_sc_hd__a221o_1 _07258_ (.A1(net1064),
    .A2(net1037),
    .B1(_02803_),
    .B2(net1078),
    .C1(_02802_),
    .X(_02804_));
 sky130_fd_sc_hd__a21o_1 _07259_ (.A1(net1062),
    .A2(_02799_),
    .B1(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__a21o_1 _07260_ (.A1(_02795_),
    .A2(_02796_),
    .B1(_02805_),
    .X(_06745_));
 sky130_fd_sc_hd__or2_1 _07261_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .X(_02806_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _07263_ (.A(_02806_),
    .B(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__a21o_1 _07264_ (.A1(_02792_),
    .A2(_02795_),
    .B1(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__nand3_1 _07265_ (.A(_02792_),
    .B(_02795_),
    .C(_02808_),
    .Y(_02810_));
 sky130_fd_sc_hd__and2_2 _07266_ (.A(latched_is_lb),
    .B(_02799_),
    .X(_02811_));
 sky130_fd_sc_hd__o21a_1 _07267_ (.A1(_02367_),
    .A2(latched_is_lh),
    .B1(net942),
    .X(_02812_));
 sky130_fd_sc_hd__o221a_1 _07268_ (.A1(net17),
    .A2(_02689_),
    .B1(_02694_),
    .B2(net31),
    .C1(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__o21a_1 _07269_ (.A1(_02811_),
    .A2(_02813_),
    .B1(net1060),
    .X(_02814_));
 sky130_fd_sc_hd__a22o_1 _07270_ (.A1(\count_instr[40] ),
    .A2(net1131),
    .B1(net1136),
    .B2(\count_instr[8] ),
    .X(_02815_));
 sky130_fd_sc_hd__a211o_1 _07271_ (.A1(net1139),
    .A2(\count_cycle[40] ),
    .B1(net976),
    .C1(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__o211a_1 _07272_ (.A1(\count_cycle[8] ),
    .A2(net971),
    .B1(net841),
    .C1(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_1 _07273_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[8] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[8] ),
    .S(net1110),
    .X(_02818_));
 sky130_fd_sc_hd__a221o_1 _07274_ (.A1(net1064),
    .A2(net1034),
    .B1(_02818_),
    .B2(net1079),
    .C1(_02817_),
    .X(_02819_));
 sky130_fd_sc_hd__or2_1 _07275_ (.A(_02814_),
    .B(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__a31o_1 _07276_ (.A1(net1071),
    .A2(_02809_),
    .A3(_02810_),
    .B1(_02820_),
    .X(_06746_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_02821_));
 sky130_fd_sc_hd__nor2_1 _07278_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_02822_));
 sky130_fd_sc_hd__or2_1 _07279_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .X(_02823_));
 sky130_fd_sc_hd__nand2_1 _07280_ (.A(_02821_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__a21o_1 _07281_ (.A1(_02807_),
    .A2(_02809_),
    .B1(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(net1071),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__a31o_1 _07283_ (.A1(_02807_),
    .A2(_02809_),
    .A3(_02824_),
    .B1(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__o221a_1 _07284_ (.A1(net18),
    .A2(_02689_),
    .B1(_02694_),
    .B2(net32),
    .C1(_02812_),
    .X(_02828_));
 sky130_fd_sc_hd__o21a_1 _07285_ (.A1(_02811_),
    .A2(_02828_),
    .B1(net1060),
    .X(_02829_));
 sky130_fd_sc_hd__a22o_1 _07286_ (.A1(\count_instr[41] ),
    .A2(net1130),
    .B1(net1135),
    .B2(\count_instr[9] ),
    .X(_02830_));
 sky130_fd_sc_hd__a211o_1 _07287_ (.A1(net1139),
    .A2(\count_cycle[41] ),
    .B1(net976),
    .C1(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__o211a_1 _07288_ (.A1(\count_cycle[9] ),
    .A2(net971),
    .B1(net841),
    .C1(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _07289_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[9] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[9] ),
    .S(net1110),
    .X(_02833_));
 sky130_fd_sc_hd__a221o_1 _07290_ (.A1(net1063),
    .A2(net1031),
    .B1(_02833_),
    .B2(net1077),
    .C1(_02829_),
    .X(_02834_));
 sky130_fd_sc_hd__or3b_1 _07291_ (.A(_02834_),
    .B(_02832_),
    .C_N(_02827_),
    .X(_06747_));
 sky130_fd_sc_hd__xnor2_1 _07292_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .Y(_02835_));
 sky130_fd_sc_hd__and3_1 _07293_ (.A(_02821_),
    .B(_02825_),
    .C(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__a21oi_1 _07294_ (.A1(_02821_),
    .A2(_02825_),
    .B1(_02835_),
    .Y(_02837_));
 sky130_fd_sc_hd__or3_1 _07295_ (.A(net991),
    .B(_02836_),
    .C(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__o221a_1 _07296_ (.A1(net19),
    .A2(_02689_),
    .B1(_02694_),
    .B2(net2),
    .C1(_02812_),
    .X(_02839_));
 sky130_fd_sc_hd__o21a_1 _07297_ (.A1(_02811_),
    .A2(_02839_),
    .B1(net1060),
    .X(_02840_));
 sky130_fd_sc_hd__a22o_1 _07298_ (.A1(\count_instr[42] ),
    .A2(net1131),
    .B1(net1135),
    .B2(\count_instr[10] ),
    .X(_02841_));
 sky130_fd_sc_hd__a211o_1 _07299_ (.A1(net1139),
    .A2(\count_cycle[42] ),
    .B1(net976),
    .C1(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__o211a_1 _07300_ (.A1(\count_cycle[10] ),
    .A2(net972),
    .B1(net841),
    .C1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _07301_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[10] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[10] ),
    .S(net1110),
    .X(_02844_));
 sky130_fd_sc_hd__a221o_1 _07302_ (.A1(net1063),
    .A2(net1029),
    .B1(_02844_),
    .B2(net1077),
    .C1(_02840_),
    .X(_02845_));
 sky130_fd_sc_hd__or3b_1 _07303_ (.A(_02845_),
    .B(_02843_),
    .C_N(_02838_),
    .X(_06717_));
 sky130_fd_sc_hd__nand2_1 _07304_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .Y(_02846_));
 sky130_fd_sc_hd__or2_1 _07305_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .X(_02847_));
 sky130_fd_sc_hd__nand2_1 _07306_ (.A(_02846_),
    .B(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hd__a21o_1 _07307_ (.A1(\reg_pc[10] ),
    .A2(\decoded_imm[10] ),
    .B1(_02837_),
    .X(_02849_));
 sky130_fd_sc_hd__xor2_1 _07308_ (.A(_02848_),
    .B(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__nor2_1 _07309_ (.A(net991),
    .B(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__o221a_1 _07310_ (.A1(net20),
    .A2(_02689_),
    .B1(_02694_),
    .B2(net3),
    .C1(_02812_),
    .X(_02852_));
 sky130_fd_sc_hd__o21a_1 _07311_ (.A1(_02811_),
    .A2(_02852_),
    .B1(net1060),
    .X(_02853_));
 sky130_fd_sc_hd__a22o_1 _07312_ (.A1(\count_instr[43] ),
    .A2(net1131),
    .B1(net1135),
    .B2(\count_instr[11] ),
    .X(_02854_));
 sky130_fd_sc_hd__a211o_1 _07313_ (.A1(net1139),
    .A2(\count_cycle[43] ),
    .B1(net976),
    .C1(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__o211a_1 _07314_ (.A1(\count_cycle[11] ),
    .A2(net971),
    .B1(net841),
    .C1(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__mux2_1 _07315_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[11] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[11] ),
    .S(net1110),
    .X(_02857_));
 sky130_fd_sc_hd__a221o_1 _07316_ (.A1(net1063),
    .A2(net1028),
    .B1(_02857_),
    .B2(net1077),
    .C1(_02853_),
    .X(_02858_));
 sky130_fd_sc_hd__or3_1 _07317_ (.A(_02851_),
    .B(_02856_),
    .C(_02858_),
    .X(_06718_));
 sky130_fd_sc_hd__or3_1 _07318_ (.A(_02824_),
    .B(_02835_),
    .C(_02848_),
    .X(_02859_));
 sky130_fd_sc_hd__a211o_1 _07319_ (.A1(_02792_),
    .A2(_02795_),
    .B1(_02808_),
    .C1(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__o21a_1 _07320_ (.A1(_02807_),
    .A2(_02822_),
    .B1(_02821_),
    .X(_02861_));
 sky130_fd_sc_hd__o31ai_1 _07321_ (.A1(_02835_),
    .A2(_02848_),
    .A3(_02861_),
    .B1(_02846_),
    .Y(_02862_));
 sky130_fd_sc_hd__a31o_1 _07322_ (.A1(\reg_pc[10] ),
    .A2(\decoded_imm[10] ),
    .A3(_02847_),
    .B1(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__inv_2 _07323_ (.A(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__xor2_1 _07324_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .X(_02865_));
 sky130_fd_sc_hd__inv_2 _07325_ (.A(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__a21o_1 _07326_ (.A1(_02860_),
    .A2(_02864_),
    .B1(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__or3b_1 _07327_ (.A(_02863_),
    .B(_02865_),
    .C_N(_02860_),
    .X(_02868_));
 sky130_fd_sc_hd__o221a_1 _07328_ (.A1(net21),
    .A2(_02689_),
    .B1(_02694_),
    .B2(net4),
    .C1(_02812_),
    .X(_02869_));
 sky130_fd_sc_hd__o21a_1 _07329_ (.A1(_02811_),
    .A2(_02869_),
    .B1(net1060),
    .X(_02870_));
 sky130_fd_sc_hd__a22o_1 _07330_ (.A1(\count_instr[44] ),
    .A2(net1131),
    .B1(net1136),
    .B2(\count_instr[12] ),
    .X(_02871_));
 sky130_fd_sc_hd__a211o_1 _07331_ (.A1(net1140),
    .A2(\count_cycle[44] ),
    .B1(net977),
    .C1(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__or2_1 _07332_ (.A(\count_cycle[12] ),
    .B(net972),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _07333_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[12] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[12] ),
    .S(net1110),
    .X(_02874_));
 sky130_fd_sc_hd__a221o_1 _07334_ (.A1(net1063),
    .A2(net1026),
    .B1(_02874_),
    .B2(net1077),
    .C1(_02870_),
    .X(_02875_));
 sky130_fd_sc_hd__a31o_1 _07335_ (.A1(net1071),
    .A2(_02867_),
    .A3(_02868_),
    .B1(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__a31o_2 _07336_ (.A1(net841),
    .A2(_02872_),
    .A3(_02873_),
    .B1(_02876_),
    .X(_06719_));
 sky130_fd_sc_hd__and2_1 _07337_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .X(_02877_));
 sky130_fd_sc_hd__nand2_1 _07338_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .Y(_02878_));
 sky130_fd_sc_hd__nor2_1 _07339_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .Y(_02879_));
 sky130_fd_sc_hd__nor2_1 _07340_ (.A(_02877_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__a21bo_1 _07341_ (.A1(\reg_pc[12] ),
    .A2(\decoded_imm[12] ),
    .B1_N(_02867_),
    .X(_02881_));
 sky130_fd_sc_hd__or2_1 _07342_ (.A(_02880_),
    .B(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(_02880_),
    .B(_02881_),
    .Y(_02883_));
 sky130_fd_sc_hd__o221a_1 _07344_ (.A1(net22),
    .A2(_02689_),
    .B1(_02694_),
    .B2(net5),
    .C1(_02812_),
    .X(_02884_));
 sky130_fd_sc_hd__o21a_1 _07345_ (.A1(_02811_),
    .A2(_02884_),
    .B1(net1060),
    .X(_02885_));
 sky130_fd_sc_hd__a22o_1 _07346_ (.A1(\count_instr[45] ),
    .A2(net1131),
    .B1(net1136),
    .B2(\count_instr[13] ),
    .X(_02886_));
 sky130_fd_sc_hd__a211o_1 _07347_ (.A1(net1140),
    .A2(\count_cycle[45] ),
    .B1(net977),
    .C1(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__o211a_1 _07348_ (.A1(\count_cycle[13] ),
    .A2(net971),
    .B1(net841),
    .C1(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _07349_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[13] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[13] ),
    .S(net1110),
    .X(_02889_));
 sky130_fd_sc_hd__a221o_1 _07350_ (.A1(net1063),
    .A2(net1024),
    .B1(_02889_),
    .B2(net1077),
    .C1(_02885_),
    .X(_02890_));
 sky130_fd_sc_hd__a31o_1 _07351_ (.A1(net1071),
    .A2(_02882_),
    .A3(_02883_),
    .B1(_02888_),
    .X(_02891_));
 sky130_fd_sc_hd__or2_1 _07352_ (.A(_02890_),
    .B(_02891_),
    .X(_06720_));
 sky130_fd_sc_hd__xor2_1 _07353_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .X(_02892_));
 sky130_fd_sc_hd__nand2b_1 _07354_ (.A_N(_02879_),
    .B(_02881_),
    .Y(_02893_));
 sky130_fd_sc_hd__a31o_1 _07355_ (.A1(\reg_pc[12] ),
    .A2(\decoded_imm[12] ),
    .A3(_02880_),
    .B1(_02877_),
    .X(_02894_));
 sky130_fd_sc_hd__a21bo_1 _07356_ (.A1(_02878_),
    .A2(_02893_),
    .B1_N(_02892_),
    .X(_02895_));
 sky130_fd_sc_hd__or3b_1 _07357_ (.A(_02877_),
    .B(_02892_),
    .C_N(_02893_),
    .X(_02896_));
 sky130_fd_sc_hd__o221a_1 _07358_ (.A1(net24),
    .A2(_02689_),
    .B1(_02694_),
    .B2(net6),
    .C1(_02812_),
    .X(_02897_));
 sky130_fd_sc_hd__o21a_1 _07359_ (.A1(_02811_),
    .A2(_02897_),
    .B1(net1060),
    .X(_02898_));
 sky130_fd_sc_hd__a22o_1 _07360_ (.A1(\count_instr[46] ),
    .A2(net1130),
    .B1(net1136),
    .B2(\count_instr[14] ),
    .X(_02899_));
 sky130_fd_sc_hd__a211o_1 _07361_ (.A1(net1140),
    .A2(\count_cycle[46] ),
    .B1(net977),
    .C1(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__o211a_1 _07362_ (.A1(\count_cycle[14] ),
    .A2(net971),
    .B1(net841),
    .C1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _07363_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[14] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[14] ),
    .S(net1110),
    .X(_02902_));
 sky130_fd_sc_hd__a221o_1 _07364_ (.A1(net1064),
    .A2(net1022),
    .B1(_02902_),
    .B2(net1079),
    .C1(_02901_),
    .X(_02903_));
 sky130_fd_sc_hd__or2_1 _07365_ (.A(_02898_),
    .B(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__a31o_1 _07366_ (.A1(net1071),
    .A2(_02895_),
    .A3(_02896_),
    .B1(_02904_),
    .X(_06721_));
 sky130_fd_sc_hd__or2_1 _07367_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .X(_02905_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(\reg_pc[15] ),
    .B(\decoded_imm[15] ),
    .Y(_02906_));
 sky130_fd_sc_hd__and2_1 _07369_ (.A(_02905_),
    .B(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__a21bo_1 _07370_ (.A1(\reg_pc[14] ),
    .A2(\decoded_imm[14] ),
    .B1_N(_02895_),
    .X(_02908_));
 sky130_fd_sc_hd__xor2_2 _07371_ (.A(_02907_),
    .B(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__or2_1 _07372_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .X(_02910_));
 sky130_fd_sc_hd__a21o_1 _07373_ (.A1(net1054),
    .A2(_02797_),
    .B1(net938),
    .X(_02911_));
 sky130_fd_sc_hd__o21a_1 _07374_ (.A1(net7),
    .A2(_02694_),
    .B1(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__a21oi_1 _07375_ (.A1(latched_is_lh),
    .A2(_02912_),
    .B1(_02811_),
    .Y(_02913_));
 sky130_fd_sc_hd__a21o_1 _07376_ (.A1(net936),
    .A2(_02913_),
    .B1(_02387_),
    .X(_02914_));
 sky130_fd_sc_hd__o21ba_1 _07377_ (.A1(net936),
    .A2(_02912_),
    .B1_N(net358),
    .X(_02915_));
 sky130_fd_sc_hd__a22o_1 _07378_ (.A1(\count_instr[47] ),
    .A2(net1132),
    .B1(net1140),
    .B2(\count_cycle[47] ),
    .X(_02916_));
 sky130_fd_sc_hd__a211o_1 _07379_ (.A1(\count_instr[15] ),
    .A2(net1136),
    .B1(net977),
    .C1(_02916_),
    .X(_02917_));
 sky130_fd_sc_hd__or2_1 _07380_ (.A(\count_cycle[15] ),
    .B(net971),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _07381_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[15] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[15] ),
    .S(net1110),
    .X(_02919_));
 sky130_fd_sc_hd__a221o_1 _07382_ (.A1(net1063),
    .A2(net1020),
    .B1(_02919_),
    .B2(net1078),
    .C1(_02915_),
    .X(_02920_));
 sky130_fd_sc_hd__a32o_1 _07383_ (.A1(net842),
    .A2(_02917_),
    .A3(_02918_),
    .B1(_02909_),
    .B2(net1071),
    .X(_02921_));
 sky130_fd_sc_hd__or2_1 _07384_ (.A(_02920_),
    .B(_02921_),
    .X(_06722_));
 sky130_fd_sc_hd__or2_1 _07385_ (.A(\reg_pc[16] ),
    .B(\decoded_imm[16] ),
    .X(_02922_));
 sky130_fd_sc_hd__nand2_1 _07386_ (.A(\reg_pc[16] ),
    .B(\decoded_imm[16] ),
    .Y(_02923_));
 sky130_fd_sc_hd__nand2_1 _07387_ (.A(_02922_),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand3_1 _07388_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .C(_02905_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand3_1 _07389_ (.A(_02880_),
    .B(_02892_),
    .C(_02907_),
    .Y(_02926_));
 sky130_fd_sc_hd__a211o_1 _07390_ (.A1(_02860_),
    .A2(_02864_),
    .B1(_02866_),
    .C1(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__nand3_1 _07391_ (.A(_02892_),
    .B(_02894_),
    .C(_02907_),
    .Y(_02928_));
 sky130_fd_sc_hd__and4_1 _07392_ (.A(_02906_),
    .B(_02925_),
    .C(_02927_),
    .D(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__or2_1 _07393_ (.A(_02924_),
    .B(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__nand2_1 _07394_ (.A(_02924_),
    .B(_02929_),
    .Y(_02931_));
 sky130_fd_sc_hd__a21oi_1 _07395_ (.A1(net8),
    .A2(net939),
    .B1(net936),
    .Y(_02932_));
 sky130_fd_sc_hd__a22o_1 _07396_ (.A1(\count_instr[48] ),
    .A2(net1132),
    .B1(net1140),
    .B2(\count_cycle[48] ),
    .X(_02933_));
 sky130_fd_sc_hd__a211o_1 _07397_ (.A1(\count_instr[16] ),
    .A2(net1136),
    .B1(net977),
    .C1(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__o211a_1 _07398_ (.A1(\count_cycle[16] ),
    .A2(net974),
    .B1(net844),
    .C1(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_1 _07399_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[16] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[16] ),
    .S(net1111),
    .X(_02936_));
 sky130_fd_sc_hd__a221o_1 _07400_ (.A1(net1065),
    .A2(net1018),
    .B1(_02936_),
    .B2(net1079),
    .C1(_02935_),
    .X(_02937_));
 sky130_fd_sc_hd__o21bai_2 _07401_ (.A1(net358),
    .A2(_02932_),
    .B1_N(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__a31o_1 _07402_ (.A1(net1071),
    .A2(_02930_),
    .A3(_02931_),
    .B1(_02938_),
    .X(_06723_));
 sky130_fd_sc_hd__nand2_1 _07403_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_02939_));
 sky130_fd_sc_hd__or2_1 _07404_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .X(_02940_));
 sky130_fd_sc_hd__nand2_1 _07405_ (.A(_02939_),
    .B(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__a21oi_1 _07406_ (.A1(_02923_),
    .A2(_02930_),
    .B1(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__a311o_1 _07407_ (.A1(_02923_),
    .A2(_02930_),
    .A3(_02941_),
    .B1(_02942_),
    .C1(net991),
    .X(_02943_));
 sky130_fd_sc_hd__a21oi_1 _07408_ (.A1(net9),
    .A2(net939),
    .B1(net936),
    .Y(_02944_));
 sky130_fd_sc_hd__nor2_1 _07409_ (.A(net358),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__a22o_1 _07410_ (.A1(\count_instr[49] ),
    .A2(net1132),
    .B1(net1140),
    .B2(\count_cycle[49] ),
    .X(_02946_));
 sky130_fd_sc_hd__a211o_1 _07411_ (.A1(\count_instr[17] ),
    .A2(net1136),
    .B1(net977),
    .C1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__o211a_1 _07412_ (.A1(\count_cycle[17] ),
    .A2(net974),
    .B1(net844),
    .C1(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _07413_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[17] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[17] ),
    .S(net1111),
    .X(_02949_));
 sky130_fd_sc_hd__a221o_1 _07414_ (.A1(net1065),
    .A2(net1016),
    .B1(_02949_),
    .B2(net1079),
    .C1(_02948_),
    .X(_02950_));
 sky130_fd_sc_hd__or3b_1 _07415_ (.A(_02950_),
    .B(_02945_),
    .C_N(_02943_),
    .X(_06724_));
 sky130_fd_sc_hd__nand2_1 _07416_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .Y(_02951_));
 sky130_fd_sc_hd__or2_1 _07417_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .X(_02952_));
 sky130_fd_sc_hd__nand2_1 _07418_ (.A(_02951_),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__o21ai_1 _07419_ (.A1(_02923_),
    .A2(_02941_),
    .B1(_02939_),
    .Y(_02954_));
 sky130_fd_sc_hd__and2b_1 _07420_ (.A_N(_02942_),
    .B(_02939_),
    .X(_02955_));
 sky130_fd_sc_hd__or2_1 _07421_ (.A(_02953_),
    .B(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__nand2_1 _07422_ (.A(_02953_),
    .B(_02955_),
    .Y(_02957_));
 sky130_fd_sc_hd__a21oi_1 _07423_ (.A1(net10),
    .A2(net939),
    .B1(net936),
    .Y(_02958_));
 sky130_fd_sc_hd__a22o_1 _07424_ (.A1(\count_instr[50] ),
    .A2(net1132),
    .B1(net1140),
    .B2(\count_cycle[50] ),
    .X(_02959_));
 sky130_fd_sc_hd__a211o_1 _07425_ (.A1(\count_instr[18] ),
    .A2(net1136),
    .B1(net977),
    .C1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__o211a_1 _07426_ (.A1(\count_cycle[18] ),
    .A2(net974),
    .B1(net844),
    .C1(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _07427_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[18] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[18] ),
    .S(net1111),
    .X(_02962_));
 sky130_fd_sc_hd__a221o_1 _07428_ (.A1(net1065),
    .A2(net1014),
    .B1(_02962_),
    .B2(net1079),
    .C1(_02961_),
    .X(_02963_));
 sky130_fd_sc_hd__o21bai_1 _07429_ (.A1(net358),
    .A2(_02958_),
    .B1_N(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__a31o_1 _07430_ (.A1(net1074),
    .A2(_02956_),
    .A3(_02957_),
    .B1(_02964_),
    .X(_06725_));
 sky130_fd_sc_hd__xnor2_1 _07431_ (.A(\reg_pc[19] ),
    .B(\decoded_imm[19] ),
    .Y(_02965_));
 sky130_fd_sc_hd__nand3_1 _07432_ (.A(_02951_),
    .B(_02956_),
    .C(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__a21o_1 _07433_ (.A1(_02951_),
    .A2(_02956_),
    .B1(_02965_),
    .X(_02967_));
 sky130_fd_sc_hd__a21oi_1 _07434_ (.A1(net11),
    .A2(net939),
    .B1(net936),
    .Y(_02968_));
 sky130_fd_sc_hd__a22o_1 _07435_ (.A1(\count_instr[51] ),
    .A2(net1132),
    .B1(net1142),
    .B2(\count_cycle[51] ),
    .X(_02969_));
 sky130_fd_sc_hd__a211o_1 _07436_ (.A1(\count_instr[19] ),
    .A2(net1138),
    .B1(net978),
    .C1(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__o211a_1 _07437_ (.A1(\count_cycle[19] ),
    .A2(net973),
    .B1(net843),
    .C1(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _07438_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[19] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[19] ),
    .S(net1111),
    .X(_02972_));
 sky130_fd_sc_hd__a221o_1 _07439_ (.A1(net1065),
    .A2(net1012),
    .B1(_02972_),
    .B2(net1078),
    .C1(_02971_),
    .X(_02973_));
 sky130_fd_sc_hd__o21bai_1 _07440_ (.A1(net358),
    .A2(_02968_),
    .B1_N(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__a31o_1 _07441_ (.A1(net1074),
    .A2(_02966_),
    .A3(_02967_),
    .B1(_02974_),
    .X(_06726_));
 sky130_fd_sc_hd__or2_1 _07442_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .X(_02975_));
 sky130_fd_sc_hd__nand2_1 _07443_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .Y(_02976_));
 sky130_fd_sc_hd__and2_1 _07444_ (.A(_02975_),
    .B(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__nor2_1 _07445_ (.A(_02953_),
    .B(_02965_),
    .Y(_02978_));
 sky130_fd_sc_hd__o211a_1 _07446_ (.A1(\reg_pc[19] ),
    .A2(\decoded_imm[19] ),
    .B1(\decoded_imm[18] ),
    .C1(\reg_pc[18] ),
    .X(_02979_));
 sky130_fd_sc_hd__a221o_1 _07447_ (.A1(\reg_pc[19] ),
    .A2(\decoded_imm[19] ),
    .B1(_02954_),
    .B2(_02978_),
    .C1(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__inv_2 _07448_ (.A(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__o41a_1 _07449_ (.A1(_02930_),
    .A2(_02941_),
    .A3(_02953_),
    .A4(_02965_),
    .B1(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__nand2b_1 _07450_ (.A_N(_02982_),
    .B(_02977_),
    .Y(_02983_));
 sky130_fd_sc_hd__xnor2_1 _07451_ (.A(_02977_),
    .B(_02982_),
    .Y(_02984_));
 sky130_fd_sc_hd__a21oi_1 _07452_ (.A1(net13),
    .A2(net939),
    .B1(net936),
    .Y(_02985_));
 sky130_fd_sc_hd__a22o_1 _07453_ (.A1(\count_instr[20] ),
    .A2(net1138),
    .B1(\count_cycle[52] ),
    .B2(net1142),
    .X(_02986_));
 sky130_fd_sc_hd__a211o_1 _07454_ (.A1(\count_instr[52] ),
    .A2(net1134),
    .B1(net978),
    .C1(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__o211a_1 _07455_ (.A1(\count_cycle[20] ),
    .A2(net974),
    .B1(net844),
    .C1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _07456_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[20] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[20] ),
    .S(net1112),
    .X(_02989_));
 sky130_fd_sc_hd__a221o_1 _07457_ (.A1(net1067),
    .A2(net1010),
    .B1(_02989_),
    .B2(net1086),
    .C1(_02988_),
    .X(_02990_));
 sky130_fd_sc_hd__o21bai_1 _07458_ (.A1(net358),
    .A2(_02985_),
    .B1_N(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__a21o_1 _07459_ (.A1(net1073),
    .A2(_02984_),
    .B1(_02991_),
    .X(_06728_));
 sky130_fd_sc_hd__or2_1 _07460_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .X(_02992_));
 sky130_fd_sc_hd__nand2_1 _07461_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .Y(_02993_));
 sky130_fd_sc_hd__and2_1 _07462_ (.A(_02992_),
    .B(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__nand2_1 _07463_ (.A(_02992_),
    .B(_02993_),
    .Y(_02995_));
 sky130_fd_sc_hd__nand2_1 _07464_ (.A(_02976_),
    .B(_02983_),
    .Y(_02996_));
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(_02994_),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__o211a_1 _07466_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_02997_),
    .C1(net1073),
    .X(_02998_));
 sky130_fd_sc_hd__a21oi_1 _07467_ (.A1(net14),
    .A2(net938),
    .B1(net936),
    .Y(_02999_));
 sky130_fd_sc_hd__nor2_1 _07468_ (.A(net358),
    .B(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__a22o_1 _07469_ (.A1(\count_instr[53] ),
    .A2(net1134),
    .B1(net1142),
    .B2(\count_cycle[53] ),
    .X(_03001_));
 sky130_fd_sc_hd__a211o_1 _07470_ (.A1(\count_instr[21] ),
    .A2(net1138),
    .B1(net978),
    .C1(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__o211a_1 _07471_ (.A1(\count_cycle[21] ),
    .A2(net973),
    .B1(net844),
    .C1(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__mux2_1 _07472_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[21] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[21] ),
    .S(net1112),
    .X(_03004_));
 sky130_fd_sc_hd__a221o_1 _07473_ (.A1(net1066),
    .A2(net1009),
    .B1(_03004_),
    .B2(net1086),
    .C1(_03003_),
    .X(_03005_));
 sky130_fd_sc_hd__or3_1 _07474_ (.A(_02998_),
    .B(_03000_),
    .C(_03005_),
    .X(_06729_));
 sky130_fd_sc_hd__or2_1 _07475_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .X(_03006_));
 sky130_fd_sc_hd__nand2_1 _07476_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _07477_ (.A(_03006_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__o21a_1 _07478_ (.A1(_02976_),
    .A2(_02995_),
    .B1(_02993_),
    .X(_03009_));
 sky130_fd_sc_hd__a21o_1 _07479_ (.A1(_02993_),
    .A2(_02997_),
    .B1(_03008_),
    .X(_03010_));
 sky130_fd_sc_hd__nand3_1 _07480_ (.A(_02993_),
    .B(_02997_),
    .C(_03008_),
    .Y(_03011_));
 sky130_fd_sc_hd__a21oi_1 _07481_ (.A1(net15),
    .A2(net938),
    .B1(net936),
    .Y(_03012_));
 sky130_fd_sc_hd__a22o_1 _07482_ (.A1(\count_instr[54] ),
    .A2(net1133),
    .B1(net1141),
    .B2(\count_cycle[54] ),
    .X(_03013_));
 sky130_fd_sc_hd__a211o_1 _07483_ (.A1(\count_instr[22] ),
    .A2(net1137),
    .B1(net978),
    .C1(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__o211a_1 _07484_ (.A1(\count_cycle[22] ),
    .A2(net973),
    .B1(net843),
    .C1(_03014_),
    .X(_03015_));
 sky130_fd_sc_hd__mux2_1 _07485_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[22] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[22] ),
    .S(net1112),
    .X(_03016_));
 sky130_fd_sc_hd__a221o_1 _07486_ (.A1(net1067),
    .A2(net1007),
    .B1(_03016_),
    .B2(net1082),
    .C1(_03015_),
    .X(_03017_));
 sky130_fd_sc_hd__o21bai_1 _07487_ (.A1(net358),
    .A2(_03012_),
    .B1_N(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__a31o_1 _07488_ (.A1(net1073),
    .A2(_03010_),
    .A3(_03011_),
    .B1(_03018_),
    .X(_06730_));
 sky130_fd_sc_hd__nor2_1 _07489_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .Y(_03019_));
 sky130_fd_sc_hd__nand2_1 _07490_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .Y(_03020_));
 sky130_fd_sc_hd__nand2b_1 _07491_ (.A_N(_03019_),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__nand3_1 _07492_ (.A(_03007_),
    .B(_03010_),
    .C(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__a21o_1 _07493_ (.A1(_03007_),
    .A2(_03010_),
    .B1(_03021_),
    .X(_03023_));
 sky130_fd_sc_hd__a21oi_1 _07494_ (.A1(net16),
    .A2(net938),
    .B1(net936),
    .Y(_03024_));
 sky130_fd_sc_hd__a22o_1 _07495_ (.A1(\count_instr[55] ),
    .A2(net1133),
    .B1(net1141),
    .B2(\count_cycle[55] ),
    .X(_03025_));
 sky130_fd_sc_hd__a211o_1 _07496_ (.A1(\count_instr[23] ),
    .A2(net1137),
    .B1(net979),
    .C1(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__o211a_1 _07497_ (.A1(\count_cycle[23] ),
    .A2(net973),
    .B1(net843),
    .C1(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _07498_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[23] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[23] ),
    .S(net1112),
    .X(_03028_));
 sky130_fd_sc_hd__a221o_1 _07499_ (.A1(net1067),
    .A2(net1006),
    .B1(_03028_),
    .B2(net1082),
    .C1(_03027_),
    .X(_03029_));
 sky130_fd_sc_hd__o21bai_1 _07500_ (.A1(net358),
    .A2(_03024_),
    .B1_N(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__a31o_1 _07501_ (.A1(net1073),
    .A2(_03022_),
    .A3(_03023_),
    .B1(_03030_),
    .X(_06731_));
 sky130_fd_sc_hd__or2_1 _07502_ (.A(_03008_),
    .B(_03021_),
    .X(_03031_));
 sky130_fd_sc_hd__o221a_1 _07503_ (.A1(_03007_),
    .A2(_03019_),
    .B1(_03031_),
    .B2(_03009_),
    .C1(_03020_),
    .X(_03032_));
 sky130_fd_sc_hd__o31a_1 _07504_ (.A1(_02983_),
    .A2(_02995_),
    .A3(_03031_),
    .B1(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__or2_1 _07505_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .X(_03034_));
 sky130_fd_sc_hd__nand2_1 _07506_ (.A(\reg_pc[24] ),
    .B(\decoded_imm[24] ),
    .Y(_03035_));
 sky130_fd_sc_hd__nand2_1 _07507_ (.A(_03034_),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__or2_1 _07508_ (.A(_03033_),
    .B(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__nand2_1 _07509_ (.A(_03033_),
    .B(_03036_),
    .Y(_03038_));
 sky130_fd_sc_hd__a21oi_1 _07510_ (.A1(net17),
    .A2(net938),
    .B1(net937),
    .Y(_03039_));
 sky130_fd_sc_hd__a22o_1 _07511_ (.A1(\count_instr[56] ),
    .A2(net1133),
    .B1(net1137),
    .B2(\count_instr[24] ),
    .X(_03040_));
 sky130_fd_sc_hd__a211o_1 _07512_ (.A1(net1141),
    .A2(\count_cycle[56] ),
    .B1(net979),
    .C1(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__o211a_1 _07513_ (.A1(\count_cycle[24] ),
    .A2(net973),
    .B1(net843),
    .C1(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _07514_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[24] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[24] ),
    .S(net1112),
    .X(_03043_));
 sky130_fd_sc_hd__a221o_1 _07515_ (.A1(net1067),
    .A2(net1005),
    .B1(_03043_),
    .B2(net1082),
    .C1(_03042_),
    .X(_03044_));
 sky130_fd_sc_hd__o21bai_1 _07516_ (.A1(net358),
    .A2(_03039_),
    .B1_N(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__a31o_1 _07517_ (.A1(net1073),
    .A2(_03037_),
    .A3(_03038_),
    .B1(_03045_),
    .X(_06732_));
 sky130_fd_sc_hd__nor2_1 _07518_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_03046_));
 sky130_fd_sc_hd__nand2_1 _07519_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_03047_));
 sky130_fd_sc_hd__nand2b_1 _07520_ (.A_N(_03046_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__a21o_1 _07521_ (.A1(_03035_),
    .A2(_03037_),
    .B1(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__nand3_1 _07522_ (.A(_03035_),
    .B(_03037_),
    .C(_03048_),
    .Y(_03050_));
 sky130_fd_sc_hd__a21oi_1 _07523_ (.A1(net18),
    .A2(net938),
    .B1(net937),
    .Y(_03051_));
 sky130_fd_sc_hd__a22o_1 _07524_ (.A1(\count_instr[57] ),
    .A2(net1133),
    .B1(net1141),
    .B2(\count_cycle[57] ),
    .X(_03052_));
 sky130_fd_sc_hd__a211o_1 _07525_ (.A1(\count_instr[25] ),
    .A2(net1137),
    .B1(net979),
    .C1(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__o211a_1 _07526_ (.A1(\count_cycle[25] ),
    .A2(net973),
    .B1(net843),
    .C1(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__mux2_1 _07527_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[25] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[25] ),
    .S(net1113),
    .X(_03055_));
 sky130_fd_sc_hd__a221o_1 _07528_ (.A1(net1069),
    .A2(net1003),
    .B1(_03055_),
    .B2(net1085),
    .C1(_03054_),
    .X(_03056_));
 sky130_fd_sc_hd__o21bai_1 _07529_ (.A1(net359),
    .A2(_03051_),
    .B1_N(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__a31o_1 _07530_ (.A1(net1073),
    .A2(_03049_),
    .A3(_03050_),
    .B1(_03057_),
    .X(_06733_));
 sky130_fd_sc_hd__nand2_1 _07531_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .Y(_03058_));
 sky130_fd_sc_hd__or2_1 _07532_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .X(_03059_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(_03058_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__a21o_1 _07534_ (.A1(_03047_),
    .A2(_03049_),
    .B1(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__nand3_1 _07535_ (.A(_03047_),
    .B(_03049_),
    .C(_03060_),
    .Y(_03062_));
 sky130_fd_sc_hd__a21oi_1 _07536_ (.A1(net19),
    .A2(net938),
    .B1(net937),
    .Y(_03063_));
 sky130_fd_sc_hd__nor2_1 _07537_ (.A(net359),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__mux2_1 _07538_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[26] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[26] ),
    .S(net1113),
    .X(_03065_));
 sky130_fd_sc_hd__a22o_1 _07539_ (.A1(net1069),
    .A2(net1000),
    .B1(_03065_),
    .B2(net1085),
    .X(_03066_));
 sky130_fd_sc_hd__or2_1 _07540_ (.A(_02702_),
    .B(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__a31o_1 _07541_ (.A1(net1073),
    .A2(_03061_),
    .A3(_03062_),
    .B1(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__a22o_1 _07542_ (.A1(\count_instr[58] ),
    .A2(net1133),
    .B1(net1137),
    .B2(\count_instr[26] ),
    .X(_03069_));
 sky130_fd_sc_hd__a221o_1 _07543_ (.A1(net1142),
    .A2(\count_cycle[58] ),
    .B1(\count_cycle[26] ),
    .B2(net978),
    .C1(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__o22a_1 _07544_ (.A1(_03064_),
    .A2(_03068_),
    .B1(_03070_),
    .B2(_02703_),
    .X(_06734_));
 sky130_fd_sc_hd__nor2_1 _07545_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_03071_));
 sky130_fd_sc_hd__nand2_1 _07546_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_03072_));
 sky130_fd_sc_hd__nand2b_1 _07547_ (.A_N(_03071_),
    .B(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__nand3_1 _07548_ (.A(_03058_),
    .B(_03061_),
    .C(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__a21o_1 _07549_ (.A1(_03058_),
    .A2(_03061_),
    .B1(_03073_),
    .X(_03075_));
 sky130_fd_sc_hd__a21oi_1 _07550_ (.A1(net20),
    .A2(net938),
    .B1(net937),
    .Y(_03076_));
 sky130_fd_sc_hd__a22o_1 _07551_ (.A1(\count_instr[59] ),
    .A2(net1133),
    .B1(net1141),
    .B2(\count_cycle[59] ),
    .X(_03077_));
 sky130_fd_sc_hd__a211o_1 _07552_ (.A1(\count_instr[27] ),
    .A2(net1138),
    .B1(net978),
    .C1(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__o211a_1 _07553_ (.A1(\count_cycle[27] ),
    .A2(net973),
    .B1(net843),
    .C1(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_1 _07554_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[27] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[27] ),
    .S(net1113),
    .X(_03080_));
 sky130_fd_sc_hd__a221o_1 _07555_ (.A1(net1069),
    .A2(net999),
    .B1(_03080_),
    .B2(net1085),
    .C1(_03079_),
    .X(_03081_));
 sky130_fd_sc_hd__o21bai_1 _07556_ (.A1(net359),
    .A2(_03076_),
    .B1_N(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__a31o_1 _07557_ (.A1(net1072),
    .A2(_03074_),
    .A3(_03075_),
    .B1(_03082_),
    .X(_06735_));
 sky130_fd_sc_hd__or2_1 _07558_ (.A(_03060_),
    .B(_03073_),
    .X(_03083_));
 sky130_fd_sc_hd__o21a_1 _07559_ (.A1(_03035_),
    .A2(_03046_),
    .B1(_03047_),
    .X(_03084_));
 sky130_fd_sc_hd__o221a_1 _07560_ (.A1(_03058_),
    .A2(_03071_),
    .B1(_03083_),
    .B2(_03084_),
    .C1(_03072_),
    .X(_03085_));
 sky130_fd_sc_hd__o31a_1 _07561_ (.A1(_03037_),
    .A2(_03048_),
    .A3(_03083_),
    .B1(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__or2_1 _07562_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .X(_03087_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_03088_));
 sky130_fd_sc_hd__nand2_1 _07564_ (.A(_03087_),
    .B(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__or2_1 _07565_ (.A(_03086_),
    .B(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__nand2_1 _07566_ (.A(_03086_),
    .B(_03089_),
    .Y(_03091_));
 sky130_fd_sc_hd__a21oi_1 _07567_ (.A1(net21),
    .A2(net939),
    .B1(net937),
    .Y(_03092_));
 sky130_fd_sc_hd__a22o_1 _07568_ (.A1(\count_instr[60] ),
    .A2(net1134),
    .B1(net1141),
    .B2(\count_cycle[60] ),
    .X(_03093_));
 sky130_fd_sc_hd__a211o_1 _07569_ (.A1(\count_instr[28] ),
    .A2(net1137),
    .B1(net978),
    .C1(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__o211a_1 _07570_ (.A1(\count_cycle[28] ),
    .A2(net973),
    .B1(net843),
    .C1(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__mux2_1 _07571_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[28] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[28] ),
    .S(net1112),
    .X(_03096_));
 sky130_fd_sc_hd__a221o_1 _07572_ (.A1(net1068),
    .A2(net996),
    .B1(_03096_),
    .B2(net1085),
    .C1(_03095_),
    .X(_03097_));
 sky130_fd_sc_hd__o21bai_1 _07573_ (.A1(net359),
    .A2(_03092_),
    .B1_N(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__a31o_1 _07574_ (.A1(net1072),
    .A2(_03090_),
    .A3(_03091_),
    .B1(_03098_),
    .X(_06736_));
 sky130_fd_sc_hd__nor2_1 _07575_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .Y(_03099_));
 sky130_fd_sc_hd__and2_1 _07576_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .X(_03100_));
 sky130_fd_sc_hd__o21ai_1 _07577_ (.A1(_03086_),
    .A2(_03089_),
    .B1(_03088_),
    .Y(_03101_));
 sky130_fd_sc_hd__o21bai_1 _07578_ (.A1(_03099_),
    .A2(_03100_),
    .B1_N(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__or3b_1 _07579_ (.A(_03099_),
    .B(_03100_),
    .C_N(_03101_),
    .X(_03103_));
 sky130_fd_sc_hd__a21oi_1 _07580_ (.A1(net22),
    .A2(net938),
    .B1(net937),
    .Y(_03104_));
 sky130_fd_sc_hd__nor2_1 _07581_ (.A(net359),
    .B(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__a22o_1 _07582_ (.A1(\count_instr[61] ),
    .A2(net1133),
    .B1(net1137),
    .B2(\count_instr[29] ),
    .X(_03106_));
 sky130_fd_sc_hd__a211o_1 _07583_ (.A1(net1141),
    .A2(\count_cycle[61] ),
    .B1(net978),
    .C1(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__o211a_1 _07584_ (.A1(\count_cycle[29] ),
    .A2(net973),
    .B1(net843),
    .C1(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__mux2_1 _07585_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[29] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[29] ),
    .S(net1113),
    .X(_03109_));
 sky130_fd_sc_hd__a221o_1 _07586_ (.A1(net1068),
    .A2(net994),
    .B1(_03109_),
    .B2(net1084),
    .C1(_03105_),
    .X(_03110_));
 sky130_fd_sc_hd__a31o_1 _07587_ (.A1(net1072),
    .A2(_03102_),
    .A3(_03103_),
    .B1(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__or2_1 _07588_ (.A(_03108_),
    .B(_03111_),
    .X(_06737_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .Y(_03112_));
 sky130_fd_sc_hd__or2_1 _07590_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .X(_03113_));
 sky130_fd_sc_hd__and2b_1 _07591_ (.A_N(_03099_),
    .B(_03101_),
    .X(_03114_));
 sky130_fd_sc_hd__o211a_1 _07592_ (.A1(_03100_),
    .A2(_03114_),
    .B1(_03113_),
    .C1(_03112_),
    .X(_03115_));
 sky130_fd_sc_hd__a211o_1 _07593_ (.A1(_03112_),
    .A2(_03113_),
    .B1(_03114_),
    .C1(_03100_),
    .X(_03116_));
 sky130_fd_sc_hd__and3b_1 _07594_ (.A_N(_03115_),
    .B(_03116_),
    .C(net1072),
    .X(_03117_));
 sky130_fd_sc_hd__a21oi_1 _07595_ (.A1(net24),
    .A2(net939),
    .B1(net937),
    .Y(_03118_));
 sky130_fd_sc_hd__nor2_1 _07596_ (.A(net359),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__a22o_1 _07597_ (.A1(\count_instr[62] ),
    .A2(net1133),
    .B1(net1141),
    .B2(\count_cycle[62] ),
    .X(_03120_));
 sky130_fd_sc_hd__a211o_1 _07598_ (.A1(\count_instr[30] ),
    .A2(net1137),
    .B1(net978),
    .C1(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__o211a_1 _07599_ (.A1(\count_cycle[30] ),
    .A2(net974),
    .B1(net843),
    .C1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_1 _07600_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[30] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[30] ),
    .S(net1112),
    .X(_03123_));
 sky130_fd_sc_hd__a221o_1 _07601_ (.A1(net1069),
    .A2(net992),
    .B1(_03123_),
    .B2(net1085),
    .C1(_03122_),
    .X(_03124_));
 sky130_fd_sc_hd__or3_1 _07602_ (.A(_03117_),
    .B(_03119_),
    .C(_03124_),
    .X(_06739_));
 sky130_fd_sc_hd__a21oi_1 _07603_ (.A1(\reg_pc[30] ),
    .A2(\decoded_imm[30] ),
    .B1(_03115_),
    .Y(_03125_));
 sky130_fd_sc_hd__xnor2_1 _07604_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_03126_));
 sky130_fd_sc_hd__xnor2_1 _07605_ (.A(_03125_),
    .B(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__a21oi_1 _07606_ (.A1(net25),
    .A2(net939),
    .B1(net937),
    .Y(_03128_));
 sky130_fd_sc_hd__a22o_1 _07607_ (.A1(\count_instr[63] ),
    .A2(net1133),
    .B1(net1141),
    .B2(\count_cycle[63] ),
    .X(_03129_));
 sky130_fd_sc_hd__a211o_1 _07608_ (.A1(\count_instr[31] ),
    .A2(net1137),
    .B1(net978),
    .C1(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__o211a_1 _07609_ (.A1(\count_cycle[31] ),
    .A2(net973),
    .B1(net843),
    .C1(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__mux2_1 _07610_ (.A0(\genblk1.genblk1.pcpi_mul.pcpi_rd[31] ),
    .A1(\genblk2.pcpi_div.pcpi_rd[31] ),
    .S(net1112),
    .X(_03132_));
 sky130_fd_sc_hd__a221o_1 _07611_ (.A1(net1188),
    .A2(net1069),
    .B1(_03132_),
    .B2(net1085),
    .C1(_03131_),
    .X(_03133_));
 sky130_fd_sc_hd__o21ba_1 _07612_ (.A1(net359),
    .A2(_03128_),
    .B1_N(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__o21ai_1 _07613_ (.A1(net991),
    .A2(_03127_),
    .B1(_03134_),
    .Y(_06740_));
 sky130_fd_sc_hd__or2_1 _07614_ (.A(net1080),
    .B(\decoded_imm_j[17] ),
    .X(_03135_));
 sky130_fd_sc_hd__o21ai_2 _07615_ (.A1(net986),
    .A2(\decoded_imm_j[2] ),
    .B1(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__o21a_2 _07616_ (.A1(net986),
    .A2(\decoded_imm_j[2] ),
    .B1(_03135_),
    .X(_03137_));
 sky130_fd_sc_hd__or2_1 _07617_ (.A(net986),
    .B(\decoded_imm_j[11] ),
    .X(_03138_));
 sky130_fd_sc_hd__o21a_1 _07618_ (.A1(net1080),
    .A2(\decoded_imm_j[15] ),
    .B1(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__o21ai_1 _07619_ (.A1(net1080),
    .A2(\decoded_imm_j[15] ),
    .B1(_03138_),
    .Y(_03140_));
 sky130_fd_sc_hd__or2_1 _07620_ (.A(net1080),
    .B(\decoded_imm_j[16] ),
    .X(_03141_));
 sky130_fd_sc_hd__o21ai_1 _07621_ (.A1(net986),
    .A2(\decoded_imm_j[1] ),
    .B1(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__o21a_2 _07622_ (.A1(net986),
    .A2(\decoded_imm_j[1] ),
    .B1(_03141_),
    .X(_03143_));
 sky130_fd_sc_hd__mux2_1 _07623_ (.A0(\cpuregs[6][2] ),
    .A1(\cpuregs[7][2] ),
    .S(net700),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_1 _07624_ (.A0(\cpuregs[4][2] ),
    .A1(\cpuregs[5][2] ),
    .S(net700),
    .X(_03145_));
 sky130_fd_sc_hd__mux2_1 _07625_ (.A0(_03144_),
    .A1(_03145_),
    .S(net819),
    .X(_03146_));
 sky130_fd_sc_hd__or2_1 _07626_ (.A(\cpuregs[0][2] ),
    .B(net700),
    .X(_03147_));
 sky130_fd_sc_hd__nor2_4 _07627_ (.A(net822),
    .B(net796),
    .Y(_03148_));
 sky130_fd_sc_hd__o211a_1 _07628_ (.A1(\cpuregs[1][2] ),
    .A2(net641),
    .B1(_03147_),
    .C1(net614),
    .X(_03149_));
 sky130_fd_sc_hd__or2_1 _07629_ (.A(net1080),
    .B(\decoded_imm_j[18] ),
    .X(_03150_));
 sky130_fd_sc_hd__o21ai_1 _07630_ (.A1(net986),
    .A2(\decoded_imm_j[3] ),
    .B1(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__o21a_2 _07631_ (.A1(net986),
    .A2(\decoded_imm_j[3] ),
    .B1(_03150_),
    .X(_03152_));
 sky130_fd_sc_hd__nor2_2 _07632_ (.A(net824),
    .B(net810),
    .Y(_03153_));
 sky130_fd_sc_hd__or2_1 _07633_ (.A(\cpuregs[2][2] ),
    .B(net699),
    .X(_03154_));
 sky130_fd_sc_hd__o211a_1 _07634_ (.A1(\cpuregs[3][2] ),
    .A2(net640),
    .B1(net601),
    .C1(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__nand2_4 _07635_ (.A(net623),
    .B(net788),
    .Y(_03156_));
 sky130_fd_sc_hd__or3_1 _07636_ (.A(_03149_),
    .B(net785),
    .C(_03155_),
    .X(_03157_));
 sky130_fd_sc_hd__a21o_1 _07637_ (.A1(net835),
    .A2(_03146_),
    .B1(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__mux2_1 _07638_ (.A0(\cpuregs[12][2] ),
    .A1(\cpuregs[13][2] ),
    .S(net700),
    .X(_03159_));
 sky130_fd_sc_hd__mux2_1 _07639_ (.A0(\cpuregs[14][2] ),
    .A1(\cpuregs[15][2] ),
    .S(net700),
    .X(_03160_));
 sky130_fd_sc_hd__or2_1 _07640_ (.A(net819),
    .B(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__o211a_1 _07641_ (.A1(net807),
    .A2(_03159_),
    .B1(_03161_),
    .C1(net835),
    .X(_03162_));
 sky130_fd_sc_hd__or2_1 _07642_ (.A(\cpuregs[8][2] ),
    .B(net700),
    .X(_03163_));
 sky130_fd_sc_hd__o211a_1 _07643_ (.A1(\cpuregs[9][2] ),
    .A2(net640),
    .B1(net614),
    .C1(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__or2_1 _07644_ (.A(\cpuregs[10][2] ),
    .B(net699),
    .X(_03165_));
 sky130_fd_sc_hd__o211a_1 _07645_ (.A1(\cpuregs[11][2] ),
    .A2(net640),
    .B1(net601),
    .C1(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__or3_1 _07646_ (.A(net794),
    .B(_03164_),
    .C(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__or2_1 _07647_ (.A(net1080),
    .B(\decoded_imm_j[19] ),
    .X(_03168_));
 sky130_fd_sc_hd__o21ai_1 _07648_ (.A1(net986),
    .A2(\decoded_imm_j[4] ),
    .B1(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__o21a_2 _07649_ (.A1(net986),
    .A2(\decoded_imm_j[4] ),
    .B1(_03168_),
    .X(_03170_));
 sky130_fd_sc_hd__o31a_4 _07650_ (.A1(net825),
    .A2(net799),
    .A3(net552),
    .B1(net776),
    .X(_03171_));
 sky130_fd_sc_hd__o211a_1 _07651_ (.A1(_03162_),
    .A2(_03167_),
    .B1(_03171_),
    .C1(_03158_),
    .X(_03172_));
 sky130_fd_sc_hd__mux2_1 _07652_ (.A0(\cpuregs[20][2] ),
    .A1(\cpuregs[21][2] ),
    .S(net697),
    .X(_03173_));
 sky130_fd_sc_hd__mux2_1 _07653_ (.A0(\cpuregs[22][2] ),
    .A1(\cpuregs[23][2] ),
    .S(net701),
    .X(_03174_));
 sky130_fd_sc_hd__mux2_1 _07654_ (.A0(_03173_),
    .A1(_03174_),
    .S(net807),
    .X(_03175_));
 sky130_fd_sc_hd__or2_1 _07655_ (.A(\cpuregs[16][2] ),
    .B(net699),
    .X(_03176_));
 sky130_fd_sc_hd__o211a_1 _07656_ (.A1(\cpuregs[17][2] ),
    .A2(net641),
    .B1(net614),
    .C1(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__o21a_1 _07657_ (.A1(\cpuregs[19][2] ),
    .A2(net641),
    .B1(net601),
    .X(_03178_));
 sky130_fd_sc_hd__o22a_1 _07658_ (.A1(\cpuregs[18][2] ),
    .A2(net555),
    .B1(_03178_),
    .B2(net785),
    .X(_03179_));
 sky130_fd_sc_hd__a211o_1 _07659_ (.A1(net837),
    .A2(_03175_),
    .B1(_03177_),
    .C1(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_1 _07660_ (.A0(\cpuregs[28][2] ),
    .A1(\cpuregs[29][2] ),
    .S(net701),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _07661_ (.A0(\cpuregs[30][2] ),
    .A1(\cpuregs[31][2] ),
    .S(net701),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_1 _07662_ (.A0(_03181_),
    .A1(_03182_),
    .S(net807),
    .X(_03183_));
 sky130_fd_sc_hd__or2_1 _07663_ (.A(\cpuregs[24][2] ),
    .B(net700),
    .X(_03184_));
 sky130_fd_sc_hd__o211a_1 _07664_ (.A1(\cpuregs[25][2] ),
    .A2(net641),
    .B1(net614),
    .C1(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__or2_1 _07665_ (.A(\cpuregs[26][2] ),
    .B(net700),
    .X(_03186_));
 sky130_fd_sc_hd__o211a_1 _07666_ (.A1(\cpuregs[27][2] ),
    .A2(net641),
    .B1(net601),
    .C1(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__a2111o_1 _07667_ (.A1(net837),
    .A2(_03183_),
    .B1(_03185_),
    .C1(_03187_),
    .D1(net794),
    .X(_03188_));
 sky130_fd_sc_hd__a31o_1 _07668_ (.A1(net775),
    .A2(_03180_),
    .A3(_03188_),
    .B1(_03172_),
    .X(_03189_));
 sky130_fd_sc_hd__and2_1 _07669_ (.A(net1080),
    .B(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__o21ai_1 _07670_ (.A1(_02475_),
    .A2(_02476_),
    .B1(net1066),
    .Y(_03191_));
 sky130_fd_sc_hd__inv_2 _07671_ (.A(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__a221o_1 _07672_ (.A1(\decoded_imm_j[2] ),
    .A2(_02701_),
    .B1(_03192_),
    .B2(_02386_),
    .C1(_03190_),
    .X(_06748_));
 sky130_fd_sc_hd__mux2_1 _07673_ (.A0(\cpuregs[6][3] ),
    .A1(\cpuregs[7][3] ),
    .S(net662),
    .X(_03193_));
 sky130_fd_sc_hd__or2_1 _07674_ (.A(\cpuregs[4][3] ),
    .B(net662),
    .X(_03194_));
 sky130_fd_sc_hd__o211a_1 _07675_ (.A1(\cpuregs[5][3] ),
    .A2(net623),
    .B1(net811),
    .C1(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__a211o_1 _07676_ (.A1(net801),
    .A2(_03193_),
    .B1(_03195_),
    .C1(net838),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_1 _07677_ (.A0(\cpuregs[2][3] ),
    .A1(\cpuregs[3][3] ),
    .S(net675),
    .X(_03197_));
 sky130_fd_sc_hd__nor2_1 _07678_ (.A(net618),
    .B(net796),
    .Y(_03198_));
 sky130_fd_sc_hd__a221o_1 _07679_ (.A1(net801),
    .A2(_03197_),
    .B1(net549),
    .B2(\cpuregs[1][3] ),
    .C1(net829),
    .X(_03199_));
 sky130_fd_sc_hd__a21o_1 _07680_ (.A1(_03196_),
    .A2(_03199_),
    .B1(net781),
    .X(_03200_));
 sky130_fd_sc_hd__mux2_1 _07681_ (.A0(\cpuregs[14][3] ),
    .A1(\cpuregs[15][3] ),
    .S(net660),
    .X(_03201_));
 sky130_fd_sc_hd__mux2_1 _07682_ (.A0(\cpuregs[12][3] ),
    .A1(\cpuregs[13][3] ),
    .S(net660),
    .X(_03202_));
 sky130_fd_sc_hd__or2_1 _07683_ (.A(net798),
    .B(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__o211a_1 _07684_ (.A1(net810),
    .A2(_03201_),
    .B1(_03203_),
    .C1(net825),
    .X(_03204_));
 sky130_fd_sc_hd__or2_1 _07685_ (.A(\cpuregs[8][3] ),
    .B(net662),
    .X(_03205_));
 sky130_fd_sc_hd__o211a_1 _07686_ (.A1(\cpuregs[9][3] ),
    .A2(net623),
    .B1(net606),
    .C1(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__or2_1 _07687_ (.A(\cpuregs[10][3] ),
    .B(net661),
    .X(_03207_));
 sky130_fd_sc_hd__o211a_1 _07688_ (.A1(\cpuregs[11][3] ),
    .A2(net623),
    .B1(net592),
    .C1(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__o41a_1 _07689_ (.A1(net788),
    .A2(_03204_),
    .A3(_03206_),
    .A4(_03208_),
    .B1(net776),
    .X(_03209_));
 sky130_fd_sc_hd__mux2_1 _07690_ (.A0(\cpuregs[28][3] ),
    .A1(\cpuregs[29][3] ),
    .S(net677),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _07691_ (.A0(\cpuregs[30][3] ),
    .A1(\cpuregs[31][3] ),
    .S(net677),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _07692_ (.A0(_03210_),
    .A1(_03211_),
    .S(net802),
    .X(_03212_));
 sky130_fd_sc_hd__or2_1 _07693_ (.A(\cpuregs[24][3] ),
    .B(net677),
    .X(_03213_));
 sky130_fd_sc_hd__o211a_1 _07694_ (.A1(\cpuregs[25][3] ),
    .A2(net629),
    .B1(net609),
    .C1(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__or2_1 _07695_ (.A(\cpuregs[26][3] ),
    .B(net677),
    .X(_03215_));
 sky130_fd_sc_hd__o211a_1 _07696_ (.A1(\cpuregs[27][3] ),
    .A2(net629),
    .B1(net595),
    .C1(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__a2111o_1 _07697_ (.A1(net829),
    .A2(_03212_),
    .B1(_03214_),
    .C1(_03216_),
    .D1(net790),
    .X(_03217_));
 sky130_fd_sc_hd__mux2_1 _07698_ (.A0(\cpuregs[20][3] ),
    .A1(\cpuregs[21][3] ),
    .S(net674),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_1 _07699_ (.A0(\cpuregs[22][3] ),
    .A1(\cpuregs[23][3] ),
    .S(net674),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _07700_ (.A0(_03218_),
    .A1(_03219_),
    .S(net801),
    .X(_03220_));
 sky130_fd_sc_hd__or2_1 _07701_ (.A(\cpuregs[16][3] ),
    .B(net676),
    .X(_03221_));
 sky130_fd_sc_hd__o211a_1 _07702_ (.A1(\cpuregs[17][3] ),
    .A2(net630),
    .B1(_03148_),
    .C1(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__o21a_1 _07703_ (.A1(\cpuregs[19][3] ),
    .A2(net630),
    .B1(net595),
    .X(_03223_));
 sky130_fd_sc_hd__o22a_1 _07704_ (.A1(\cpuregs[18][3] ),
    .A2(net552),
    .B1(_03223_),
    .B2(net781),
    .X(_03224_));
 sky130_fd_sc_hd__a211o_1 _07705_ (.A1(net829),
    .A2(_03220_),
    .B1(_03222_),
    .C1(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__and3_1 _07706_ (.A(net772),
    .B(_03217_),
    .C(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__a21oi_4 _07707_ (.A1(_03200_),
    .A2(_03209_),
    .B1(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__nor2_1 _07708_ (.A(net987),
    .B(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_1 _07709_ (.A(\reg_sh[3] ),
    .B(\reg_sh[2] ),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _07710_ (.A(_02473_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__a221o_1 _07711_ (.A1(\decoded_imm_j[3] ),
    .A2(_02701_),
    .B1(_03192_),
    .B2(_03230_),
    .C1(_03228_),
    .X(_06749_));
 sky130_fd_sc_hd__mux2_1 _07712_ (.A0(\cpuregs[6][4] ),
    .A1(\cpuregs[7][4] ),
    .S(net698),
    .X(_03231_));
 sky130_fd_sc_hd__or2_1 _07713_ (.A(\cpuregs[4][4] ),
    .B(net698),
    .X(_03232_));
 sky130_fd_sc_hd__o211a_1 _07714_ (.A1(\cpuregs[5][4] ),
    .A2(net640),
    .B1(net819),
    .C1(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__a211o_1 _07715_ (.A1(net807),
    .A2(_03231_),
    .B1(_03233_),
    .C1(net839),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _07716_ (.A0(\cpuregs[2][4] ),
    .A1(\cpuregs[3][4] ),
    .S(net697),
    .X(_03235_));
 sky130_fd_sc_hd__a221o_1 _07717_ (.A1(\cpuregs[1][4] ),
    .A2(net551),
    .B1(_03235_),
    .B2(net807),
    .C1(net835),
    .X(_03236_));
 sky130_fd_sc_hd__a21o_1 _07718_ (.A1(_03234_),
    .A2(_03236_),
    .B1(net785),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _07719_ (.A0(\cpuregs[14][4] ),
    .A1(\cpuregs[15][4] ),
    .S(net698),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _07720_ (.A0(\cpuregs[12][4] ),
    .A1(\cpuregs[13][4] ),
    .S(net698),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _07721_ (.A0(_03238_),
    .A1(_03239_),
    .S(net819),
    .X(_03240_));
 sky130_fd_sc_hd__or2_1 _07722_ (.A(\cpuregs[8][4] ),
    .B(net697),
    .X(_03241_));
 sky130_fd_sc_hd__o211a_1 _07723_ (.A1(\cpuregs[9][4] ),
    .A2(net640),
    .B1(net614),
    .C1(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__or2_1 _07724_ (.A(\cpuregs[10][4] ),
    .B(net697),
    .X(_03243_));
 sky130_fd_sc_hd__o211a_1 _07725_ (.A1(\cpuregs[11][4] ),
    .A2(net640),
    .B1(net601),
    .C1(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__a211o_1 _07726_ (.A1(net835),
    .A2(_03240_),
    .B1(_03242_),
    .C1(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__o211a_1 _07727_ (.A1(net794),
    .A2(_03245_),
    .B1(_03237_),
    .C1(net778),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _07728_ (.A0(\cpuregs[30][4] ),
    .A1(\cpuregs[31][4] ),
    .S(net678),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _07729_ (.A0(\cpuregs[28][4] ),
    .A1(\cpuregs[29][4] ),
    .S(net701),
    .X(_03248_));
 sky130_fd_sc_hd__mux2_1 _07730_ (.A0(_03247_),
    .A1(_03248_),
    .S(net819),
    .X(_03249_));
 sky130_fd_sc_hd__or2_1 _07731_ (.A(\cpuregs[24][4] ),
    .B(net698),
    .X(_03250_));
 sky130_fd_sc_hd__o211a_1 _07732_ (.A1(\cpuregs[25][4] ),
    .A2(net641),
    .B1(net614),
    .C1(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__or2_1 _07733_ (.A(\cpuregs[26][4] ),
    .B(net698),
    .X(_03252_));
 sky130_fd_sc_hd__o211a_1 _07734_ (.A1(\cpuregs[27][4] ),
    .A2(net631),
    .B1(net595),
    .C1(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__a2111o_1 _07735_ (.A1(net835),
    .A2(_03249_),
    .B1(_03251_),
    .C1(_03253_),
    .D1(net794),
    .X(_03254_));
 sky130_fd_sc_hd__mux2_1 _07736_ (.A0(\cpuregs[20][4] ),
    .A1(\cpuregs[21][4] ),
    .S(net701),
    .X(_03255_));
 sky130_fd_sc_hd__mux2_1 _07737_ (.A0(\cpuregs[22][4] ),
    .A1(\cpuregs[23][4] ),
    .S(net701),
    .X(_03256_));
 sky130_fd_sc_hd__mux2_1 _07738_ (.A0(_03255_),
    .A1(_03256_),
    .S(net807),
    .X(_03257_));
 sky130_fd_sc_hd__or2_1 _07739_ (.A(\cpuregs[16][4] ),
    .B(net698),
    .X(_03258_));
 sky130_fd_sc_hd__o211a_1 _07740_ (.A1(\cpuregs[17][4] ),
    .A2(net641),
    .B1(net614),
    .C1(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__o21a_1 _07741_ (.A1(\cpuregs[19][4] ),
    .A2(net641),
    .B1(net601),
    .X(_03260_));
 sky130_fd_sc_hd__o22a_1 _07742_ (.A1(\cpuregs[18][4] ),
    .A2(net555),
    .B1(_03260_),
    .B2(net785),
    .X(_03261_));
 sky130_fd_sc_hd__a211o_1 _07743_ (.A1(net835),
    .A2(_03257_),
    .B1(_03259_),
    .C1(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__a31oi_4 _07744_ (.A1(net775),
    .A2(_03254_),
    .A3(_03262_),
    .B1(_03246_),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_1 _07745_ (.A(net987),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__a32o_1 _07746_ (.A1(net1066),
    .A2(\reg_sh[4] ),
    .A3(_02473_),
    .B1(_02701_),
    .B2(\decoded_imm_j[4] ),
    .X(_03265_));
 sky130_fd_sc_hd__or3_1 _07747_ (.A(_02478_),
    .B(_03264_),
    .C(_03265_),
    .X(_06750_));
 sky130_fd_sc_hd__nand2_1 _07748_ (.A(net255),
    .B(net996),
    .Y(_03266_));
 sky130_fd_sc_hd__or2_1 _07749_ (.A(net255),
    .B(net996),
    .X(_03267_));
 sky130_fd_sc_hd__nand2_1 _07750_ (.A(_03266_),
    .B(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__or2_1 _07751_ (.A(net252),
    .B(net1002),
    .X(_03269_));
 sky130_fd_sc_hd__nand2_1 _07752_ (.A(net252),
    .B(net1002),
    .Y(_03270_));
 sky130_fd_sc_hd__and2_1 _07753_ (.A(_03269_),
    .B(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__nand2_1 _07754_ (.A(_03269_),
    .B(_03270_),
    .Y(_03272_));
 sky130_fd_sc_hd__and2_1 _07755_ (.A(net1176),
    .B(net1044),
    .X(_03273_));
 sky130_fd_sc_hd__nor2_1 _07756_ (.A(net1176),
    .B(net1044),
    .Y(_03274_));
 sky130_fd_sc_hd__nor2_1 _07757_ (.A(_03273_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__and2_1 _07758_ (.A(net1177),
    .B(net1045),
    .X(_03276_));
 sky130_fd_sc_hd__or2_1 _07759_ (.A(net1177),
    .B(net1045),
    .X(_03277_));
 sky130_fd_sc_hd__nand2b_2 _07760_ (.A_N(_03276_),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__xor2_1 _07761_ (.A(net1181),
    .B(net1053),
    .X(_03279_));
 sky130_fd_sc_hd__nand2_1 _07762_ (.A(net1171),
    .B(net1039),
    .Y(_03280_));
 sky130_fd_sc_hd__inv_2 _07763_ (.A(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__nor2_1 _07764_ (.A(net1171),
    .B(net1039),
    .Y(_03282_));
 sky130_fd_sc_hd__nor2_1 _07765_ (.A(_03281_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__or2_1 _07766_ (.A(net1047),
    .B(net1178),
    .X(_03284_));
 sky130_fd_sc_hd__xor2_2 _07767_ (.A(net1047),
    .B(net1178),
    .X(_03285_));
 sky130_fd_sc_hd__or2_1 _07768_ (.A(net1163),
    .B(net1024),
    .X(_03286_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(net1163),
    .B(net1024),
    .Y(_03287_));
 sky130_fd_sc_hd__and2_2 _07770_ (.A(_03286_),
    .B(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__nand2_1 _07771_ (.A(net254),
    .B(net998),
    .Y(_03289_));
 sky130_fd_sc_hd__or2_1 _07772_ (.A(net254),
    .B(net998),
    .X(_03290_));
 sky130_fd_sc_hd__and2_1 _07773_ (.A(_03289_),
    .B(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__and2_1 _07774_ (.A(net251),
    .B(net1004),
    .X(_03292_));
 sky130_fd_sc_hd__nor2_1 _07775_ (.A(net251),
    .B(net1004),
    .Y(_03293_));
 sky130_fd_sc_hd__nor2_1 _07776_ (.A(_03292_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__nand2_1 _07777_ (.A(net253),
    .B(net1000),
    .Y(_03295_));
 sky130_fd_sc_hd__or2_1 _07778_ (.A(net253),
    .B(net1000),
    .X(_03296_));
 sky130_fd_sc_hd__and2_1 _07779_ (.A(_03295_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__nand2_1 _07780_ (.A(net1164),
    .B(net1026),
    .Y(_03298_));
 sky130_fd_sc_hd__nor2_1 _07781_ (.A(net1164),
    .B(net1026),
    .Y(_03299_));
 sky130_fd_sc_hd__or2_1 _07782_ (.A(net1164),
    .B(net1026),
    .X(_03300_));
 sky130_fd_sc_hd__and2_1 _07783_ (.A(_03298_),
    .B(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__nand2_1 _07784_ (.A(_03298_),
    .B(_03300_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand2_1 _07785_ (.A(net1174),
    .B(net1042),
    .Y(_03303_));
 sky130_fd_sc_hd__nor2_1 _07786_ (.A(net1174),
    .B(net1042),
    .Y(_03304_));
 sky130_fd_sc_hd__or2_1 _07787_ (.A(net1174),
    .B(net1043),
    .X(_03305_));
 sky130_fd_sc_hd__and2_1 _07788_ (.A(_03303_),
    .B(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__nand2_1 _07789_ (.A(_03303_),
    .B(_03305_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand2_1 _07790_ (.A(net1172),
    .B(net1040),
    .Y(_03308_));
 sky130_fd_sc_hd__nor2_1 _07791_ (.A(net1172),
    .B(net1041),
    .Y(_03309_));
 sky130_fd_sc_hd__inv_2 _07792_ (.A(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand2_1 _07793_ (.A(_03308_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand2_1 _07794_ (.A(net256),
    .B(net994),
    .Y(_03312_));
 sky130_fd_sc_hd__or2_1 _07795_ (.A(net256),
    .B(net994),
    .X(_03313_));
 sky130_fd_sc_hd__nand2_1 _07796_ (.A(_03312_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__nand2_1 _07797_ (.A(net1169),
    .B(net1035),
    .Y(_03315_));
 sky130_fd_sc_hd__inv_2 _07798_ (.A(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__nor2_1 _07799_ (.A(net1169),
    .B(net1036),
    .Y(_03317_));
 sky130_fd_sc_hd__nor2_1 _07800_ (.A(_03316_),
    .B(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__and2_1 _07801_ (.A(net1158),
    .B(net1007),
    .X(_03319_));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(net1158),
    .B(net1007),
    .Y(_03320_));
 sky130_fd_sc_hd__nor2_1 _07803_ (.A(net1158),
    .B(net1007),
    .Y(_03321_));
 sky130_fd_sc_hd__or2_1 _07804_ (.A(net1158),
    .B(net1008),
    .X(_03322_));
 sky130_fd_sc_hd__nor2_1 _07805_ (.A(_03319_),
    .B(_03321_),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(_03320_),
    .B(_03322_),
    .Y(_03324_));
 sky130_fd_sc_hd__nand2_1 _07807_ (.A(net250),
    .B(net1006),
    .Y(_03325_));
 sky130_fd_sc_hd__or2_1 _07808_ (.A(net250),
    .B(net1006),
    .X(_03326_));
 sky130_fd_sc_hd__and2_1 _07809_ (.A(_03325_),
    .B(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__and2_1 _07810_ (.A(net247),
    .B(net1010),
    .X(_03328_));
 sky130_fd_sc_hd__nor2_1 _07811_ (.A(net247),
    .B(net1010),
    .Y(_03329_));
 sky130_fd_sc_hd__nor2_1 _07812_ (.A(_03328_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__or2_1 _07813_ (.A(net248),
    .B(net1009),
    .X(_03331_));
 sky130_fd_sc_hd__nand2_1 _07814_ (.A(net248),
    .B(net1009),
    .Y(_03332_));
 sky130_fd_sc_hd__and2_1 _07815_ (.A(_03331_),
    .B(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__inv_2 _07816_ (.A(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__or4_1 _07817_ (.A(_03323_),
    .B(_03327_),
    .C(_03330_),
    .D(_03333_),
    .X(_03335_));
 sky130_fd_sc_hd__xor2_2 _07818_ (.A(net1159),
    .B(net1012),
    .X(_03336_));
 sky130_fd_sc_hd__and2_1 _07819_ (.A(net244),
    .B(net1014),
    .X(_03337_));
 sky130_fd_sc_hd__nor2_1 _07820_ (.A(net244),
    .B(net1014),
    .Y(_03338_));
 sky130_fd_sc_hd__nor2_1 _07821_ (.A(_03337_),
    .B(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__or2_1 _07822_ (.A(_03336_),
    .B(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__nor2_1 _07823_ (.A(_02395_),
    .B(_02407_),
    .Y(_03341_));
 sky130_fd_sc_hd__nor2_1 _07824_ (.A(net1161),
    .B(net1018),
    .Y(_03342_));
 sky130_fd_sc_hd__nor2_1 _07825_ (.A(_03341_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__or2_1 _07826_ (.A(net1160),
    .B(net1016),
    .X(_03344_));
 sky130_fd_sc_hd__and2_1 _07827_ (.A(net1160),
    .B(net1016),
    .X(_03345_));
 sky130_fd_sc_hd__nand2_1 _07828_ (.A(net1160),
    .B(net1016),
    .Y(_03346_));
 sky130_fd_sc_hd__and2_1 _07829_ (.A(_03344_),
    .B(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__or3_1 _07830_ (.A(_03340_),
    .B(_03343_),
    .C(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__or2_1 _07831_ (.A(net1167),
    .B(net1031),
    .X(_03349_));
 sky130_fd_sc_hd__nand2_1 _07832_ (.A(net1167),
    .B(net1031),
    .Y(_03350_));
 sky130_fd_sc_hd__and2_1 _07833_ (.A(_03349_),
    .B(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__nand2_1 _07834_ (.A(net1168),
    .B(net1033),
    .Y(_03352_));
 sky130_fd_sc_hd__or2_1 _07835_ (.A(net1168),
    .B(net1033),
    .X(_03353_));
 sky130_fd_sc_hd__and2_1 _07836_ (.A(_03352_),
    .B(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__inv_2 _07837_ (.A(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__or2_1 _07838_ (.A(_03351_),
    .B(_03354_),
    .X(_03356_));
 sky130_fd_sc_hd__nand2_1 _07839_ (.A(net1166),
    .B(net1029),
    .Y(_03357_));
 sky130_fd_sc_hd__nor2_1 _07840_ (.A(net1166),
    .B(net1029),
    .Y(_03358_));
 sky130_fd_sc_hd__or2_1 _07841_ (.A(net1166),
    .B(net1029),
    .X(_03359_));
 sky130_fd_sc_hd__nand2_2 _07842_ (.A(_03357_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(net1165),
    .B(net1028),
    .Y(_03361_));
 sky130_fd_sc_hd__nor2_1 _07844_ (.A(net1165),
    .B(net1028),
    .Y(_03362_));
 sky130_fd_sc_hd__or2_1 _07845_ (.A(net1165),
    .B(net1028),
    .X(_03363_));
 sky130_fd_sc_hd__nand2_2 _07846_ (.A(_03361_),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand2_1 _07847_ (.A(_03360_),
    .B(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__nand2_1 _07848_ (.A(net1188),
    .B(net1157),
    .Y(_03366_));
 sky130_fd_sc_hd__or2_1 _07849_ (.A(net1188),
    .B(net1157),
    .X(_03367_));
 sky130_fd_sc_hd__and2_2 _07850_ (.A(_03366_),
    .B(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__inv_2 _07851_ (.A(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__and2_1 _07852_ (.A(net258),
    .B(net992),
    .X(_03370_));
 sky130_fd_sc_hd__nor2_1 _07853_ (.A(net258),
    .B(net992),
    .Y(_03371_));
 sky130_fd_sc_hd__or2_1 _07854_ (.A(_03370_),
    .B(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__and2_1 _07855_ (.A(_03369_),
    .B(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__and2_1 _07856_ (.A(net1162),
    .B(net1020),
    .X(_03374_));
 sky130_fd_sc_hd__or2_1 _07857_ (.A(net1162),
    .B(net1020),
    .X(_03375_));
 sky130_fd_sc_hd__nand2b_2 _07858_ (.A_N(_03374_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__and2_1 _07859_ (.A(net240),
    .B(net1022),
    .X(_03377_));
 sky130_fd_sc_hd__nor2_1 _07860_ (.A(net240),
    .B(net1022),
    .Y(_03378_));
 sky130_fd_sc_hd__or2_2 _07861_ (.A(_03377_),
    .B(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(_03291_),
    .B(_03297_),
    .Y(_03380_));
 sky130_fd_sc_hd__and3_1 _07863_ (.A(_03268_),
    .B(_03314_),
    .C(_03373_),
    .X(_03381_));
 sky130_fd_sc_hd__or4bb_1 _07864_ (.A(_03271_),
    .B(_03294_),
    .C_N(_03380_),
    .D_N(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__nand2_1 _07865_ (.A(_03278_),
    .B(_03311_),
    .Y(_03383_));
 sky130_fd_sc_hd__or2_1 _07866_ (.A(_03283_),
    .B(_03318_),
    .X(_03384_));
 sky130_fd_sc_hd__or3_1 _07867_ (.A(_03275_),
    .B(_03279_),
    .C(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__or4_1 _07868_ (.A(_03285_),
    .B(_03306_),
    .C(_03383_),
    .D(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__or4bb_1 _07869_ (.A(_03288_),
    .B(_03301_),
    .C_N(_03376_),
    .D_N(_03379_),
    .X(_03387_));
 sky130_fd_sc_hd__or4_1 _07870_ (.A(_03335_),
    .B(_03348_),
    .C(_03356_),
    .D(_03365_),
    .X(_03388_));
 sky130_fd_sc_hd__or4_2 _07871_ (.A(_03382_),
    .B(_03386_),
    .C(_03387_),
    .D(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__nor2_1 _07872_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .Y(_03390_));
 sky130_fd_sc_hd__and4_1 _07873_ (.A(_02365_),
    .B(_02366_),
    .C(_02413_),
    .D(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__and2_1 _07874_ (.A(_03389_),
    .B(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__and2b_1 _07875_ (.A_N(net1157),
    .B(net1188),
    .X(_03393_));
 sky130_fd_sc_hd__nand2b_1 _07876_ (.A_N(net258),
    .B(net992),
    .Y(_03394_));
 sky130_fd_sc_hd__nor2_1 _07877_ (.A(_03368_),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__and2b_1 _07878_ (.A_N(net253),
    .B(net1001),
    .X(_03396_));
 sky130_fd_sc_hd__or2_1 _07879_ (.A(net1160),
    .B(_02408_),
    .X(_03397_));
 sky130_fd_sc_hd__o31a_1 _07880_ (.A1(net1161),
    .A2(_02407_),
    .A3(_03347_),
    .B1(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__or2_1 _07881_ (.A(net1159),
    .B(_02409_),
    .X(_03399_));
 sky130_fd_sc_hd__nand2b_1 _07882_ (.A_N(net244),
    .B(net1015),
    .Y(_03400_));
 sky130_fd_sc_hd__o221a_1 _07883_ (.A1(_03340_),
    .A2(_03398_),
    .B1(_03400_),
    .B2(_03336_),
    .C1(_03399_),
    .X(_03401_));
 sky130_fd_sc_hd__and2b_1 _07884_ (.A_N(net247),
    .B(net1010),
    .X(_03402_));
 sky130_fd_sc_hd__nand2_1 _07885_ (.A(_03334_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__o21ai_1 _07886_ (.A1(net248),
    .A2(_02410_),
    .B1(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__and2b_1 _07887_ (.A_N(net1158),
    .B(net1008),
    .X(_03405_));
 sky130_fd_sc_hd__a21oi_1 _07888_ (.A1(_03324_),
    .A2(_03404_),
    .B1(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__or2_1 _07889_ (.A(_03327_),
    .B(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__o221a_1 _07890_ (.A1(net250),
    .A2(_02411_),
    .B1(_03335_),
    .B2(_03401_),
    .C1(_03407_),
    .X(_03408_));
 sky130_fd_sc_hd__and2b_1 _07891_ (.A_N(net1162),
    .B(net1020),
    .X(_03409_));
 sky130_fd_sc_hd__a31o_1 _07892_ (.A1(_02394_),
    .A2(net1022),
    .A3(_03376_),
    .B1(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__and2b_1 _07893_ (.A_N(net1166),
    .B(net1030),
    .X(_03411_));
 sky130_fd_sc_hd__or2_1 _07894_ (.A(net1167),
    .B(_02403_),
    .X(_03412_));
 sky130_fd_sc_hd__nand2b_1 _07895_ (.A_N(net1168),
    .B(net1033),
    .Y(_03413_));
 sky130_fd_sc_hd__o21ai_1 _07896_ (.A1(_03351_),
    .A2(_03413_),
    .B1(_03412_),
    .Y(_03414_));
 sky130_fd_sc_hd__a21o_1 _07897_ (.A1(_03360_),
    .A2(_03414_),
    .B1(_03411_),
    .X(_03415_));
 sky130_fd_sc_hd__nand2_1 _07898_ (.A(_03364_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__o21a_1 _07899_ (.A1(net1165),
    .A2(_02404_),
    .B1(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__and2b_1 _07900_ (.A_N(net1172),
    .B(net1041),
    .X(_03418_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(net1176),
    .B(_02402_),
    .Y(_03419_));
 sky130_fd_sc_hd__and2b_1 _07902_ (.A_N(net1177),
    .B(net1046),
    .X(_03420_));
 sky130_fd_sc_hd__nand2b_1 _07903_ (.A_N(net1178),
    .B(net1049),
    .Y(_03421_));
 sky130_fd_sc_hd__and2b_1 _07904_ (.A_N(net1051),
    .B(net1180),
    .X(_03422_));
 sky130_fd_sc_hd__o21ai_1 _07905_ (.A1(_03285_),
    .A2(_03422_),
    .B1(_03421_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21oi_1 _07906_ (.A1(_03278_),
    .A2(_03423_),
    .B1(_03420_),
    .Y(_03424_));
 sky130_fd_sc_hd__a221o_1 _07907_ (.A1(_02392_),
    .A2(net228),
    .B1(_03278_),
    .B2(_03423_),
    .C1(_03420_),
    .X(_03425_));
 sky130_fd_sc_hd__a32o_1 _07908_ (.A1(_03307_),
    .A2(_03419_),
    .A3(_03425_),
    .B1(net1043),
    .B2(_02393_),
    .X(_03426_));
 sky130_fd_sc_hd__a21oi_1 _07909_ (.A1(_03311_),
    .A2(_03426_),
    .B1(_03418_),
    .Y(_03427_));
 sky130_fd_sc_hd__or2_1 _07910_ (.A(_03283_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__nand2b_1 _07911_ (.A_N(net1171),
    .B(net1039),
    .Y(_03429_));
 sky130_fd_sc_hd__nand2b_1 _07912_ (.A_N(net1169),
    .B(net1036),
    .Y(_03430_));
 sky130_fd_sc_hd__o221a_1 _07913_ (.A1(_03384_),
    .A2(_03427_),
    .B1(_03429_),
    .B2(_03318_),
    .C1(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__o31ai_1 _07914_ (.A1(_03356_),
    .A2(_03365_),
    .A3(_03431_),
    .B1(_03417_),
    .Y(_03432_));
 sky130_fd_sc_hd__nand2_1 _07915_ (.A(_03302_),
    .B(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__o21a_1 _07916_ (.A1(net1164),
    .A2(_02405_),
    .B1(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__or3_1 _07917_ (.A(net1164),
    .B(_02405_),
    .C(_03288_),
    .X(_03435_));
 sky130_fd_sc_hd__o221ai_4 _07918_ (.A1(net1163),
    .A2(_02406_),
    .B1(_03288_),
    .B2(_03433_),
    .C1(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__a31oi_4 _07919_ (.A1(_03376_),
    .A2(_03379_),
    .A3(_03436_),
    .B1(_03410_),
    .Y(_03437_));
 sky130_fd_sc_hd__o31a_1 _07920_ (.A1(_03335_),
    .A2(_03348_),
    .A3(_03437_),
    .B1(_03408_),
    .X(_03438_));
 sky130_fd_sc_hd__nor2_1 _07921_ (.A(_03294_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__and2b_1 _07922_ (.A_N(net252),
    .B(net1002),
    .X(_03440_));
 sky130_fd_sc_hd__a31o_1 _07923_ (.A1(_02396_),
    .A2(net1004),
    .A3(_03272_),
    .B1(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__a21oi_1 _07924_ (.A1(_03272_),
    .A2(_03439_),
    .B1(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__o21ba_1 _07925_ (.A1(_03297_),
    .A2(_03442_),
    .B1_N(_03396_),
    .X(_03443_));
 sky130_fd_sc_hd__and3_1 _07926_ (.A(_03272_),
    .B(_03380_),
    .C(_03439_),
    .X(_03444_));
 sky130_fd_sc_hd__and2b_1 _07927_ (.A_N(_03291_),
    .B(_03396_),
    .X(_03445_));
 sky130_fd_sc_hd__a221o_1 _07928_ (.A1(_02397_),
    .A2(net998),
    .B1(_03380_),
    .B2(_03441_),
    .C1(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__o21a_1 _07929_ (.A1(_03444_),
    .A2(_03446_),
    .B1(_03268_),
    .X(_03447_));
 sky130_fd_sc_hd__a22o_1 _07930_ (.A1(_02399_),
    .A2(net996),
    .B1(net994),
    .B2(_02398_),
    .X(_03448_));
 sky130_fd_sc_hd__o22a_1 _07931_ (.A1(_02398_),
    .A2(net995),
    .B1(_03447_),
    .B2(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__nand2_1 _07932_ (.A(_03373_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__or3b_1 _07933_ (.A(_03393_),
    .B(_03395_),
    .C_N(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__a31o_1 _07934_ (.A1(_03369_),
    .A2(_03394_),
    .A3(_03450_),
    .B1(_03393_),
    .X(_03452_));
 sky130_fd_sc_hd__or2_1 _07935_ (.A(_02366_),
    .B(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__mux2_1 _07936_ (.A0(_02413_),
    .A1(_02365_),
    .S(_03451_),
    .X(_03454_));
 sky130_fd_sc_hd__a221oi_1 _07937_ (.A1(instr_bne),
    .A2(_03389_),
    .B1(_03452_),
    .B2(is_slti_blt_slt),
    .C1(_03391_),
    .Y(_03455_));
 sky130_fd_sc_hd__a31o_1 _07938_ (.A1(_03453_),
    .A2(_03454_),
    .A3(_03455_),
    .B1(_03392_),
    .X(_03456_));
 sky130_fd_sc_hd__inv_2 _07939_ (.A(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__a21oi_1 _07940_ (.A1(_02377_),
    .A2(_02384_),
    .B1(net969),
    .Y(_03458_));
 sky130_fd_sc_hd__nor2_2 _07941_ (.A(instr_and),
    .B(instr_andi),
    .Y(_03459_));
 sky130_fd_sc_hd__or2_1 _07942_ (.A(instr_and),
    .B(instr_andi),
    .X(_03460_));
 sky130_fd_sc_hd__a31o_1 _07943_ (.A1(net1181),
    .A2(net1053),
    .A3(net933),
    .B1(_03458_),
    .X(_03461_));
 sky130_fd_sc_hd__nor2_2 _07944_ (.A(instr_xor),
    .B(instr_xori),
    .Y(_03462_));
 sky130_fd_sc_hd__or2_1 _07945_ (.A(instr_xor),
    .B(instr_xori),
    .X(_03463_));
 sky130_fd_sc_hd__and4b_2 _07946_ (.A_N(is_compare),
    .B(net969),
    .C(net935),
    .D(net931),
    .X(_03464_));
 sky130_fd_sc_hd__or4_4 _07947_ (.A(is_compare),
    .B(_02433_),
    .C(net933),
    .D(net928),
    .X(_03465_));
 sky130_fd_sc_hd__o21a_1 _07948_ (.A1(net929),
    .A2(net771),
    .B1(_03279_),
    .X(_03466_));
 sky130_fd_sc_hd__a211o_1 _07949_ (.A1(net3052),
    .A2(_03457_),
    .B1(_03461_),
    .C1(_03466_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__and3_1 _07950_ (.A(net1047),
    .B(net1178),
    .C(net932),
    .X(_03467_));
 sky130_fd_sc_hd__a221o_1 _07951_ (.A1(net967),
    .A2(_03284_),
    .B1(_03285_),
    .B2(net928),
    .C1(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__xnor2_1 _07952_ (.A(_03285_),
    .B(_03422_),
    .Y(_03469_));
 sky130_fd_sc_hd__o21ai_1 _07953_ (.A1(net1143),
    .A2(_02377_),
    .B1(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__or3_1 _07954_ (.A(net1144),
    .B(_02377_),
    .C(_03469_),
    .X(_03471_));
 sky130_fd_sc_hd__a31o_1 _07955_ (.A1(net771),
    .A2(_03470_),
    .A3(_03471_),
    .B1(_03468_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__nor2_1 _07956_ (.A(_03278_),
    .B(net930),
    .Y(_03472_));
 sky130_fd_sc_hd__a221o_1 _07957_ (.A1(net967),
    .A2(_03277_),
    .B1(net932),
    .B2(_03276_),
    .C1(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__a22o_1 _07958_ (.A1(net1180),
    .A2(net1051),
    .B1(net1178),
    .B2(net1049),
    .X(_03474_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(_03284_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__mux2_1 _07960_ (.A0(_03423_),
    .A1(_03475_),
    .S(net989),
    .X(_03476_));
 sky130_fd_sc_hd__or2_1 _07961_ (.A(_03278_),
    .B(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__nand2_1 _07962_ (.A(_03278_),
    .B(_03476_),
    .Y(_03478_));
 sky130_fd_sc_hd__a31o_1 _07963_ (.A1(net771),
    .A2(_03477_),
    .A3(_03478_),
    .B1(_03473_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__o21a_1 _07964_ (.A1(_03273_),
    .A2(net930),
    .B1(net968),
    .X(_03479_));
 sky130_fd_sc_hd__nor2_1 _07965_ (.A(_03274_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__a31o_1 _07966_ (.A1(_03277_),
    .A2(_03284_),
    .A3(_03474_),
    .B1(_03276_),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _07967_ (.A0(_03424_),
    .A1(_03481_),
    .S(net989),
    .X(_03482_));
 sky130_fd_sc_hd__a21oi_1 _07968_ (.A1(_03275_),
    .A2(_03482_),
    .B1(_03465_),
    .Y(_03483_));
 sky130_fd_sc_hd__o21a_1 _07969_ (.A1(_03275_),
    .A2(_03482_),
    .B1(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__a211o_1 _07970_ (.A1(_03273_),
    .A2(net932),
    .B1(_03480_),
    .C1(_03484_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__o22a_1 _07971_ (.A1(net968),
    .A2(_03304_),
    .B1(net934),
    .B2(_03303_),
    .X(_03485_));
 sky130_fd_sc_hd__o21ai_1 _07972_ (.A1(_03307_),
    .A2(net930),
    .B1(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__a311oi_2 _07973_ (.A1(_03277_),
    .A2(_03284_),
    .A3(_03474_),
    .B1(_03276_),
    .C1(_03273_),
    .Y(_03487_));
 sky130_fd_sc_hd__a21o_1 _07974_ (.A1(_03419_),
    .A2(_03425_),
    .B1(net989),
    .X(_03488_));
 sky130_fd_sc_hd__o31ai_1 _07975_ (.A1(net1144),
    .A2(_03274_),
    .A3(_03487_),
    .B1(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(_03306_),
    .B(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__o21a_1 _07977_ (.A1(_03306_),
    .A2(_03489_),
    .B1(net770),
    .X(_03491_));
 sky130_fd_sc_hd__a21o_1 _07978_ (.A1(_03490_),
    .A2(_03491_),
    .B1(_03486_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__or2_1 _07979_ (.A(_03308_),
    .B(net934),
    .X(_03492_));
 sky130_fd_sc_hd__o221a_1 _07980_ (.A1(net968),
    .A2(_03309_),
    .B1(_03311_),
    .B2(net930),
    .C1(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__or3_1 _07981_ (.A(_03274_),
    .B(_03304_),
    .C(_03487_),
    .X(_03494_));
 sky130_fd_sc_hd__and3_1 _07982_ (.A(net988),
    .B(_03303_),
    .C(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__a21o_1 _07983_ (.A1(net1143),
    .A2(_03426_),
    .B1(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__o21ai_1 _07984_ (.A1(_03311_),
    .A2(_03496_),
    .B1(net771),
    .Y(_03497_));
 sky130_fd_sc_hd__a21o_1 _07985_ (.A1(_03311_),
    .A2(_03496_),
    .B1(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__nand2_1 _07986_ (.A(_03493_),
    .B(_03498_),
    .Y(\alu_out[5] ));
 sky130_fd_sc_hd__nand2_1 _07987_ (.A(_03283_),
    .B(net928),
    .Y(_03499_));
 sky130_fd_sc_hd__o221a_1 _07988_ (.A1(net968),
    .A2(_03282_),
    .B1(net934),
    .B2(_03280_),
    .C1(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__a31o_1 _07989_ (.A1(_03303_),
    .A2(_03308_),
    .A3(_03494_),
    .B1(_03309_),
    .X(_03501_));
 sky130_fd_sc_hd__nand2_1 _07990_ (.A(net988),
    .B(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__o21a_1 _07991_ (.A1(net988),
    .A2(_03427_),
    .B1(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__o21ai_1 _07992_ (.A1(_03283_),
    .A2(_03503_),
    .B1(net770),
    .Y(_03504_));
 sky130_fd_sc_hd__a21o_1 _07993_ (.A1(_03283_),
    .A2(_03503_),
    .B1(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__nand2_1 _07994_ (.A(_03500_),
    .B(_03505_),
    .Y(\alu_out[6] ));
 sky130_fd_sc_hd__nand2_1 _07995_ (.A(_03318_),
    .B(net928),
    .Y(_03506_));
 sky130_fd_sc_hd__o221a_1 _07996_ (.A1(net968),
    .A2(_03317_),
    .B1(net934),
    .B2(_03315_),
    .C1(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__a21o_1 _07997_ (.A1(_03280_),
    .A2(_03501_),
    .B1(_03282_),
    .X(_03508_));
 sky130_fd_sc_hd__nor2_1 _07998_ (.A(net1143),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__a31o_1 _07999_ (.A1(net1143),
    .A2(_03428_),
    .A3(_03429_),
    .B1(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__nor2_1 _08000_ (.A(_03318_),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__a21o_1 _08001_ (.A1(_03318_),
    .A2(_03510_),
    .B1(_03465_),
    .X(_03512_));
 sky130_fd_sc_hd__o21ai_1 _08002_ (.A1(_03511_),
    .A2(_03512_),
    .B1(_03507_),
    .Y(\alu_out[7] ));
 sky130_fd_sc_hd__nor2_1 _08003_ (.A(_03352_),
    .B(net934),
    .Y(_03513_));
 sky130_fd_sc_hd__a221o_1 _08004_ (.A1(net967),
    .A2(_03353_),
    .B1(_03354_),
    .B2(net928),
    .C1(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__a21oi_1 _08005_ (.A1(_03315_),
    .A2(_03508_),
    .B1(_03317_),
    .Y(_03515_));
 sky130_fd_sc_hd__mux2_1 _08006_ (.A0(_03431_),
    .A1(_03515_),
    .S(net988),
    .X(_03516_));
 sky130_fd_sc_hd__nand2_1 _08007_ (.A(_03354_),
    .B(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__or2_1 _08008_ (.A(_03354_),
    .B(_03516_),
    .X(_03518_));
 sky130_fd_sc_hd__a31o_1 _08009_ (.A1(net770),
    .A2(_03517_),
    .A3(_03518_),
    .B1(_03514_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__nor2_1 _08010_ (.A(_03350_),
    .B(net934),
    .Y(_03519_));
 sky130_fd_sc_hd__a221o_1 _08011_ (.A1(net967),
    .A2(_03349_),
    .B1(_03351_),
    .B2(net928),
    .C1(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__o21a_1 _08012_ (.A1(_03354_),
    .A2(_03431_),
    .B1(_03413_),
    .X(_03521_));
 sky130_fd_sc_hd__a211oi_2 _08013_ (.A1(_03315_),
    .A2(_03508_),
    .B1(_03355_),
    .C1(_03317_),
    .Y(_03522_));
 sky130_fd_sc_hd__a211o_1 _08014_ (.A1(net1168),
    .A2(net1033),
    .B1(_03522_),
    .C1(net1143),
    .X(_03523_));
 sky130_fd_sc_hd__o21ai_1 _08015_ (.A1(net988),
    .A2(_03521_),
    .B1(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__xnor2_1 _08016_ (.A(_03351_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__a21o_1 _08017_ (.A1(net770),
    .A2(_03525_),
    .B1(_03520_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__or2_1 _08018_ (.A(_03357_),
    .B(net934),
    .X(_03526_));
 sky130_fd_sc_hd__o221a_1 _08019_ (.A1(net968),
    .A2(_03358_),
    .B1(_03360_),
    .B2(net930),
    .C1(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__nand2_1 _08020_ (.A(_03350_),
    .B(_03352_),
    .Y(_03528_));
 sky130_fd_sc_hd__o21ai_1 _08021_ (.A1(_03522_),
    .A2(_03528_),
    .B1(_03349_),
    .Y(_03529_));
 sky130_fd_sc_hd__o21bai_1 _08022_ (.A1(_03356_),
    .A2(_03431_),
    .B1_N(_03414_),
    .Y(_03530_));
 sky130_fd_sc_hd__mux2_1 _08023_ (.A0(_03529_),
    .A1(_03530_),
    .S(net1143),
    .X(_03531_));
 sky130_fd_sc_hd__nor2_1 _08024_ (.A(_03360_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__a21o_1 _08025_ (.A1(_03360_),
    .A2(_03531_),
    .B1(_03465_),
    .X(_03533_));
 sky130_fd_sc_hd__o21ai_1 _08026_ (.A1(_03532_),
    .A2(_03533_),
    .B1(_03527_),
    .Y(\alu_out[10] ));
 sky130_fd_sc_hd__or2_1 _08027_ (.A(_03364_),
    .B(net930),
    .X(_03534_));
 sky130_fd_sc_hd__o221a_1 _08028_ (.A1(net968),
    .A2(_03362_),
    .B1(net934),
    .B2(_03361_),
    .C1(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__a21o_1 _08029_ (.A1(_03360_),
    .A2(_03530_),
    .B1(_03411_),
    .X(_03536_));
 sky130_fd_sc_hd__o211a_1 _08030_ (.A1(_03358_),
    .A2(_03529_),
    .B1(net988),
    .C1(_03357_),
    .X(_03537_));
 sky130_fd_sc_hd__a21o_1 _08031_ (.A1(net1143),
    .A2(_03536_),
    .B1(_03537_),
    .X(_03538_));
 sky130_fd_sc_hd__o21ai_1 _08032_ (.A1(_03364_),
    .A2(_03538_),
    .B1(net770),
    .Y(_03539_));
 sky130_fd_sc_hd__a21o_1 _08033_ (.A1(_03364_),
    .A2(_03538_),
    .B1(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__nand2_1 _08034_ (.A(_03535_),
    .B(_03540_),
    .Y(\alu_out[11] ));
 sky130_fd_sc_hd__o22a_1 _08035_ (.A1(net968),
    .A2(_03299_),
    .B1(net934),
    .B2(_03298_),
    .X(_03541_));
 sky130_fd_sc_hd__o21ai_1 _08036_ (.A1(_03302_),
    .A2(net930),
    .B1(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand2_1 _08037_ (.A(_03351_),
    .B(_03522_),
    .Y(_03543_));
 sky130_fd_sc_hd__or4bb_1 _08038_ (.A(_03360_),
    .B(_03364_),
    .C_N(_03528_),
    .D_N(_03349_),
    .X(_03544_));
 sky130_fd_sc_hd__o211a_1 _08039_ (.A1(_03357_),
    .A2(_03362_),
    .B1(_03544_),
    .C1(_03361_),
    .X(_03545_));
 sky130_fd_sc_hd__o31a_1 _08040_ (.A1(_03360_),
    .A2(_03364_),
    .A3(_03543_),
    .B1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_1 _08041_ (.A0(_03432_),
    .A1(_03546_),
    .S(net988),
    .X(_03547_));
 sky130_fd_sc_hd__nand2_1 _08042_ (.A(_03302_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__or2_1 _08043_ (.A(_03302_),
    .B(_03547_),
    .X(_03549_));
 sky130_fd_sc_hd__a31o_1 _08044_ (.A1(net770),
    .A2(_03548_),
    .A3(_03549_),
    .B1(_03542_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__nor2_1 _08045_ (.A(_03287_),
    .B(net934),
    .Y(_03550_));
 sky130_fd_sc_hd__a221o_1 _08046_ (.A1(net967),
    .A2(_03286_),
    .B1(_03288_),
    .B2(net928),
    .C1(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__o21ai_1 _08047_ (.A1(_03299_),
    .A2(_03546_),
    .B1(_03298_),
    .Y(_03552_));
 sky130_fd_sc_hd__mux2_1 _08048_ (.A0(_03434_),
    .A1(_03552_),
    .S(net988),
    .X(_03553_));
 sky130_fd_sc_hd__or2_1 _08049_ (.A(_03288_),
    .B(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_03288_),
    .B(_03553_),
    .Y(_03555_));
 sky130_fd_sc_hd__a31o_1 _08051_ (.A1(net770),
    .A2(_03554_),
    .A3(_03555_),
    .B1(_03551_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__o2bb2a_1 _08052_ (.A1_N(_03377_),
    .A2_N(net932),
    .B1(_03378_),
    .B2(net968),
    .X(_03556_));
 sky130_fd_sc_hd__o21ai_1 _08053_ (.A1(_03379_),
    .A2(net930),
    .B1(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__nand2_1 _08054_ (.A(_03288_),
    .B(_03301_),
    .Y(_03558_));
 sky130_fd_sc_hd__nand2_1 _08055_ (.A(_03287_),
    .B(_03298_),
    .Y(_03559_));
 sky130_fd_sc_hd__o2bb2a_1 _08056_ (.A1_N(_03286_),
    .A2_N(_03559_),
    .B1(_03558_),
    .B2(_03546_),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_1 _08057_ (.A0(_03436_),
    .A1(_03560_),
    .S(net988),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_1 _08058_ (.A(_03379_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__or2_1 _08059_ (.A(_03379_),
    .B(_03561_),
    .X(_03563_));
 sky130_fd_sc_hd__a31o_1 _08060_ (.A1(net770),
    .A2(_03562_),
    .A3(_03563_),
    .B1(_03557_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__nor2_1 _08061_ (.A(_03376_),
    .B(net930),
    .Y(_03564_));
 sky130_fd_sc_hd__a221o_1 _08062_ (.A1(net967),
    .A2(_03375_),
    .B1(net932),
    .B2(_03374_),
    .C1(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__and2_1 _08063_ (.A(_03379_),
    .B(_03436_),
    .X(_03566_));
 sky130_fd_sc_hd__a21o_1 _08064_ (.A1(_02394_),
    .A2(net1023),
    .B1(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__o21ba_1 _08065_ (.A1(_03378_),
    .A2(_03560_),
    .B1_N(_03377_),
    .X(_03568_));
 sky130_fd_sc_hd__mux2_1 _08066_ (.A0(_03567_),
    .A1(_03568_),
    .S(net988),
    .X(_03569_));
 sky130_fd_sc_hd__or2_1 _08067_ (.A(_03376_),
    .B(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__nand2_1 _08068_ (.A(_03376_),
    .B(_03569_),
    .Y(_03571_));
 sky130_fd_sc_hd__a31o_1 _08069_ (.A1(net770),
    .A2(_03570_),
    .A3(_03571_),
    .B1(_03565_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__nor2_1 _08070_ (.A(net968),
    .B(_03342_),
    .Y(_03572_));
 sky130_fd_sc_hd__a221o_1 _08071_ (.A1(_03341_),
    .A2(net932),
    .B1(net928),
    .B2(_03343_),
    .C1(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__nor3_1 _08072_ (.A(_03379_),
    .B(_03546_),
    .C(_03558_),
    .Y(_03574_));
 sky130_fd_sc_hd__and3b_1 _08073_ (.A_N(_03379_),
    .B(_03559_),
    .C(_03286_),
    .X(_03575_));
 sky130_fd_sc_hd__o41a_1 _08074_ (.A1(_03374_),
    .A2(_03377_),
    .A3(_03574_),
    .A4(_03575_),
    .B1(_03375_),
    .X(_03576_));
 sky130_fd_sc_hd__mux2_1 _08075_ (.A0(_03437_),
    .A1(_03576_),
    .S(net989),
    .X(_03577_));
 sky130_fd_sc_hd__or2_1 _08076_ (.A(_03343_),
    .B(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nand2_1 _08077_ (.A(_03343_),
    .B(_03577_),
    .Y(_03579_));
 sky130_fd_sc_hd__a31o_1 _08078_ (.A1(net771),
    .A2(_03578_),
    .A3(_03579_),
    .B1(_03573_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__a21o_1 _08079_ (.A1(_03346_),
    .A2(net928),
    .B1(net967),
    .X(_03580_));
 sky130_fd_sc_hd__nor2_1 _08080_ (.A(_03341_),
    .B(_03576_),
    .Y(_03581_));
 sky130_fd_sc_hd__or2_1 _08081_ (.A(_03343_),
    .B(_03437_),
    .X(_03582_));
 sky130_fd_sc_hd__o211ai_1 _08082_ (.A1(net1161),
    .A2(_02407_),
    .B1(_03582_),
    .C1(net1143),
    .Y(_03583_));
 sky130_fd_sc_hd__o31a_1 _08083_ (.A1(net1143),
    .A2(_03342_),
    .A3(_03581_),
    .B1(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__xnor2_1 _08084_ (.A(_03347_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__a22o_1 _08085_ (.A1(_03345_),
    .A2(net932),
    .B1(net770),
    .B2(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__a21o_1 _08086_ (.A1(_03344_),
    .A2(_03580_),
    .B1(_03586_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__nor2_1 _08087_ (.A(_03337_),
    .B(net930),
    .Y(_03587_));
 sky130_fd_sc_hd__o21ba_1 _08088_ (.A1(net967),
    .A2(_03587_),
    .B1_N(_03338_),
    .X(_03588_));
 sky130_fd_sc_hd__o21a_1 _08089_ (.A1(_03347_),
    .A2(_03582_),
    .B1(_03398_),
    .X(_03589_));
 sky130_fd_sc_hd__and3_1 _08090_ (.A(_03343_),
    .B(_03347_),
    .C(_03576_),
    .X(_03590_));
 sky130_fd_sc_hd__a31o_1 _08091_ (.A1(net1161),
    .A2(net1018),
    .A3(_03344_),
    .B1(_03345_),
    .X(_03591_));
 sky130_fd_sc_hd__inv_2 _08092_ (.A(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__nor2_1 _08093_ (.A(_03590_),
    .B(_03591_),
    .Y(_03593_));
 sky130_fd_sc_hd__inv_2 _08094_ (.A(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__mux2_1 _08095_ (.A0(_03589_),
    .A1(_03594_),
    .S(net989),
    .X(_03595_));
 sky130_fd_sc_hd__a21oi_1 _08096_ (.A1(_03339_),
    .A2(_03595_),
    .B1(_03465_),
    .Y(_03596_));
 sky130_fd_sc_hd__o21a_1 _08097_ (.A1(_03339_),
    .A2(_03595_),
    .B1(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__a211o_1 _08098_ (.A1(_03337_),
    .A2(net932),
    .B1(_03588_),
    .C1(_03597_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__o21a_1 _08099_ (.A1(net1159),
    .A2(net1012),
    .B1(net967),
    .X(_03598_));
 sky130_fd_sc_hd__a31o_1 _08100_ (.A1(net1159),
    .A2(net1013),
    .A3(net932),
    .B1(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__o21ai_1 _08101_ (.A1(_03339_),
    .A2(_03589_),
    .B1(_03400_),
    .Y(_03600_));
 sky130_fd_sc_hd__or2_1 _08102_ (.A(_03338_),
    .B(_03593_),
    .X(_03601_));
 sky130_fd_sc_hd__nor2_1 _08103_ (.A(net1144),
    .B(_03337_),
    .Y(_03602_));
 sky130_fd_sc_hd__a22o_1 _08104_ (.A1(net1144),
    .A2(_03600_),
    .B1(_03601_),
    .B2(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__xor2_1 _08105_ (.A(_03336_),
    .B(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__nor2_1 _08106_ (.A(_03465_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__a211o_1 _08107_ (.A1(_03336_),
    .A2(net928),
    .B1(_03599_),
    .C1(_03605_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__o21a_1 _08108_ (.A1(_03328_),
    .A2(net931),
    .B1(net969),
    .X(_03606_));
 sky130_fd_sc_hd__a2bb2o_1 _08109_ (.A1_N(_03329_),
    .A2_N(_03606_),
    .B1(net933),
    .B2(_03328_),
    .X(_03607_));
 sky130_fd_sc_hd__nand2_1 _08110_ (.A(_03336_),
    .B(_03339_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21a_1 _08111_ (.A1(net1159),
    .A2(net1013),
    .B1(_03337_),
    .X(_03609_));
 sky130_fd_sc_hd__a21oi_1 _08112_ (.A1(net1159),
    .A2(net1013),
    .B1(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__o21a_1 _08113_ (.A1(_03593_),
    .A2(_03608_),
    .B1(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__inv_2 _08114_ (.A(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__o21a_1 _08115_ (.A1(_03348_),
    .A2(_03437_),
    .B1(_03401_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _08116_ (.A0(_03612_),
    .A1(_03613_),
    .S(net1143),
    .X(_03614_));
 sky130_fd_sc_hd__nand2_1 _08117_ (.A(_03330_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__o21a_1 _08118_ (.A1(_03330_),
    .A2(_03614_),
    .B1(net771),
    .X(_03616_));
 sky130_fd_sc_hd__a21o_1 _08119_ (.A1(_03615_),
    .A2(_03616_),
    .B1(_03607_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__nor2_1 _08120_ (.A(_03332_),
    .B(net935),
    .Y(_03617_));
 sky130_fd_sc_hd__a221o_1 _08121_ (.A1(net966),
    .A2(_03331_),
    .B1(_03333_),
    .B2(net929),
    .C1(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__nor2_1 _08122_ (.A(_03330_),
    .B(_03613_),
    .Y(_03619_));
 sky130_fd_sc_hd__o21ai_1 _08123_ (.A1(_03402_),
    .A2(_03619_),
    .B1(net1144),
    .Y(_03620_));
 sky130_fd_sc_hd__nor2_1 _08124_ (.A(_03329_),
    .B(_03611_),
    .Y(_03621_));
 sky130_fd_sc_hd__o31a_1 _08125_ (.A1(net1144),
    .A2(_03328_),
    .A3(_03621_),
    .B1(_03620_),
    .X(_03622_));
 sky130_fd_sc_hd__xnor2_1 _08126_ (.A(_03334_),
    .B(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__a21o_1 _08127_ (.A1(_03464_),
    .A2(_03623_),
    .B1(_03618_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__nand2_1 _08128_ (.A(_03319_),
    .B(net932),
    .Y(_03624_));
 sky130_fd_sc_hd__o221a_1 _08129_ (.A1(net969),
    .A2(_03321_),
    .B1(_03324_),
    .B2(net931),
    .C1(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__nand2_1 _08130_ (.A(_03330_),
    .B(_03333_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand2b_1 _08131_ (.A_N(_03328_),
    .B(_03332_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand2_1 _08132_ (.A(_03331_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__o21ai_1 _08133_ (.A1(_03611_),
    .A2(_03626_),
    .B1(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__a21oi_1 _08134_ (.A1(_03334_),
    .A2(_03619_),
    .B1(_03404_),
    .Y(_03630_));
 sky130_fd_sc_hd__mux2_1 _08135_ (.A0(_03629_),
    .A1(_03630_),
    .S(net1144),
    .X(_03631_));
 sky130_fd_sc_hd__xnor2_1 _08136_ (.A(_03323_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__o21ai_2 _08137_ (.A1(_03465_),
    .A2(_03632_),
    .B1(_03625_),
    .Y(\alu_out[22] ));
 sky130_fd_sc_hd__nor2_1 _08138_ (.A(_03325_),
    .B(net935),
    .Y(_03633_));
 sky130_fd_sc_hd__a221o_1 _08139_ (.A1(net966),
    .A2(_03326_),
    .B1(_03327_),
    .B2(net929),
    .C1(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__o21ba_1 _08140_ (.A1(_03323_),
    .A2(_03630_),
    .B1_N(_03405_),
    .X(_03635_));
 sky130_fd_sc_hd__a21o_1 _08141_ (.A1(_03322_),
    .A2(_03629_),
    .B1(_03319_),
    .X(_03636_));
 sky130_fd_sc_hd__mux2_1 _08142_ (.A0(_03635_),
    .A1(_03636_),
    .S(_02364_),
    .X(_03637_));
 sky130_fd_sc_hd__or2_1 _08143_ (.A(_03327_),
    .B(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__nand2_1 _08144_ (.A(_03327_),
    .B(_03637_),
    .Y(_03639_));
 sky130_fd_sc_hd__a31o_1 _08145_ (.A1(_03464_),
    .A2(_03638_),
    .A3(_03639_),
    .B1(_03634_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__nor2_1 _08146_ (.A(_03292_),
    .B(net931),
    .Y(_03640_));
 sky130_fd_sc_hd__o21ba_1 _08147_ (.A1(net966),
    .A2(_03640_),
    .B1_N(_03293_),
    .X(_03641_));
 sky130_fd_sc_hd__o21a_1 _08148_ (.A1(_03592_),
    .A2(_03608_),
    .B1(_03610_),
    .X(_03642_));
 sky130_fd_sc_hd__and2_1 _08149_ (.A(_03323_),
    .B(_03327_),
    .X(_03643_));
 sky130_fd_sc_hd__nand2_1 _08150_ (.A(_03320_),
    .B(_03325_),
    .Y(_03644_));
 sky130_fd_sc_hd__o21ai_1 _08151_ (.A1(_03626_),
    .A2(_03642_),
    .B1(_03628_),
    .Y(_03645_));
 sky130_fd_sc_hd__a22o_1 _08152_ (.A1(_03326_),
    .A2(_03644_),
    .B1(_03645_),
    .B2(_03643_),
    .X(_03646_));
 sky130_fd_sc_hd__nor2_1 _08153_ (.A(_03608_),
    .B(_03626_),
    .Y(_03647_));
 sky130_fd_sc_hd__a31o_1 _08154_ (.A1(_03590_),
    .A2(_03643_),
    .A3(_03647_),
    .B1(_03646_),
    .X(_03648_));
 sky130_fd_sc_hd__mux2_1 _08155_ (.A0(_03438_),
    .A1(_03648_),
    .S(net990),
    .X(_03649_));
 sky130_fd_sc_hd__o21ai_1 _08156_ (.A1(_03294_),
    .A2(_03649_),
    .B1(net771),
    .Y(_03650_));
 sky130_fd_sc_hd__a21oi_1 _08157_ (.A1(_03294_),
    .A2(_03649_),
    .B1(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__a211o_1 _08158_ (.A1(_03292_),
    .A2(net933),
    .B1(_03641_),
    .C1(_03651_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__o2bb2a_1 _08159_ (.A1_N(net966),
    .A2_N(_03269_),
    .B1(_03270_),
    .B2(net935),
    .X(_03652_));
 sky130_fd_sc_hd__o21a_1 _08160_ (.A1(_03272_),
    .A2(net931),
    .B1(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__a211o_1 _08161_ (.A1(_02396_),
    .A2(net1004),
    .B1(_03439_),
    .C1(net990),
    .X(_03654_));
 sky130_fd_sc_hd__nor2_1 _08162_ (.A(_03292_),
    .B(_03648_),
    .Y(_03655_));
 sky130_fd_sc_hd__o31a_1 _08163_ (.A1(net1145),
    .A2(_03293_),
    .A3(_03655_),
    .B1(_03654_),
    .X(_03656_));
 sky130_fd_sc_hd__nor2_1 _08164_ (.A(_03272_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__a21o_1 _08165_ (.A1(_03272_),
    .A2(_03656_),
    .B1(_03465_),
    .X(_03658_));
 sky130_fd_sc_hd__o21ai_1 _08166_ (.A1(_03657_),
    .A2(_03658_),
    .B1(_03653_),
    .Y(\alu_out[25] ));
 sky130_fd_sc_hd__nor2_1 _08167_ (.A(_03295_),
    .B(net935),
    .Y(_03659_));
 sky130_fd_sc_hd__a221o_1 _08168_ (.A1(net966),
    .A2(_03296_),
    .B1(_03297_),
    .B2(net929),
    .C1(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__and3_1 _08169_ (.A(_03271_),
    .B(_03294_),
    .C(_03648_),
    .X(_03661_));
 sky130_fd_sc_hd__a21o_1 _08170_ (.A1(net252),
    .A2(net1002),
    .B1(_03292_),
    .X(_03662_));
 sky130_fd_sc_hd__a21o_1 _08171_ (.A1(_03269_),
    .A2(_03662_),
    .B1(_03661_),
    .X(_03663_));
 sky130_fd_sc_hd__mux2_1 _08172_ (.A0(_03442_),
    .A1(_03663_),
    .S(net990),
    .X(_03664_));
 sky130_fd_sc_hd__o21ai_1 _08173_ (.A1(_03297_),
    .A2(_03664_),
    .B1(_03464_),
    .Y(_03665_));
 sky130_fd_sc_hd__a21oi_1 _08174_ (.A1(_03297_),
    .A2(_03664_),
    .B1(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__or2_1 _08175_ (.A(_03660_),
    .B(_03666_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__nor2_1 _08176_ (.A(_03289_),
    .B(net935),
    .Y(_03667_));
 sky130_fd_sc_hd__a221o_1 _08177_ (.A1(net966),
    .A2(_03290_),
    .B1(_03291_),
    .B2(net929),
    .C1(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__a21bo_1 _08178_ (.A1(_03296_),
    .A2(_03663_),
    .B1_N(_03295_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _08179_ (.A0(_03443_),
    .A1(_03669_),
    .S(net990),
    .X(_03670_));
 sky130_fd_sc_hd__or2_1 _08180_ (.A(_03291_),
    .B(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__nand2_1 _08181_ (.A(_03291_),
    .B(_03670_),
    .Y(_03672_));
 sky130_fd_sc_hd__a31o_1 _08182_ (.A1(net771),
    .A2(_03671_),
    .A3(_03672_),
    .B1(_03668_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__a21o_1 _08183_ (.A1(_03266_),
    .A2(net929),
    .B1(net966),
    .X(_03673_));
 sky130_fd_sc_hd__nand2_1 _08184_ (.A(_03289_),
    .B(_03295_),
    .Y(_03674_));
 sky130_fd_sc_hd__a32oi_2 _08185_ (.A1(_03291_),
    .A2(_03297_),
    .A3(_03663_),
    .B1(_03674_),
    .B2(_03290_),
    .Y(_03675_));
 sky130_fd_sc_hd__or3_1 _08186_ (.A(net990),
    .B(_03444_),
    .C(_03446_),
    .X(_03676_));
 sky130_fd_sc_hd__o21ai_1 _08187_ (.A1(net1145),
    .A2(_03675_),
    .B1(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__xnor2_1 _08188_ (.A(_03268_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__a2bb2o_1 _08189_ (.A1_N(_03266_),
    .A2_N(net935),
    .B1(net771),
    .B2(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__a21o_1 _08190_ (.A1(_03267_),
    .A2(_03673_),
    .B1(_03679_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__a21o_1 _08191_ (.A1(_03312_),
    .A2(net929),
    .B1(net966),
    .X(_03680_));
 sky130_fd_sc_hd__o2bb2a_1 _08192_ (.A1_N(_03313_),
    .A2_N(_03680_),
    .B1(net935),
    .B2(_03312_),
    .X(_03681_));
 sky130_fd_sc_hd__a21bo_1 _08193_ (.A1(_03266_),
    .A2(_03675_),
    .B1_N(_03267_),
    .X(_03682_));
 sky130_fd_sc_hd__a21o_1 _08194_ (.A1(_02399_),
    .A2(net997),
    .B1(net990),
    .X(_03683_));
 sky130_fd_sc_hd__o22a_1 _08195_ (.A1(net1145),
    .A2(_03682_),
    .B1(_03683_),
    .B2(_03447_),
    .X(_03684_));
 sky130_fd_sc_hd__xnor2_1 _08196_ (.A(_03314_),
    .B(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__o21ai_2 _08197_ (.A1(_03465_),
    .A2(_03685_),
    .B1(_03681_),
    .Y(\alu_out[29] ));
 sky130_fd_sc_hd__o21a_1 _08198_ (.A1(_03370_),
    .A2(net931),
    .B1(net969),
    .X(_03686_));
 sky130_fd_sc_hd__nor2_1 _08199_ (.A(_03371_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__a21bo_1 _08200_ (.A1(_03312_),
    .A2(_03682_),
    .B1_N(_03313_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _08201_ (.A0(_03449_),
    .A1(_03688_),
    .S(net990),
    .X(_03689_));
 sky130_fd_sc_hd__a21oi_1 _08202_ (.A1(_03372_),
    .A2(_03689_),
    .B1(_03465_),
    .Y(_03690_));
 sky130_fd_sc_hd__o21a_1 _08203_ (.A1(_03372_),
    .A2(_03689_),
    .B1(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__a211o_1 _08204_ (.A1(_03370_),
    .A2(net933),
    .B1(_03687_),
    .C1(_03691_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__nor2_1 _08205_ (.A(_03366_),
    .B(net935),
    .Y(_03692_));
 sky130_fd_sc_hd__a221o_1 _08206_ (.A1(net966),
    .A2(_03367_),
    .B1(_03368_),
    .B2(net929),
    .C1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__nand2_1 _08207_ (.A(_03372_),
    .B(_03449_),
    .Y(_03694_));
 sky130_fd_sc_hd__a21o_1 _08208_ (.A1(_03394_),
    .A2(_03694_),
    .B1(net990),
    .X(_03695_));
 sky130_fd_sc_hd__nor2_1 _08209_ (.A(_03371_),
    .B(_03688_),
    .Y(_03696_));
 sky130_fd_sc_hd__o31a_1 _08210_ (.A1(net1145),
    .A2(_03370_),
    .A3(_03696_),
    .B1(_03695_),
    .X(_03697_));
 sky130_fd_sc_hd__or2_1 _08211_ (.A(_03368_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__a21oi_1 _08212_ (.A1(_03368_),
    .A2(_03697_),
    .B1(_03465_),
    .Y(_03699_));
 sky130_fd_sc_hd__a21o_1 _08213_ (.A1(_03698_),
    .A2(_03699_),
    .B1(_03693_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__a22o_4 _08214_ (.A1(_02383_),
    .A2(net1053),
    .B1(_02689_),
    .B2(net942),
    .X(net131));
 sky130_fd_sc_hd__a211o_2 _08215_ (.A1(net1050),
    .A2(_02384_),
    .B1(_02688_),
    .C1(net940),
    .X(net132));
 sky130_fd_sc_hd__a211o_2 _08216_ (.A1(net1050),
    .A2(net1053),
    .B1(_02688_),
    .C1(net940),
    .X(net133));
 sky130_fd_sc_hd__a22o_1 _08217_ (.A1(net1181),
    .A2(net1056),
    .B1(net265),
    .B2(net1054),
    .X(_03700_));
 sky130_fd_sc_hd__a22o_1 _08218_ (.A1(net1180),
    .A2(net1059),
    .B1(net1168),
    .B2(net942),
    .X(net127));
 sky130_fd_sc_hd__a22o_1 _08219_ (.A1(net1058),
    .A2(net1179),
    .B1(net266),
    .B2(net1054),
    .X(_03701_));
 sky130_fd_sc_hd__a22o_1 _08220_ (.A1(net1059),
    .A2(net1178),
    .B1(net1167),
    .B2(net942),
    .X(net128));
 sky130_fd_sc_hd__a22o_1 _08221_ (.A1(net1056),
    .A2(net1177),
    .B1(net236),
    .B2(net1055),
    .X(_03702_));
 sky130_fd_sc_hd__a22o_1 _08222_ (.A1(net1056),
    .A2(net1177),
    .B1(net236),
    .B2(net942),
    .X(net98));
 sky130_fd_sc_hd__a22o_1 _08223_ (.A1(net1058),
    .A2(net1176),
    .B1(net237),
    .B2(net1055),
    .X(_03703_));
 sky130_fd_sc_hd__a22o_1 _08224_ (.A1(net1059),
    .A2(net1176),
    .B1(net1165),
    .B2(net942),
    .X(net99));
 sky130_fd_sc_hd__a22o_1 _08225_ (.A1(net1058),
    .A2(net1175),
    .B1(net238),
    .B2(net1055),
    .X(_03704_));
 sky130_fd_sc_hd__a22o_1 _08226_ (.A1(net1059),
    .A2(net1174),
    .B1(net1164),
    .B2(net942),
    .X(net100));
 sky130_fd_sc_hd__a22o_1 _08227_ (.A1(net1056),
    .A2(net1173),
    .B1(net239),
    .B2(net1054),
    .X(_03705_));
 sky130_fd_sc_hd__a22o_1 _08228_ (.A1(net1056),
    .A2(net1173),
    .B1(net239),
    .B2(net942),
    .X(net101));
 sky130_fd_sc_hd__a22o_1 _08229_ (.A1(net1056),
    .A2(net1171),
    .B1(net240),
    .B2(net1055),
    .X(_03706_));
 sky130_fd_sc_hd__a22o_2 _08230_ (.A1(net1056),
    .A2(net1171),
    .B1(net240),
    .B2(net942),
    .X(net102));
 sky130_fd_sc_hd__a22o_1 _08231_ (.A1(net1056),
    .A2(net1170),
    .B1(net1162),
    .B2(net1055),
    .X(_03707_));
 sky130_fd_sc_hd__a22o_1 _08232_ (.A1(net1056),
    .A2(net1169),
    .B1(net1162),
    .B2(_02690_),
    .X(net103));
 sky130_fd_sc_hd__mux2_1 _08233_ (.A0(net1180),
    .A1(net1161),
    .S(net940),
    .X(net104));
 sky130_fd_sc_hd__mux2_1 _08234_ (.A0(net1178),
    .A1(net1160),
    .S(net940),
    .X(net105));
 sky130_fd_sc_hd__mux2_1 _08235_ (.A0(net1177),
    .A1(net244),
    .S(net940),
    .X(net106));
 sky130_fd_sc_hd__mux2_1 _08236_ (.A0(net1176),
    .A1(net1159),
    .S(net940),
    .X(net107));
 sky130_fd_sc_hd__mux2_1 _08237_ (.A0(net1175),
    .A1(net247),
    .S(net940),
    .X(net109));
 sky130_fd_sc_hd__mux2_1 _08238_ (.A0(net1172),
    .A1(net248),
    .S(net940),
    .X(net110));
 sky130_fd_sc_hd__mux2_1 _08239_ (.A0(net1171),
    .A1(net1158),
    .S(net940),
    .X(net111));
 sky130_fd_sc_hd__mux2_1 _08240_ (.A0(net1170),
    .A1(net250),
    .S(net941),
    .X(net112));
 sky130_fd_sc_hd__a21o_1 _08241_ (.A1(net251),
    .A2(net941),
    .B1(_03700_),
    .X(net113));
 sky130_fd_sc_hd__a21o_1 _08242_ (.A1(net252),
    .A2(net941),
    .B1(_03701_),
    .X(net114));
 sky130_fd_sc_hd__a21o_1 _08243_ (.A1(net253),
    .A2(net941),
    .B1(_03702_),
    .X(net115));
 sky130_fd_sc_hd__a21o_1 _08244_ (.A1(net254),
    .A2(net941),
    .B1(_03703_),
    .X(net116));
 sky130_fd_sc_hd__a21o_1 _08245_ (.A1(net255),
    .A2(net941),
    .B1(_03704_),
    .X(net117));
 sky130_fd_sc_hd__a21o_1 _08246_ (.A1(net256),
    .A2(net941),
    .B1(_03705_),
    .X(net118));
 sky130_fd_sc_hd__a21o_1 _08247_ (.A1(net258),
    .A2(net941),
    .B1(_03706_),
    .X(net120));
 sky130_fd_sc_hd__a21o_1 _08248_ (.A1(net1157),
    .A2(net940),
    .B1(_03707_),
    .X(net121));
 sky130_fd_sc_hd__nand2_1 _08249_ (.A(latched_branch),
    .B(latched_store),
    .Y(_03708_));
 sky130_fd_sc_hd__mux2_1 _08250_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(net923),
    .X(_03709_));
 sky130_fd_sc_hd__mux2_4 _08251_ (.A0(net1045),
    .A1(_03709_),
    .S(net981),
    .X(net86));
 sky130_fd_sc_hd__mux2_1 _08252_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(net922),
    .X(_03710_));
 sky130_fd_sc_hd__mux2_2 _08253_ (.A0(net1044),
    .A1(_03710_),
    .S(net981),
    .X(net89));
 sky130_fd_sc_hd__mux2_1 _08254_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(net923),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_2 _08255_ (.A0(net1042),
    .A1(_03711_),
    .S(net981),
    .X(net90));
 sky130_fd_sc_hd__mux2_1 _08256_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(net923),
    .X(_03712_));
 sky130_fd_sc_hd__mux2_2 _08257_ (.A0(net1040),
    .A1(_03712_),
    .S(net980),
    .X(net91));
 sky130_fd_sc_hd__mux2_1 _08258_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(net921),
    .X(_03713_));
 sky130_fd_sc_hd__mux2_2 _08259_ (.A0(net1038),
    .A1(_03713_),
    .S(net980),
    .X(net92));
 sky130_fd_sc_hd__mux2_1 _08260_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(net921),
    .X(_03714_));
 sky130_fd_sc_hd__mux2_2 _08261_ (.A0(net1035),
    .A1(_03714_),
    .S(net980),
    .X(net93));
 sky130_fd_sc_hd__mux2_1 _08262_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(net921),
    .X(_03715_));
 sky130_fd_sc_hd__mux2_1 _08263_ (.A0(net1033),
    .A1(_03715_),
    .S(net980),
    .X(net94));
 sky130_fd_sc_hd__mux2_1 _08264_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(net921),
    .X(_03716_));
 sky130_fd_sc_hd__mux2_1 _08265_ (.A0(net1031),
    .A1(_03716_),
    .S(net980),
    .X(net95));
 sky130_fd_sc_hd__mux2_1 _08266_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(net921),
    .X(_03717_));
 sky130_fd_sc_hd__mux2_1 _08267_ (.A0(net1029),
    .A1(_03717_),
    .S(net981),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _08268_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(net920),
    .X(_03718_));
 sky130_fd_sc_hd__mux2_1 _08269_ (.A0(net1028),
    .A1(_03718_),
    .S(net980),
    .X(net67));
 sky130_fd_sc_hd__mux2_1 _08270_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(net920),
    .X(_03719_));
 sky130_fd_sc_hd__mux2_1 _08271_ (.A0(net1026),
    .A1(_03719_),
    .S(net980),
    .X(net68));
 sky130_fd_sc_hd__mux2_1 _08272_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(net920),
    .X(_03720_));
 sky130_fd_sc_hd__mux2_1 _08273_ (.A0(net1024),
    .A1(_03720_),
    .S(net980),
    .X(net69));
 sky130_fd_sc_hd__mux2_1 _08274_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(net920),
    .X(_03721_));
 sky130_fd_sc_hd__mux2_1 _08275_ (.A0(net1022),
    .A1(_03721_),
    .S(net980),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _08276_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(net921),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_2 _08277_ (.A0(net1020),
    .A1(_03722_),
    .S(net980),
    .X(net71));
 sky130_fd_sc_hd__mux2_1 _08278_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(net922),
    .X(_03723_));
 sky130_fd_sc_hd__mux2_2 _08279_ (.A0(net1018),
    .A1(_03723_),
    .S(net981),
    .X(net72));
 sky130_fd_sc_hd__mux2_1 _08280_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(net922),
    .X(_03724_));
 sky130_fd_sc_hd__mux2_2 _08281_ (.A0(net1017),
    .A1(_03724_),
    .S(net981),
    .X(net73));
 sky130_fd_sc_hd__mux2_1 _08282_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(net922),
    .X(_03725_));
 sky130_fd_sc_hd__mux2_2 _08283_ (.A0(net1014),
    .A1(_03725_),
    .S(net981),
    .X(net74));
 sky130_fd_sc_hd__mux2_1 _08284_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(net922),
    .X(_03726_));
 sky130_fd_sc_hd__mux2_2 _08285_ (.A0(net1012),
    .A1(_03726_),
    .S(net981),
    .X(net75));
 sky130_fd_sc_hd__mux2_1 _08286_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(net926),
    .X(_03727_));
 sky130_fd_sc_hd__mux2_2 _08287_ (.A0(net1010),
    .A1(_03727_),
    .S(net981),
    .X(net76));
 sky130_fd_sc_hd__mux2_1 _08288_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(net926),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_2 _08289_ (.A0(net1009),
    .A1(_03728_),
    .S(net982),
    .X(net77));
 sky130_fd_sc_hd__mux2_1 _08290_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(net926),
    .X(_03729_));
 sky130_fd_sc_hd__mux2_2 _08291_ (.A0(net1007),
    .A1(_03729_),
    .S(net982),
    .X(net78));
 sky130_fd_sc_hd__mux2_1 _08292_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(net926),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_2 _08293_ (.A0(net1006),
    .A1(_03730_),
    .S(net982),
    .X(net79));
 sky130_fd_sc_hd__mux2_1 _08294_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(net925),
    .X(_03731_));
 sky130_fd_sc_hd__mux2_2 _08295_ (.A0(net1004),
    .A1(_03731_),
    .S(net982),
    .X(net80));
 sky130_fd_sc_hd__mux2_1 _08296_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(net925),
    .X(_03732_));
 sky130_fd_sc_hd__mux2_1 _08297_ (.A0(net1002),
    .A1(_03732_),
    .S(net982),
    .X(net81));
 sky130_fd_sc_hd__mux2_1 _08298_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(net924),
    .X(_03733_));
 sky130_fd_sc_hd__mux2_2 _08299_ (.A0(net1000),
    .A1(_03733_),
    .S(net982),
    .X(net82));
 sky130_fd_sc_hd__mux2_1 _08300_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(net925),
    .X(_03734_));
 sky130_fd_sc_hd__mux2_2 _08301_ (.A0(net998),
    .A1(_03734_),
    .S(net983),
    .X(net83));
 sky130_fd_sc_hd__mux2_1 _08302_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(net925),
    .X(_03735_));
 sky130_fd_sc_hd__mux2_2 _08303_ (.A0(net996),
    .A1(_03735_),
    .S(net982),
    .X(net84));
 sky130_fd_sc_hd__mux2_1 _08304_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(net924),
    .X(_03736_));
 sky130_fd_sc_hd__mux2_1 _08305_ (.A0(net994),
    .A1(_03736_),
    .S(net982),
    .X(net85));
 sky130_fd_sc_hd__mux2_1 _08306_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(net924),
    .X(_03737_));
 sky130_fd_sc_hd__mux2_1 _08307_ (.A0(net992),
    .A1(_03737_),
    .S(net982),
    .X(net87));
 sky130_fd_sc_hd__mux2_1 _08308_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(net924),
    .X(_03738_));
 sky130_fd_sc_hd__mux2_2 _08309_ (.A0(net1188),
    .A1(_03738_),
    .S(net983),
    .X(net88));
 sky130_fd_sc_hd__nor2_1 _08310_ (.A(net991),
    .B(_03456_),
    .Y(_03739_));
 sky130_fd_sc_hd__nor2_1 _08311_ (.A(_02486_),
    .B(_03456_),
    .Y(_03740_));
 sky130_fd_sc_hd__nor2_1 _08312_ (.A(_02369_),
    .B(_02452_),
    .Y(_03741_));
 sky130_fd_sc_hd__o2bb2a_1 _08313_ (.A1_N(net961),
    .A2_N(_03740_),
    .B1(net548),
    .B2(_00814_),
    .X(_00000_));
 sky130_fd_sc_hd__or3b_1 _08314_ (.A(\latched_rd[2] ),
    .B(\latched_rd[3] ),
    .C_N(\latched_rd[4] ),
    .X(_03742_));
 sky130_fd_sc_hd__o21ai_4 _08315_ (.A1(latched_branch),
    .A2(latched_store),
    .B1(net850),
    .Y(_03743_));
 sky130_fd_sc_hd__or3_1 _08316_ (.A(\latched_rd[2] ),
    .B(\latched_rd[4] ),
    .C(\latched_rd[3] ),
    .X(_03744_));
 sky130_fd_sc_hd__or3b_4 _08317_ (.A(\latched_rd[0] ),
    .B(_03743_),
    .C_N(\latched_rd[1] ),
    .X(_03745_));
 sky130_fd_sc_hd__or2_4 _08318_ (.A(_03742_),
    .B(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__or2_4 _08319_ (.A(latched_branch),
    .B(_02368_),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_1 _08320_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(net1155),
    .X(_03748_));
 sky130_fd_sc_hd__and2b_2 _08321_ (.A_N(net768),
    .B(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__mux2_1 _08322_ (.A0(net587),
    .A1(net2216),
    .S(net530),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _08323_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(net1154),
    .X(_03750_));
 sky130_fd_sc_hd__mux2_4 _08324_ (.A0(_03750_),
    .A1(\reg_pc[1] ),
    .S(net768),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_1 _08325_ (.A0(net584),
    .A1(net2523),
    .S(net530),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _08326_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(net1154),
    .X(_03752_));
 sky130_fd_sc_hd__mux2_2 _08327_ (.A0(_03752_),
    .A1(_02371_),
    .S(net767),
    .X(_03753_));
 sky130_fd_sc_hd__mux2_1 _08328_ (.A0(net581),
    .A1(net2206),
    .S(net531),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _08329_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(net1154),
    .X(_03754_));
 sky130_fd_sc_hd__xor2_1 _08330_ (.A(\reg_pc[3] ),
    .B(\reg_pc[2] ),
    .X(_03755_));
 sky130_fd_sc_hd__mux2_2 _08331_ (.A0(_03754_),
    .A1(_03755_),
    .S(net767),
    .X(_03756_));
 sky130_fd_sc_hd__mux2_1 _08332_ (.A0(net577),
    .A1(net2474),
    .S(net528),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _08333_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(net1154),
    .X(_03757_));
 sky130_fd_sc_hd__and3_1 _08334_ (.A(\reg_pc[4] ),
    .B(\reg_pc[3] ),
    .C(\reg_pc[2] ),
    .X(_03758_));
 sky130_fd_sc_hd__a21oi_1 _08335_ (.A1(\reg_pc[3] ),
    .A2(\reg_pc[2] ),
    .B1(\reg_pc[4] ),
    .Y(_03759_));
 sky130_fd_sc_hd__nor2_1 _08336_ (.A(_03758_),
    .B(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__mux2_2 _08337_ (.A0(_03757_),
    .A1(_03760_),
    .S(net767),
    .X(_03761_));
 sky130_fd_sc_hd__mux2_1 _08338_ (.A0(net573),
    .A1(net2440),
    .S(net531),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _08339_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(net1154),
    .X(_03762_));
 sky130_fd_sc_hd__nor2_1 _08340_ (.A(\reg_pc[5] ),
    .B(_03758_),
    .Y(_03763_));
 sky130_fd_sc_hd__and2_1 _08341_ (.A(\reg_pc[5] ),
    .B(_03758_),
    .X(_03764_));
 sky130_fd_sc_hd__nor2_1 _08342_ (.A(_03763_),
    .B(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__mux2_1 _08343_ (.A0(_03762_),
    .A1(_03765_),
    .S(net767),
    .X(_03766_));
 sky130_fd_sc_hd__mux2_1 _08344_ (.A0(net542),
    .A1(net2537),
    .S(net528),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _08345_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(net1153),
    .X(_03767_));
 sky130_fd_sc_hd__xor2_1 _08346_ (.A(\reg_pc[6] ),
    .B(_03764_),
    .X(_03768_));
 sky130_fd_sc_hd__mux2_1 _08347_ (.A0(_03767_),
    .A1(_03768_),
    .S(net766),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_1 _08348_ (.A0(net539),
    .A1(net2279),
    .S(net528),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _08349_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(net1153),
    .X(_03770_));
 sky130_fd_sc_hd__a21oi_1 _08350_ (.A1(\reg_pc[6] ),
    .A2(_03764_),
    .B1(\reg_pc[7] ),
    .Y(_03771_));
 sky130_fd_sc_hd__and3_1 _08351_ (.A(\reg_pc[7] ),
    .B(\reg_pc[6] ),
    .C(_03764_),
    .X(_03772_));
 sky130_fd_sc_hd__nor2_1 _08352_ (.A(_03771_),
    .B(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__mux2_4 _08353_ (.A0(_03770_),
    .A1(_03773_),
    .S(net766),
    .X(_03774_));
 sky130_fd_sc_hd__mux2_1 _08354_ (.A0(net524),
    .A1(net2309),
    .S(net529),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _08355_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(net1153),
    .X(_03775_));
 sky130_fd_sc_hd__xor2_1 _08356_ (.A(\reg_pc[8] ),
    .B(_03772_),
    .X(_03776_));
 sky130_fd_sc_hd__mux2_1 _08357_ (.A0(_03775_),
    .A1(_03776_),
    .S(net766),
    .X(_03777_));
 sky130_fd_sc_hd__mux2_1 _08358_ (.A0(net520),
    .A1(net2366),
    .S(net529),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _08359_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(net1153),
    .X(_03778_));
 sky130_fd_sc_hd__a21oi_1 _08360_ (.A1(\reg_pc[8] ),
    .A2(_03772_),
    .B1(\reg_pc[9] ),
    .Y(_03779_));
 sky130_fd_sc_hd__and3_1 _08361_ (.A(\reg_pc[9] ),
    .B(\reg_pc[8] ),
    .C(_03772_),
    .X(_03780_));
 sky130_fd_sc_hd__nor2_1 _08362_ (.A(_03779_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__mux2_1 _08363_ (.A0(_03778_),
    .A1(_03781_),
    .S(net766),
    .X(_03782_));
 sky130_fd_sc_hd__mux2_1 _08364_ (.A0(net409),
    .A1(net2182),
    .S(net529),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _08365_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(net1153),
    .X(_03783_));
 sky130_fd_sc_hd__xor2_1 _08366_ (.A(\reg_pc[10] ),
    .B(_03780_),
    .X(_03784_));
 sky130_fd_sc_hd__mux2_2 _08367_ (.A0(_03783_),
    .A1(_03784_),
    .S(net766),
    .X(_03785_));
 sky130_fd_sc_hd__mux2_1 _08368_ (.A0(net405),
    .A1(net2156),
    .S(net529),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _08369_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(net1153),
    .X(_03786_));
 sky130_fd_sc_hd__a21oi_1 _08370_ (.A1(\reg_pc[10] ),
    .A2(_03780_),
    .B1(\reg_pc[11] ),
    .Y(_03787_));
 sky130_fd_sc_hd__and3_1 _08371_ (.A(\reg_pc[11] ),
    .B(\reg_pc[10] ),
    .C(_03780_),
    .X(_03788_));
 sky130_fd_sc_hd__and3_1 _08372_ (.A(\reg_pc[11] ),
    .B(\reg_pc[10] ),
    .C(_03780_),
    .X(_03789_));
 sky130_fd_sc_hd__nor2_1 _08373_ (.A(_03787_),
    .B(_03788_),
    .Y(_03790_));
 sky130_fd_sc_hd__mux2_1 _08374_ (.A0(_03786_),
    .A1(_03790_),
    .S(net766),
    .X(_03791_));
 sky130_fd_sc_hd__mux2_1 _08375_ (.A0(net355),
    .A1(net2452),
    .S(net529),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _08376_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(net1153),
    .X(_03792_));
 sky130_fd_sc_hd__xor2_1 _08377_ (.A(\reg_pc[12] ),
    .B(_03788_),
    .X(_03793_));
 sky130_fd_sc_hd__mux2_1 _08378_ (.A0(_03792_),
    .A1(_03793_),
    .S(net766),
    .X(_03794_));
 sky130_fd_sc_hd__mux2_1 _08379_ (.A0(net351),
    .A1(net2370),
    .S(net528),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _08380_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(net1153),
    .X(_03795_));
 sky130_fd_sc_hd__a21oi_1 _08381_ (.A1(\reg_pc[12] ),
    .A2(_03788_),
    .B1(\reg_pc[13] ),
    .Y(_03796_));
 sky130_fd_sc_hd__and3_1 _08382_ (.A(\reg_pc[13] ),
    .B(\reg_pc[12] ),
    .C(_03789_),
    .X(_03797_));
 sky130_fd_sc_hd__nor2_1 _08383_ (.A(_03796_),
    .B(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__mux2_2 _08384_ (.A0(_03795_),
    .A1(_03798_),
    .S(net766),
    .X(_03799_));
 sky130_fd_sc_hd__mux2_1 _08385_ (.A0(net347),
    .A1(net2210),
    .S(net528),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _08386_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(net1153),
    .X(_03800_));
 sky130_fd_sc_hd__xor2_1 _08387_ (.A(\reg_pc[14] ),
    .B(_03797_),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_2 _08388_ (.A0(_03800_),
    .A1(_03801_),
    .S(net766),
    .X(_03802_));
 sky130_fd_sc_hd__mux2_1 _08389_ (.A0(net343),
    .A1(net2388),
    .S(net529),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _08390_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(net1153),
    .X(_03803_));
 sky130_fd_sc_hd__a21oi_1 _08391_ (.A1(\reg_pc[14] ),
    .A2(_03797_),
    .B1(\reg_pc[15] ),
    .Y(_03804_));
 sky130_fd_sc_hd__and3_1 _08392_ (.A(\reg_pc[15] ),
    .B(\reg_pc[14] ),
    .C(_03797_),
    .X(_03805_));
 sky130_fd_sc_hd__nor2_1 _08393_ (.A(_03804_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__mux2_4 _08394_ (.A0(_03803_),
    .A1(_03806_),
    .S(net766),
    .X(_03807_));
 sky130_fd_sc_hd__mux2_1 _08395_ (.A0(net339),
    .A1(net2204),
    .S(net528),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _08396_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(net1154),
    .X(_03808_));
 sky130_fd_sc_hd__xor2_1 _08397_ (.A(\reg_pc[16] ),
    .B(_03805_),
    .X(_03809_));
 sky130_fd_sc_hd__mux2_2 _08398_ (.A0(_03808_),
    .A1(_03809_),
    .S(net767),
    .X(_03810_));
 sky130_fd_sc_hd__mux2_1 _08399_ (.A0(net336),
    .A1(net2315),
    .S(net528),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _08400_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(net1154),
    .X(_03811_));
 sky130_fd_sc_hd__a21oi_1 _08401_ (.A1(\reg_pc[16] ),
    .A2(_03805_),
    .B1(\reg_pc[17] ),
    .Y(_03812_));
 sky130_fd_sc_hd__and3_1 _08402_ (.A(\reg_pc[17] ),
    .B(\reg_pc[16] ),
    .C(_03805_),
    .X(_03813_));
 sky130_fd_sc_hd__nor2_1 _08403_ (.A(_03812_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__mux2_2 _08404_ (.A0(_03811_),
    .A1(_03814_),
    .S(net767),
    .X(_03815_));
 sky130_fd_sc_hd__mux2_1 _08405_ (.A0(net332),
    .A1(net2131),
    .S(net528),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _08406_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(net1154),
    .X(_03816_));
 sky130_fd_sc_hd__xor2_1 _08407_ (.A(\reg_pc[18] ),
    .B(_03813_),
    .X(_03817_));
 sky130_fd_sc_hd__mux2_4 _08408_ (.A0(_03816_),
    .A1(_03817_),
    .S(net767),
    .X(_03818_));
 sky130_fd_sc_hd__mux2_1 _08409_ (.A0(net328),
    .A1(net2379),
    .S(net528),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _08410_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(net1154),
    .X(_03819_));
 sky130_fd_sc_hd__a21oi_1 _08411_ (.A1(\reg_pc[18] ),
    .A2(_03813_),
    .B1(\reg_pc[19] ),
    .Y(_03820_));
 sky130_fd_sc_hd__and3_1 _08412_ (.A(\reg_pc[19] ),
    .B(\reg_pc[18] ),
    .C(_03813_),
    .X(_03821_));
 sky130_fd_sc_hd__nor2_1 _08413_ (.A(_03820_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__mux2_1 _08414_ (.A0(_03819_),
    .A1(_03822_),
    .S(net767),
    .X(_03823_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(net324),
    .A1(net2450),
    .S(net530),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _08416_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(net1155),
    .X(_03824_));
 sky130_fd_sc_hd__xor2_1 _08417_ (.A(\reg_pc[20] ),
    .B(_03821_),
    .X(_03825_));
 sky130_fd_sc_hd__mux2_4 _08418_ (.A0(_03824_),
    .A1(_03825_),
    .S(net768),
    .X(_03826_));
 sky130_fd_sc_hd__mux2_1 _08419_ (.A0(net321),
    .A1(net2475),
    .S(net528),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _08420_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(net1155),
    .X(_03827_));
 sky130_fd_sc_hd__a21oi_1 _08421_ (.A1(\reg_pc[20] ),
    .A2(_03821_),
    .B1(\reg_pc[21] ),
    .Y(_03828_));
 sky130_fd_sc_hd__and3_1 _08422_ (.A(\reg_pc[21] ),
    .B(\reg_pc[20] ),
    .C(_03821_),
    .X(_03829_));
 sky130_fd_sc_hd__nor2_1 _08423_ (.A(_03828_),
    .B(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__mux2_1 _08424_ (.A0(_03827_),
    .A1(_03830_),
    .S(net768),
    .X(_03831_));
 sky130_fd_sc_hd__mux2_1 _08425_ (.A0(net316),
    .A1(net2146),
    .S(net530),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _08426_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(net1155),
    .X(_03832_));
 sky130_fd_sc_hd__nor2_1 _08427_ (.A(\reg_pc[22] ),
    .B(_03829_),
    .Y(_03833_));
 sky130_fd_sc_hd__and2_1 _08428_ (.A(\reg_pc[22] ),
    .B(_03829_),
    .X(_03834_));
 sky130_fd_sc_hd__nor2_1 _08429_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__mux2_1 _08430_ (.A0(_03832_),
    .A1(_03835_),
    .S(net768),
    .X(_03836_));
 sky130_fd_sc_hd__mux2_1 _08431_ (.A0(net313),
    .A1(net2222),
    .S(net530),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _08432_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(net1155),
    .X(_03837_));
 sky130_fd_sc_hd__xor2_1 _08433_ (.A(\reg_pc[23] ),
    .B(_03834_),
    .X(_03838_));
 sky130_fd_sc_hd__mux2_1 _08434_ (.A0(_03837_),
    .A1(_03838_),
    .S(net768),
    .X(_03839_));
 sky130_fd_sc_hd__mux2_1 _08435_ (.A0(net311),
    .A1(net2406),
    .S(net530),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _08436_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(net1156),
    .X(_03840_));
 sky130_fd_sc_hd__a21oi_1 _08437_ (.A1(\reg_pc[23] ),
    .A2(_03834_),
    .B1(\reg_pc[24] ),
    .Y(_03841_));
 sky130_fd_sc_hd__and3_1 _08438_ (.A(\reg_pc[24] ),
    .B(\reg_pc[23] ),
    .C(_03834_),
    .X(_03842_));
 sky130_fd_sc_hd__nor2_1 _08439_ (.A(_03841_),
    .B(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__mux2_2 _08440_ (.A0(_03840_),
    .A1(_03843_),
    .S(net768),
    .X(_03844_));
 sky130_fd_sc_hd__mux2_1 _08441_ (.A0(net306),
    .A1(net2331),
    .S(net531),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _08442_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(net1155),
    .X(_03845_));
 sky130_fd_sc_hd__nor2_1 _08443_ (.A(\reg_pc[25] ),
    .B(_03842_),
    .Y(_03846_));
 sky130_fd_sc_hd__and2_1 _08444_ (.A(\reg_pc[25] ),
    .B(_03842_),
    .X(_03847_));
 sky130_fd_sc_hd__nor2_1 _08445_ (.A(_03846_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__mux2_1 _08446_ (.A0(_03845_),
    .A1(_03848_),
    .S(net769),
    .X(_03849_));
 sky130_fd_sc_hd__mux2_1 _08447_ (.A0(net301),
    .A1(net2247),
    .S(net531),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _08448_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(net1155),
    .X(_03850_));
 sky130_fd_sc_hd__xor2_1 _08449_ (.A(\reg_pc[26] ),
    .B(_03847_),
    .X(_03851_));
 sky130_fd_sc_hd__mux2_2 _08450_ (.A0(_03850_),
    .A1(_03851_),
    .S(net768),
    .X(_03852_));
 sky130_fd_sc_hd__mux2_1 _08451_ (.A0(net297),
    .A1(net2217),
    .S(net531),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _08452_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(net1155),
    .X(_03853_));
 sky130_fd_sc_hd__a21oi_1 _08453_ (.A1(\reg_pc[26] ),
    .A2(_03847_),
    .B1(\reg_pc[27] ),
    .Y(_03854_));
 sky130_fd_sc_hd__and3_1 _08454_ (.A(\reg_pc[27] ),
    .B(\reg_pc[26] ),
    .C(_03847_),
    .X(_03855_));
 sky130_fd_sc_hd__nor2_1 _08455_ (.A(_03854_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__mux2_2 _08456_ (.A0(_03853_),
    .A1(_03856_),
    .S(net768),
    .X(_03857_));
 sky130_fd_sc_hd__mux2_1 _08457_ (.A0(net293),
    .A1(net2458),
    .S(net530),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _08458_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(net1155),
    .X(_03858_));
 sky130_fd_sc_hd__xor2_1 _08459_ (.A(\reg_pc[28] ),
    .B(_03855_),
    .X(_03859_));
 sky130_fd_sc_hd__mux2_2 _08460_ (.A0(_03858_),
    .A1(_03859_),
    .S(net768),
    .X(_03860_));
 sky130_fd_sc_hd__mux2_1 _08461_ (.A0(net289),
    .A1(net2531),
    .S(net530),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _08462_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(net1155),
    .X(_03861_));
 sky130_fd_sc_hd__a21oi_1 _08463_ (.A1(\reg_pc[28] ),
    .A2(_03855_),
    .B1(\reg_pc[29] ),
    .Y(_03862_));
 sky130_fd_sc_hd__and3_1 _08464_ (.A(\reg_pc[29] ),
    .B(\reg_pc[28] ),
    .C(_03855_),
    .X(_03863_));
 sky130_fd_sc_hd__nor2_1 _08465_ (.A(_03862_),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__mux2_1 _08466_ (.A0(_03861_),
    .A1(_03864_),
    .S(net769),
    .X(_03865_));
 sky130_fd_sc_hd__mux2_1 _08467_ (.A0(net285),
    .A1(net2493),
    .S(net531),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _08468_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(net1156),
    .X(_03866_));
 sky130_fd_sc_hd__or2_1 _08469_ (.A(\reg_pc[30] ),
    .B(_03863_),
    .X(_03867_));
 sky130_fd_sc_hd__nand2_1 _08470_ (.A(\reg_pc[30] ),
    .B(_03863_),
    .Y(_03868_));
 sky130_fd_sc_hd__and2b_1 _08471_ (.A_N(net769),
    .B(_03866_),
    .X(_03869_));
 sky130_fd_sc_hd__a31o_2 _08472_ (.A1(net769),
    .A2(_03867_),
    .A3(_03868_),
    .B1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__mux2_1 _08473_ (.A0(net283),
    .A1(net2305),
    .S(net530),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _08474_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(net1156),
    .X(_03871_));
 sky130_fd_sc_hd__xnor2_1 _08475_ (.A(\reg_pc[31] ),
    .B(_03868_),
    .Y(_03872_));
 sky130_fd_sc_hd__mux2_2 _08476_ (.A0(_03871_),
    .A1(_03872_),
    .S(net769),
    .X(_03873_));
 sky130_fd_sc_hd__mux2_1 _08477_ (.A0(net278),
    .A1(net2506),
    .S(net530),
    .X(_00081_));
 sky130_fd_sc_hd__and2_1 _08478_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1237),
    .X(_03874_));
 sky130_fd_sc_hd__nand2_1 _08479_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1223),
    .Y(_03875_));
 sky130_fd_sc_hd__and3_1 _08480_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1189),
    .C(net1237),
    .X(_03876_));
 sky130_fd_sc_hd__o21a_1 _08481_ (.A1(\genblk1.genblk1.pcpi_mul.instr_mulhsu ),
    .A2(\genblk1.genblk1.pcpi_mul.instr_mulh ),
    .B1(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__a21o_1 _08482_ (.A1(net1215),
    .A2(net1582),
    .B1(net762),
    .X(_00082_));
 sky130_fd_sc_hd__a22o_1 _08483_ (.A1(net1199),
    .A2(net2759),
    .B1(net916),
    .B2(net1181),
    .X(_00083_));
 sky130_fd_sc_hd__nand3_1 _08484_ (.A(\genblk1.genblk1.pcpi_mul.rd[0] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[1] ),
    .C(net1101),
    .Y(_03878_));
 sky130_fd_sc_hd__nor2_2 _08485_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1216),
    .Y(_03879_));
 sky130_fd_sc_hd__a21o_1 _08486_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[1] ),
    .A2(net1102),
    .B1(\genblk1.genblk1.pcpi_mul.rd[0] ),
    .X(_03880_));
 sky130_fd_sc_hd__a32o_1 _08487_ (.A1(_03878_),
    .A2(net894),
    .A3(_03880_),
    .B1(net2681),
    .B2(net1199),
    .X(_00084_));
 sky130_fd_sc_hd__a21oi_1 _08488_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[2] ),
    .A2(net1101),
    .B1(\genblk1.genblk1.pcpi_mul.rd[1] ),
    .Y(_03881_));
 sky130_fd_sc_hd__and3_1 _08489_ (.A(\genblk1.genblk1.pcpi_mul.rd[1] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[2] ),
    .C(net1101),
    .X(_03882_));
 sky130_fd_sc_hd__nor3_1 _08490_ (.A(_03878_),
    .B(_03881_),
    .C(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__inv_2 _08491_ (.A(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__o21ai_1 _08492_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03878_),
    .Y(_03885_));
 sky130_fd_sc_hd__a32o_1 _08493_ (.A1(net896),
    .A2(_03884_),
    .A3(_03885_),
    .B1(net2614),
    .B2(net1199),
    .X(_00085_));
 sky130_fd_sc_hd__a21o_1 _08494_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[3] ),
    .A2(net1098),
    .B1(\genblk1.genblk1.pcpi_mul.rd[2] ),
    .X(_03886_));
 sky130_fd_sc_hd__nand3_1 _08495_ (.A(\genblk1.genblk1.pcpi_mul.rd[2] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[3] ),
    .C(net1098),
    .Y(_03887_));
 sky130_fd_sc_hd__a211o_1 _08496_ (.A1(_03886_),
    .A2(_03887_),
    .B1(_03882_),
    .C1(net761),
    .X(_03888_));
 sky130_fd_sc_hd__o211a_1 _08497_ (.A1(_03882_),
    .A2(net761),
    .B1(_03886_),
    .C1(_03887_),
    .X(_03889_));
 sky130_fd_sc_hd__inv_2 _08498_ (.A(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__a32o_1 _08499_ (.A1(net894),
    .A2(_03888_),
    .A3(_03890_),
    .B1(net2624),
    .B2(net1199),
    .X(_00086_));
 sky130_fd_sc_hd__nand3_1 _08500_ (.A(\genblk1.genblk1.pcpi_mul.rd[3] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[4] ),
    .C(net1098),
    .Y(_03891_));
 sky130_fd_sc_hd__a21o_1 _08501_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[4] ),
    .A2(net1098),
    .B1(\genblk1.genblk1.pcpi_mul.rd[3] ),
    .X(_03892_));
 sky130_fd_sc_hd__nand2_1 _08502_ (.A(_03891_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_1 _08503_ (.A(_03887_),
    .B(_03890_),
    .Y(_03894_));
 sky130_fd_sc_hd__xnor2_1 _08504_ (.A(_03893_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__a22o_1 _08505_ (.A1(net1199),
    .A2(net2872),
    .B1(net894),
    .B2(_03895_),
    .X(_00087_));
 sky130_fd_sc_hd__nand2_1 _08506_ (.A(\genblk1.genblk1.pcpi_mul.rd[4] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[4] ),
    .Y(_03896_));
 sky130_fd_sc_hd__inv_2 _08507_ (.A(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__or2_1 _08508_ (.A(\genblk1.genblk1.pcpi_mul.rd[4] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[4] ),
    .X(_03898_));
 sky130_fd_sc_hd__a22o_1 _08509_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[5] ),
    .A2(net1098),
    .B1(_03896_),
    .B2(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__and4_1 _08510_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[5] ),
    .B(net1098),
    .C(_03896_),
    .D(_03898_),
    .X(_03900_));
 sky130_fd_sc_hd__inv_2 _08511_ (.A(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__a32o_1 _08512_ (.A1(net893),
    .A2(_03899_),
    .A3(_03901_),
    .B1(net2604),
    .B2(net1200),
    .X(_00088_));
 sky130_fd_sc_hd__a21o_1 _08513_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[6] ),
    .A2(net1096),
    .B1(\genblk1.genblk1.pcpi_mul.rd[5] ),
    .X(_03902_));
 sky130_fd_sc_hd__and3_1 _08514_ (.A(\genblk1.genblk1.pcpi_mul.rd[5] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[6] ),
    .C(net1097),
    .X(_03903_));
 sky130_fd_sc_hd__nand3_1 _08515_ (.A(\genblk1.genblk1.pcpi_mul.rd[5] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[6] ),
    .C(net1096),
    .Y(_03904_));
 sky130_fd_sc_hd__a211o_1 _08516_ (.A1(_03902_),
    .A2(_03904_),
    .B1(_03897_),
    .C1(_03900_),
    .X(_03905_));
 sky130_fd_sc_hd__o211a_1 _08517_ (.A1(_03897_),
    .A2(_03900_),
    .B1(_03902_),
    .C1(_03904_),
    .X(_03906_));
 sky130_fd_sc_hd__inv_2 _08518_ (.A(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__a32o_1 _08519_ (.A1(net892),
    .A2(_03905_),
    .A3(_03907_),
    .B1(net2773),
    .B2(net1201),
    .X(_00089_));
 sky130_fd_sc_hd__a21o_1 _08520_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[7] ),
    .A2(net1097),
    .B1(\genblk1.genblk1.pcpi_mul.rd[6] ),
    .X(_03908_));
 sky130_fd_sc_hd__nand3_1 _08521_ (.A(\genblk1.genblk1.pcpi_mul.rd[6] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[7] ),
    .C(net1097),
    .Y(_03909_));
 sky130_fd_sc_hd__a211o_1 _08522_ (.A1(_03908_),
    .A2(_03909_),
    .B1(_03903_),
    .C1(_03906_),
    .X(_03910_));
 sky130_fd_sc_hd__o211a_1 _08523_ (.A1(_03903_),
    .A2(_03906_),
    .B1(_03908_),
    .C1(_03909_),
    .X(_03911_));
 sky130_fd_sc_hd__inv_2 _08524_ (.A(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__a32o_1 _08525_ (.A1(net892),
    .A2(_03910_),
    .A3(_03912_),
    .B1(net2659),
    .B2(net1201),
    .X(_00090_));
 sky130_fd_sc_hd__nand3_1 _08526_ (.A(\genblk1.genblk1.pcpi_mul.rd[7] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[8] ),
    .C(net1095),
    .Y(_03913_));
 sky130_fd_sc_hd__a21o_1 _08527_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[8] ),
    .A2(net1095),
    .B1(\genblk1.genblk1.pcpi_mul.rd[7] ),
    .X(_03914_));
 sky130_fd_sc_hd__nand2_1 _08528_ (.A(_03913_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(_03909_),
    .B(_03912_),
    .Y(_03916_));
 sky130_fd_sc_hd__xnor2_1 _08530_ (.A(_03915_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__a22o_1 _08531_ (.A1(net1195),
    .A2(net2883),
    .B1(net888),
    .B2(_03917_),
    .X(_00091_));
 sky130_fd_sc_hd__nand2_1 _08532_ (.A(\genblk1.genblk1.pcpi_mul.rd[8] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[8] ),
    .Y(_03918_));
 sky130_fd_sc_hd__inv_2 _08533_ (.A(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__or2_1 _08534_ (.A(\genblk1.genblk1.pcpi_mul.rd[8] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[8] ),
    .X(_03920_));
 sky130_fd_sc_hd__a22o_1 _08535_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[9] ),
    .A2(net1094),
    .B1(_03918_),
    .B2(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__and4_1 _08536_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[9] ),
    .B(net1095),
    .C(_03918_),
    .D(_03920_),
    .X(_03922_));
 sky130_fd_sc_hd__inv_2 _08537_ (.A(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__a32o_1 _08538_ (.A1(net887),
    .A2(_03921_),
    .A3(_03923_),
    .B1(net2592),
    .B2(net1193),
    .X(_00092_));
 sky130_fd_sc_hd__a21o_1 _08539_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[10] ),
    .A2(net1095),
    .B1(\genblk1.genblk1.pcpi_mul.rd[9] ),
    .X(_03924_));
 sky130_fd_sc_hd__and3_1 _08540_ (.A(\genblk1.genblk1.pcpi_mul.rd[9] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[10] ),
    .C(net1091),
    .X(_03925_));
 sky130_fd_sc_hd__nand3_1 _08541_ (.A(\genblk1.genblk1.pcpi_mul.rd[9] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[10] ),
    .C(net1092),
    .Y(_03926_));
 sky130_fd_sc_hd__a211o_1 _08542_ (.A1(_03924_),
    .A2(_03926_),
    .B1(_03919_),
    .C1(_03922_),
    .X(_03927_));
 sky130_fd_sc_hd__o211a_1 _08543_ (.A1(_03919_),
    .A2(_03922_),
    .B1(_03924_),
    .C1(_03926_),
    .X(_03928_));
 sky130_fd_sc_hd__inv_2 _08544_ (.A(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__a32o_1 _08545_ (.A1(net887),
    .A2(_03927_),
    .A3(_03929_),
    .B1(net2749),
    .B2(net1193),
    .X(_00093_));
 sky130_fd_sc_hd__a21o_1 _08546_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[11] ),
    .A2(net1091),
    .B1(\genblk1.genblk1.pcpi_mul.rd[10] ),
    .X(_03930_));
 sky130_fd_sc_hd__nand3_1 _08547_ (.A(\genblk1.genblk1.pcpi_mul.rd[10] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[11] ),
    .C(net1092),
    .Y(_03931_));
 sky130_fd_sc_hd__a211o_1 _08548_ (.A1(_03930_),
    .A2(_03931_),
    .B1(_03925_),
    .C1(_03928_),
    .X(_03932_));
 sky130_fd_sc_hd__o211a_1 _08549_ (.A1(_03925_),
    .A2(_03928_),
    .B1(_03930_),
    .C1(_03931_),
    .X(_03933_));
 sky130_fd_sc_hd__inv_2 _08550_ (.A(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__a32o_1 _08551_ (.A1(net887),
    .A2(_03932_),
    .A3(_03934_),
    .B1(net2628),
    .B2(net1197),
    .X(_00094_));
 sky130_fd_sc_hd__nand3_1 _08552_ (.A(\genblk1.genblk1.pcpi_mul.rd[11] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[12] ),
    .C(net1091),
    .Y(_03935_));
 sky130_fd_sc_hd__a21o_1 _08553_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[12] ),
    .A2(net1091),
    .B1(\genblk1.genblk1.pcpi_mul.rd[11] ),
    .X(_03936_));
 sky130_fd_sc_hd__nand2_1 _08554_ (.A(_03935_),
    .B(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _08555_ (.A(_03931_),
    .B(_03934_),
    .Y(_03938_));
 sky130_fd_sc_hd__xnor2_1 _08556_ (.A(_03937_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__a22o_1 _08557_ (.A1(net1193),
    .A2(net2911),
    .B1(net886),
    .B2(_03939_),
    .X(_00095_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(\genblk1.genblk1.pcpi_mul.rd[12] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[12] ),
    .Y(_03940_));
 sky130_fd_sc_hd__inv_2 _08559_ (.A(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__or2_1 _08560_ (.A(\genblk1.genblk1.pcpi_mul.rd[12] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[12] ),
    .X(_03942_));
 sky130_fd_sc_hd__a22o_1 _08561_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[13] ),
    .A2(net1090),
    .B1(_03940_),
    .B2(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__and4_1 _08562_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[13] ),
    .B(net1090),
    .C(_03940_),
    .D(_03942_),
    .X(_03944_));
 sky130_fd_sc_hd__inv_2 _08563_ (.A(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__a32o_1 _08564_ (.A1(net885),
    .A2(_03943_),
    .A3(_03945_),
    .B1(net2574),
    .B2(net1192),
    .X(_00096_));
 sky130_fd_sc_hd__a21o_1 _08565_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[14] ),
    .A2(net1093),
    .B1(\genblk1.genblk1.pcpi_mul.rd[13] ),
    .X(_03946_));
 sky130_fd_sc_hd__and3_1 _08566_ (.A(\genblk1.genblk1.pcpi_mul.rd[13] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[14] ),
    .C(net1093),
    .X(_03947_));
 sky130_fd_sc_hd__nand3_1 _08567_ (.A(\genblk1.genblk1.pcpi_mul.rd[13] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[14] ),
    .C(net1093),
    .Y(_03948_));
 sky130_fd_sc_hd__a211o_1 _08568_ (.A1(_03946_),
    .A2(_03948_),
    .B1(_03941_),
    .C1(_03944_),
    .X(_03949_));
 sky130_fd_sc_hd__o211a_1 _08569_ (.A1(_03941_),
    .A2(_03944_),
    .B1(_03946_),
    .C1(_03948_),
    .X(_03950_));
 sky130_fd_sc_hd__inv_2 _08570_ (.A(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__a32o_1 _08571_ (.A1(net885),
    .A2(_03949_),
    .A3(_03951_),
    .B1(net2765),
    .B2(net1192),
    .X(_00097_));
 sky130_fd_sc_hd__a21o_1 _08572_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[15] ),
    .A2(net1090),
    .B1(\genblk1.genblk1.pcpi_mul.rd[14] ),
    .X(_03952_));
 sky130_fd_sc_hd__nand3_1 _08573_ (.A(\genblk1.genblk1.pcpi_mul.rd[14] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[15] ),
    .C(net1090),
    .Y(_03953_));
 sky130_fd_sc_hd__a211o_1 _08574_ (.A1(_03952_),
    .A2(_03953_),
    .B1(_03947_),
    .C1(_03950_),
    .X(_03954_));
 sky130_fd_sc_hd__o211a_1 _08575_ (.A1(_03947_),
    .A2(_03950_),
    .B1(_03952_),
    .C1(_03953_),
    .X(_03955_));
 sky130_fd_sc_hd__inv_2 _08576_ (.A(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__a32o_1 _08577_ (.A1(net891),
    .A2(_03954_),
    .A3(_03956_),
    .B1(net2626),
    .B2(net1192),
    .X(_00098_));
 sky130_fd_sc_hd__nand3_1 _08578_ (.A(\genblk1.genblk1.pcpi_mul.rd[15] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[16] ),
    .C(net1094),
    .Y(_03957_));
 sky130_fd_sc_hd__a21o_1 _08579_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[16] ),
    .A2(net1094),
    .B1(\genblk1.genblk1.pcpi_mul.rd[15] ),
    .X(_03958_));
 sky130_fd_sc_hd__nand2_1 _08580_ (.A(_03957_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__nand2_1 _08581_ (.A(_03953_),
    .B(_03956_),
    .Y(_03960_));
 sky130_fd_sc_hd__xnor2_1 _08582_ (.A(_03959_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__a22o_1 _08583_ (.A1(net1196),
    .A2(net2880),
    .B1(net890),
    .B2(_03961_),
    .X(_00099_));
 sky130_fd_sc_hd__nand2_1 _08584_ (.A(\genblk1.genblk1.pcpi_mul.rd[16] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[16] ),
    .Y(_03962_));
 sky130_fd_sc_hd__inv_2 _08585_ (.A(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__or2_1 _08586_ (.A(\genblk1.genblk1.pcpi_mul.rd[16] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[16] ),
    .X(_03964_));
 sky130_fd_sc_hd__a22o_1 _08587_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[17] ),
    .A2(net1094),
    .B1(_03962_),
    .B2(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__and4_1 _08588_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[17] ),
    .B(net1094),
    .C(_03962_),
    .D(_03964_),
    .X(_03966_));
 sky130_fd_sc_hd__inv_2 _08589_ (.A(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__a32o_1 _08590_ (.A1(net890),
    .A2(_03965_),
    .A3(_03967_),
    .B1(net2567),
    .B2(net1196),
    .X(_00100_));
 sky130_fd_sc_hd__a21o_1 _08591_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[18] ),
    .A2(net1100),
    .B1(\genblk1.genblk1.pcpi_mul.rd[17] ),
    .X(_03968_));
 sky130_fd_sc_hd__and3_1 _08592_ (.A(\genblk1.genblk1.pcpi_mul.rd[17] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[18] ),
    .C(net1096),
    .X(_03969_));
 sky130_fd_sc_hd__nand3_1 _08593_ (.A(\genblk1.genblk1.pcpi_mul.rd[17] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[18] ),
    .C(net1100),
    .Y(_03970_));
 sky130_fd_sc_hd__a211o_1 _08594_ (.A1(_03968_),
    .A2(_03970_),
    .B1(_03963_),
    .C1(_03966_),
    .X(_03971_));
 sky130_fd_sc_hd__o211a_1 _08595_ (.A1(_03963_),
    .A2(_03966_),
    .B1(_03968_),
    .C1(_03970_),
    .X(_03972_));
 sky130_fd_sc_hd__inv_2 _08596_ (.A(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__a32o_1 _08597_ (.A1(net890),
    .A2(_03971_),
    .A3(_03973_),
    .B1(net2838),
    .B2(net1196),
    .X(_00101_));
 sky130_fd_sc_hd__a21o_1 _08598_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[19] ),
    .A2(net1097),
    .B1(\genblk1.genblk1.pcpi_mul.rd[18] ),
    .X(_03974_));
 sky130_fd_sc_hd__nand3_1 _08599_ (.A(\genblk1.genblk1.pcpi_mul.rd[18] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[19] ),
    .C(net1097),
    .Y(_03975_));
 sky130_fd_sc_hd__a211o_1 _08600_ (.A1(_03974_),
    .A2(_03975_),
    .B1(_03969_),
    .C1(_03972_),
    .X(_03976_));
 sky130_fd_sc_hd__o211a_1 _08601_ (.A1(_03969_),
    .A2(_03972_),
    .B1(_03974_),
    .C1(_03975_),
    .X(_03977_));
 sky130_fd_sc_hd__inv_2 _08602_ (.A(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__a32o_1 _08603_ (.A1(net892),
    .A2(_03976_),
    .A3(_03978_),
    .B1(net2632),
    .B2(net1200),
    .X(_00102_));
 sky130_fd_sc_hd__nand3_1 _08604_ (.A(\genblk1.genblk1.pcpi_mul.rd[19] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[20] ),
    .C(net1099),
    .Y(_03979_));
 sky130_fd_sc_hd__a21o_1 _08605_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[20] ),
    .A2(net1098),
    .B1(\genblk1.genblk1.pcpi_mul.rd[19] ),
    .X(_03980_));
 sky130_fd_sc_hd__nand2_1 _08606_ (.A(_03979_),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_1 _08607_ (.A(_03975_),
    .B(_03978_),
    .Y(_03982_));
 sky130_fd_sc_hd__xnor2_1 _08608_ (.A(_03981_),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__a22o_1 _08609_ (.A1(net1203),
    .A2(net2888),
    .B1(net895),
    .B2(_03983_),
    .X(_00103_));
 sky130_fd_sc_hd__nand2_1 _08610_ (.A(\genblk1.genblk1.pcpi_mul.rd[20] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[20] ),
    .Y(_03984_));
 sky130_fd_sc_hd__inv_2 _08611_ (.A(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__or2_1 _08612_ (.A(\genblk1.genblk1.pcpi_mul.rd[20] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[20] ),
    .X(_03986_));
 sky130_fd_sc_hd__a22o_1 _08613_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[21] ),
    .A2(net1102),
    .B1(_03984_),
    .B2(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__and4_1 _08614_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[21] ),
    .B(net1102),
    .C(_03984_),
    .D(_03986_),
    .X(_03988_));
 sky130_fd_sc_hd__inv_2 _08615_ (.A(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__a32o_1 _08616_ (.A1(net895),
    .A2(_03987_),
    .A3(_03989_),
    .B1(net2559),
    .B2(net1203),
    .X(_00104_));
 sky130_fd_sc_hd__a21o_1 _08617_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[22] ),
    .A2(net1102),
    .B1(\genblk1.genblk1.pcpi_mul.rd[21] ),
    .X(_03990_));
 sky130_fd_sc_hd__and3_1 _08618_ (.A(\genblk1.genblk1.pcpi_mul.rd[21] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[22] ),
    .C(net1104),
    .X(_03991_));
 sky130_fd_sc_hd__nand3_1 _08619_ (.A(\genblk1.genblk1.pcpi_mul.rd[21] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[22] ),
    .C(net1104),
    .Y(_03992_));
 sky130_fd_sc_hd__a211o_1 _08620_ (.A1(_03990_),
    .A2(_03992_),
    .B1(_03985_),
    .C1(_03988_),
    .X(_03993_));
 sky130_fd_sc_hd__o211a_1 _08621_ (.A1(_03985_),
    .A2(_03988_),
    .B1(_03990_),
    .C1(_03992_),
    .X(_03994_));
 sky130_fd_sc_hd__inv_2 _08622_ (.A(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__a32o_1 _08623_ (.A1(net900),
    .A2(_03993_),
    .A3(_03995_),
    .B1(net2748),
    .B2(net1202),
    .X(_00105_));
 sky130_fd_sc_hd__a21o_1 _08624_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[23] ),
    .A2(net1104),
    .B1(\genblk1.genblk1.pcpi_mul.rd[22] ),
    .X(_03996_));
 sky130_fd_sc_hd__nand3_1 _08625_ (.A(\genblk1.genblk1.pcpi_mul.rd[22] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[23] ),
    .C(net1103),
    .Y(_03997_));
 sky130_fd_sc_hd__a211o_1 _08626_ (.A1(_03996_),
    .A2(_03997_),
    .B1(_03991_),
    .C1(_03994_),
    .X(_03998_));
 sky130_fd_sc_hd__o211a_1 _08627_ (.A1(_03991_),
    .A2(_03994_),
    .B1(_03996_),
    .C1(_03997_),
    .X(_03999_));
 sky130_fd_sc_hd__inv_2 _08628_ (.A(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__a32o_1 _08629_ (.A1(net903),
    .A2(_03998_),
    .A3(_04000_),
    .B1(net2660),
    .B2(net1210),
    .X(_00106_));
 sky130_fd_sc_hd__nand3_1 _08630_ (.A(\genblk1.genblk1.pcpi_mul.rd[23] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[24] ),
    .C(net1103),
    .Y(_04001_));
 sky130_fd_sc_hd__a21o_1 _08631_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[24] ),
    .A2(net1103),
    .B1(\genblk1.genblk1.pcpi_mul.rd[23] ),
    .X(_04002_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__nand2_1 _08633_ (.A(_03997_),
    .B(_04000_),
    .Y(_04004_));
 sky130_fd_sc_hd__xnor2_1 _08634_ (.A(_04003_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__a22o_1 _08635_ (.A1(net1210),
    .A2(net2897),
    .B1(net899),
    .B2(_04005_),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_1 _08636_ (.A(\genblk1.genblk1.pcpi_mul.rd[24] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[24] ),
    .Y(_04006_));
 sky130_fd_sc_hd__inv_2 _08637_ (.A(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__or2_1 _08638_ (.A(\genblk1.genblk1.pcpi_mul.rd[24] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[24] ),
    .X(_04008_));
 sky130_fd_sc_hd__a22o_1 _08639_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[25] ),
    .A2(net1103),
    .B1(_04006_),
    .B2(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__and4_1 _08640_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[25] ),
    .B(net1103),
    .C(_04006_),
    .D(_04008_),
    .X(_04010_));
 sky130_fd_sc_hd__inv_2 _08641_ (.A(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__a32o_1 _08642_ (.A1(net901),
    .A2(_04009_),
    .A3(_04011_),
    .B1(net2587),
    .B2(net1210),
    .X(_00108_));
 sky130_fd_sc_hd__a21o_1 _08643_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[26] ),
    .A2(net1105),
    .B1(\genblk1.genblk1.pcpi_mul.rd[25] ),
    .X(_04012_));
 sky130_fd_sc_hd__and3_1 _08644_ (.A(\genblk1.genblk1.pcpi_mul.rd[25] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[26] ),
    .C(net1105),
    .X(_04013_));
 sky130_fd_sc_hd__nand3_1 _08645_ (.A(\genblk1.genblk1.pcpi_mul.rd[25] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[26] ),
    .C(net1105),
    .Y(_04014_));
 sky130_fd_sc_hd__a211o_1 _08646_ (.A1(_04012_),
    .A2(_04014_),
    .B1(_04007_),
    .C1(_04010_),
    .X(_04015_));
 sky130_fd_sc_hd__o211a_1 _08647_ (.A1(_04007_),
    .A2(_04010_),
    .B1(_04012_),
    .C1(_04014_),
    .X(_04016_));
 sky130_fd_sc_hd__inv_2 _08648_ (.A(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__a32o_1 _08649_ (.A1(net902),
    .A2(_04015_),
    .A3(_04017_),
    .B1(net2781),
    .B2(net1212),
    .X(_00109_));
 sky130_fd_sc_hd__a21o_1 _08650_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[27] ),
    .A2(net1108),
    .B1(\genblk1.genblk1.pcpi_mul.rd[26] ),
    .X(_04018_));
 sky130_fd_sc_hd__nand3_1 _08651_ (.A(\genblk1.genblk1.pcpi_mul.rd[26] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[27] ),
    .C(net1105),
    .Y(_04019_));
 sky130_fd_sc_hd__a211o_1 _08652_ (.A1(_04018_),
    .A2(_04019_),
    .B1(_04013_),
    .C1(_04016_),
    .X(_04020_));
 sky130_fd_sc_hd__o211a_1 _08653_ (.A1(_04013_),
    .A2(_04016_),
    .B1(_04018_),
    .C1(_04019_),
    .X(_04021_));
 sky130_fd_sc_hd__inv_2 _08654_ (.A(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__a32o_1 _08655_ (.A1(net902),
    .A2(_04020_),
    .A3(_04022_),
    .B1(net2683),
    .B2(net1212),
    .X(_00110_));
 sky130_fd_sc_hd__nand3_1 _08656_ (.A(\genblk1.genblk1.pcpi_mul.rd[27] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[28] ),
    .C(net1105),
    .Y(_04023_));
 sky130_fd_sc_hd__a21o_1 _08657_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[28] ),
    .A2(net1105),
    .B1(\genblk1.genblk1.pcpi_mul.rd[27] ),
    .X(_04024_));
 sky130_fd_sc_hd__nand2_1 _08658_ (.A(_04023_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_04019_),
    .B(_04022_),
    .Y(_04026_));
 sky130_fd_sc_hd__xnor2_1 _08660_ (.A(_04025_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__a22o_1 _08661_ (.A1(net1212),
    .A2(net2921),
    .B1(net901),
    .B2(_04027_),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_1 _08662_ (.A(\genblk1.genblk1.pcpi_mul.rd[28] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[28] ),
    .Y(_04028_));
 sky130_fd_sc_hd__inv_2 _08663_ (.A(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__or2_1 _08664_ (.A(\genblk1.genblk1.pcpi_mul.rd[28] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[28] ),
    .X(_04030_));
 sky130_fd_sc_hd__a22o_1 _08665_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[29] ),
    .A2(net1106),
    .B1(_04028_),
    .B2(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__and4_1 _08666_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[29] ),
    .B(net1106),
    .C(_04028_),
    .D(_04030_),
    .X(_04032_));
 sky130_fd_sc_hd__inv_2 _08667_ (.A(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__a32o_1 _08668_ (.A1(net904),
    .A2(_04031_),
    .A3(_04033_),
    .B1(net2577),
    .B2(net1217),
    .X(_00112_));
 sky130_fd_sc_hd__a21o_1 _08669_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[30] ),
    .A2(net1106),
    .B1(\genblk1.genblk1.pcpi_mul.rd[29] ),
    .X(_04034_));
 sky130_fd_sc_hd__and3_1 _08670_ (.A(\genblk1.genblk1.pcpi_mul.rd[29] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[30] ),
    .C(net1106),
    .X(_04035_));
 sky130_fd_sc_hd__nand3_1 _08671_ (.A(\genblk1.genblk1.pcpi_mul.rd[29] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[30] ),
    .C(net1106),
    .Y(_04036_));
 sky130_fd_sc_hd__a211o_1 _08672_ (.A1(_04034_),
    .A2(_04036_),
    .B1(_04029_),
    .C1(_04032_),
    .X(_04037_));
 sky130_fd_sc_hd__o211a_1 _08673_ (.A1(_04029_),
    .A2(_04032_),
    .B1(_04034_),
    .C1(_04036_),
    .X(_04038_));
 sky130_fd_sc_hd__inv_2 _08674_ (.A(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__a32o_1 _08675_ (.A1(net904),
    .A2(_04037_),
    .A3(_04039_),
    .B1(net2789),
    .B2(net1217),
    .X(_00113_));
 sky130_fd_sc_hd__a21o_1 _08676_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[31] ),
    .A2(net1106),
    .B1(\genblk1.genblk1.pcpi_mul.rd[30] ),
    .X(_04040_));
 sky130_fd_sc_hd__nand3_1 _08677_ (.A(\genblk1.genblk1.pcpi_mul.rd[30] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[31] ),
    .C(net1106),
    .Y(_04041_));
 sky130_fd_sc_hd__a211o_1 _08678_ (.A1(_04040_),
    .A2(_04041_),
    .B1(_04035_),
    .C1(_04038_),
    .X(_04042_));
 sky130_fd_sc_hd__o211a_1 _08679_ (.A1(_04035_),
    .A2(_04038_),
    .B1(_04040_),
    .C1(_04041_),
    .X(_04043_));
 sky130_fd_sc_hd__inv_2 _08680_ (.A(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__a32o_1 _08681_ (.A1(net905),
    .A2(_04042_),
    .A3(_04044_),
    .B1(net2696),
    .B2(net1218),
    .X(_00114_));
 sky130_fd_sc_hd__nand3_1 _08682_ (.A(\genblk1.genblk1.pcpi_mul.rd[31] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[32] ),
    .C(net1107),
    .Y(_04045_));
 sky130_fd_sc_hd__a21o_1 _08683_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[32] ),
    .A2(net1107),
    .B1(\genblk1.genblk1.pcpi_mul.rd[31] ),
    .X(_04046_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_04045_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__nand2_1 _08685_ (.A(_04041_),
    .B(_04044_),
    .Y(_04048_));
 sky130_fd_sc_hd__xnor2_1 _08686_ (.A(_04047_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__a22o_1 _08687_ (.A1(net1218),
    .A2(net2919),
    .B1(net905),
    .B2(_04049_),
    .X(_00115_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(\genblk1.genblk1.pcpi_mul.rd[32] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[32] ),
    .Y(_04050_));
 sky130_fd_sc_hd__inv_2 _08689_ (.A(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__or2_1 _08690_ (.A(\genblk1.genblk1.pcpi_mul.rd[32] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[32] ),
    .X(_04052_));
 sky130_fd_sc_hd__a22o_1 _08691_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[33] ),
    .A2(net1101),
    .B1(_04050_),
    .B2(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__and4_1 _08692_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[33] ),
    .B(net1101),
    .C(_04050_),
    .D(_04052_),
    .X(_04054_));
 sky130_fd_sc_hd__inv_2 _08693_ (.A(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__a32o_1 _08694_ (.A1(net899),
    .A2(_04053_),
    .A3(_04055_),
    .B1(net2622),
    .B2(net1202),
    .X(_00116_));
 sky130_fd_sc_hd__a21o_1 _08695_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[34] ),
    .A2(net1101),
    .B1(\genblk1.genblk1.pcpi_mul.rd[33] ),
    .X(_04056_));
 sky130_fd_sc_hd__and3_1 _08696_ (.A(\genblk1.genblk1.pcpi_mul.rd[33] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[34] ),
    .C(net1101),
    .X(_04057_));
 sky130_fd_sc_hd__nand3_1 _08697_ (.A(\genblk1.genblk1.pcpi_mul.rd[33] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[34] ),
    .C(net1101),
    .Y(_04058_));
 sky130_fd_sc_hd__a211o_1 _08698_ (.A1(_04056_),
    .A2(_04058_),
    .B1(_04051_),
    .C1(_04054_),
    .X(_04059_));
 sky130_fd_sc_hd__o211a_1 _08699_ (.A1(_04051_),
    .A2(_04054_),
    .B1(_04056_),
    .C1(_04058_),
    .X(_04060_));
 sky130_fd_sc_hd__inv_2 _08700_ (.A(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__a32o_1 _08701_ (.A1(net894),
    .A2(_04059_),
    .A3(_04061_),
    .B1(net2918),
    .B2(net1202),
    .X(_00117_));
 sky130_fd_sc_hd__a21o_1 _08702_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[35] ),
    .A2(net1101),
    .B1(\genblk1.genblk1.pcpi_mul.rd[34] ),
    .X(_04062_));
 sky130_fd_sc_hd__nand3_1 _08703_ (.A(\genblk1.genblk1.pcpi_mul.rd[34] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[35] ),
    .C(net1101),
    .Y(_04063_));
 sky130_fd_sc_hd__a211o_1 _08704_ (.A1(_04062_),
    .A2(_04063_),
    .B1(_04057_),
    .C1(_04060_),
    .X(_04064_));
 sky130_fd_sc_hd__o211a_1 _08705_ (.A1(_04057_),
    .A2(_04060_),
    .B1(_04062_),
    .C1(_04063_),
    .X(_04065_));
 sky130_fd_sc_hd__inv_2 _08706_ (.A(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__a32o_1 _08707_ (.A1(net894),
    .A2(_04064_),
    .A3(_04066_),
    .B1(net2703),
    .B2(net1202),
    .X(_00118_));
 sky130_fd_sc_hd__nand3_1 _08708_ (.A(\genblk1.genblk1.pcpi_mul.rd[35] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[36] ),
    .C(net1098),
    .Y(_04067_));
 sky130_fd_sc_hd__a21o_1 _08709_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[36] ),
    .A2(net1098),
    .B1(\genblk1.genblk1.pcpi_mul.rd[35] ),
    .X(_04068_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_04067_),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(_04063_),
    .B(_04066_),
    .Y(_04070_));
 sky130_fd_sc_hd__xnor2_1 _08712_ (.A(_04069_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__a22o_1 _08713_ (.A1(net1200),
    .A2(net2931),
    .B1(net894),
    .B2(_04071_),
    .X(_00119_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(\genblk1.genblk1.pcpi_mul.rd[36] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[36] ),
    .Y(_04072_));
 sky130_fd_sc_hd__inv_2 _08715_ (.A(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__or2_1 _08716_ (.A(\genblk1.genblk1.pcpi_mul.rd[36] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[36] ),
    .X(_04074_));
 sky130_fd_sc_hd__a22o_1 _08717_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[37] ),
    .A2(net1099),
    .B1(_04072_),
    .B2(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__and4_1 _08718_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[37] ),
    .B(net1099),
    .C(_04072_),
    .D(_04074_),
    .X(_04076_));
 sky130_fd_sc_hd__inv_2 _08719_ (.A(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__a32o_1 _08720_ (.A1(net893),
    .A2(_04075_),
    .A3(_04077_),
    .B1(net2650),
    .B2(net1201),
    .X(_00120_));
 sky130_fd_sc_hd__a21o_1 _08721_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[38] ),
    .A2(net1099),
    .B1(\genblk1.genblk1.pcpi_mul.rd[37] ),
    .X(_04078_));
 sky130_fd_sc_hd__and3_1 _08722_ (.A(\genblk1.genblk1.pcpi_mul.rd[37] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[38] ),
    .C(net1099),
    .X(_04079_));
 sky130_fd_sc_hd__nand3_1 _08723_ (.A(\genblk1.genblk1.pcpi_mul.rd[37] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[38] ),
    .C(net1099),
    .Y(_04080_));
 sky130_fd_sc_hd__a211o_1 _08724_ (.A1(_04078_),
    .A2(_04080_),
    .B1(_04073_),
    .C1(_04076_),
    .X(_04081_));
 sky130_fd_sc_hd__o211a_1 _08725_ (.A1(_04073_),
    .A2(_04076_),
    .B1(_04078_),
    .C1(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__inv_2 _08726_ (.A(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__a32o_1 _08727_ (.A1(net892),
    .A2(_04081_),
    .A3(_04083_),
    .B1(net2869),
    .B2(net1201),
    .X(_00121_));
 sky130_fd_sc_hd__a21o_1 _08728_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[39] ),
    .A2(net1096),
    .B1(\genblk1.genblk1.pcpi_mul.rd[38] ),
    .X(_04084_));
 sky130_fd_sc_hd__nand3_1 _08729_ (.A(\genblk1.genblk1.pcpi_mul.rd[38] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[39] ),
    .C(net1096),
    .Y(_04085_));
 sky130_fd_sc_hd__a211o_1 _08730_ (.A1(_04084_),
    .A2(_04085_),
    .B1(_04079_),
    .C1(_04082_),
    .X(_04086_));
 sky130_fd_sc_hd__o211a_1 _08731_ (.A1(_04079_),
    .A2(_04082_),
    .B1(_04084_),
    .C1(_04085_),
    .X(_04087_));
 sky130_fd_sc_hd__inv_2 _08732_ (.A(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__a32o_1 _08733_ (.A1(net892),
    .A2(_04086_),
    .A3(_04088_),
    .B1(net2691),
    .B2(net1201),
    .X(_00122_));
 sky130_fd_sc_hd__nand3_1 _08734_ (.A(\genblk1.genblk1.pcpi_mul.rd[39] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[40] ),
    .C(net1094),
    .Y(_04089_));
 sky130_fd_sc_hd__a21o_1 _08735_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[40] ),
    .A2(net1094),
    .B1(\genblk1.genblk1.pcpi_mul.rd[39] ),
    .X(_04090_));
 sky130_fd_sc_hd__nand2_1 _08736_ (.A(_04089_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__nand2_1 _08737_ (.A(_04085_),
    .B(_04088_),
    .Y(_04092_));
 sky130_fd_sc_hd__xnor2_1 _08738_ (.A(_04091_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__a22o_1 _08739_ (.A1(net1197),
    .A2(net2924),
    .B1(net889),
    .B2(_04093_),
    .X(_00123_));
 sky130_fd_sc_hd__nand2_1 _08740_ (.A(\genblk1.genblk1.pcpi_mul.rd[40] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[40] ),
    .Y(_04094_));
 sky130_fd_sc_hd__inv_2 _08741_ (.A(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__or2_1 _08742_ (.A(\genblk1.genblk1.pcpi_mul.rd[40] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[40] ),
    .X(_04096_));
 sky130_fd_sc_hd__a22o_1 _08743_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[41] ),
    .A2(net1091),
    .B1(_04094_),
    .B2(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__and4_1 _08744_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[41] ),
    .B(net1092),
    .C(_04094_),
    .D(_04096_),
    .X(_04098_));
 sky130_fd_sc_hd__inv_2 _08745_ (.A(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__a32o_1 _08746_ (.A1(net887),
    .A2(_04097_),
    .A3(_04099_),
    .B1(net2598),
    .B2(net1197),
    .X(_00124_));
 sky130_fd_sc_hd__a21o_1 _08747_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[42] ),
    .A2(net1092),
    .B1(\genblk1.genblk1.pcpi_mul.rd[41] ),
    .X(_04100_));
 sky130_fd_sc_hd__and3_1 _08748_ (.A(\genblk1.genblk1.pcpi_mul.rd[41] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[42] ),
    .C(net1091),
    .X(_04101_));
 sky130_fd_sc_hd__nand3_1 _08749_ (.A(\genblk1.genblk1.pcpi_mul.rd[41] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[42] ),
    .C(net1092),
    .Y(_04102_));
 sky130_fd_sc_hd__a211o_1 _08750_ (.A1(_04100_),
    .A2(_04102_),
    .B1(_04095_),
    .C1(_04098_),
    .X(_04103_));
 sky130_fd_sc_hd__o211a_1 _08751_ (.A1(_04095_),
    .A2(_04098_),
    .B1(_04100_),
    .C1(_04102_),
    .X(_04104_));
 sky130_fd_sc_hd__inv_2 _08752_ (.A(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__a32o_1 _08753_ (.A1(net886),
    .A2(_04103_),
    .A3(_04105_),
    .B1(net2842),
    .B2(net1193),
    .X(_00125_));
 sky130_fd_sc_hd__a21o_1 _08754_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[43] ),
    .A2(net1091),
    .B1(\genblk1.genblk1.pcpi_mul.rd[42] ),
    .X(_04106_));
 sky130_fd_sc_hd__nand3_1 _08755_ (.A(\genblk1.genblk1.pcpi_mul.rd[42] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[43] ),
    .C(net1091),
    .Y(_04107_));
 sky130_fd_sc_hd__a211o_1 _08756_ (.A1(_04106_),
    .A2(_04107_),
    .B1(_04101_),
    .C1(_04104_),
    .X(_04108_));
 sky130_fd_sc_hd__o211a_1 _08757_ (.A1(_04101_),
    .A2(_04104_),
    .B1(_04106_),
    .C1(_04107_),
    .X(_04109_));
 sky130_fd_sc_hd__inv_2 _08758_ (.A(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__a32o_1 _08759_ (.A1(net886),
    .A2(_04108_),
    .A3(_04110_),
    .B1(net2682),
    .B2(net1193),
    .X(_00126_));
 sky130_fd_sc_hd__nand3_1 _08760_ (.A(\genblk1.genblk1.pcpi_mul.rd[43] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[44] ),
    .C(net1091),
    .Y(_04111_));
 sky130_fd_sc_hd__a21o_1 _08761_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[44] ),
    .A2(net1091),
    .B1(\genblk1.genblk1.pcpi_mul.rd[43] ),
    .X(_04112_));
 sky130_fd_sc_hd__nand2_1 _08762_ (.A(_04111_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand2_1 _08763_ (.A(_04107_),
    .B(_04110_),
    .Y(_04114_));
 sky130_fd_sc_hd__xnor2_1 _08764_ (.A(_04113_),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__a22o_1 _08765_ (.A1(net1193),
    .A2(net2967),
    .B1(net886),
    .B2(_04115_),
    .X(_00127_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(\genblk1.genblk1.pcpi_mul.rd[44] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[44] ),
    .Y(_04116_));
 sky130_fd_sc_hd__inv_2 _08767_ (.A(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__or2_1 _08768_ (.A(\genblk1.genblk1.pcpi_mul.rd[44] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[44] ),
    .X(_04118_));
 sky130_fd_sc_hd__a22o_1 _08769_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[45] ),
    .A2(net1090),
    .B1(_04116_),
    .B2(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__and4_1 _08770_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[45] ),
    .B(net1090),
    .C(_04116_),
    .D(_04118_),
    .X(_04120_));
 sky130_fd_sc_hd__inv_2 _08771_ (.A(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__a32o_1 _08772_ (.A1(net885),
    .A2(_04119_),
    .A3(_04121_),
    .B1(net2676),
    .B2(net1194),
    .X(_00128_));
 sky130_fd_sc_hd__a21o_1 _08773_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[46] ),
    .A2(net1090),
    .B1(\genblk1.genblk1.pcpi_mul.rd[45] ),
    .X(_04122_));
 sky130_fd_sc_hd__and3_1 _08774_ (.A(\genblk1.genblk1.pcpi_mul.rd[45] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[46] ),
    .C(net1093),
    .X(_04123_));
 sky130_fd_sc_hd__nand3_1 _08775_ (.A(\genblk1.genblk1.pcpi_mul.rd[45] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[46] ),
    .C(net1090),
    .Y(_04124_));
 sky130_fd_sc_hd__a211o_1 _08776_ (.A1(_04122_),
    .A2(_04124_),
    .B1(_04117_),
    .C1(_04120_),
    .X(_04125_));
 sky130_fd_sc_hd__o211a_1 _08777_ (.A1(_04117_),
    .A2(_04120_),
    .B1(_04122_),
    .C1(_04124_),
    .X(_04126_));
 sky130_fd_sc_hd__inv_2 _08778_ (.A(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__a32o_1 _08779_ (.A1(net885),
    .A2(_04125_),
    .A3(_04127_),
    .B1(net2871),
    .B2(net1194),
    .X(_00129_));
 sky130_fd_sc_hd__a21o_1 _08780_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[47] ),
    .A2(net1090),
    .B1(\genblk1.genblk1.pcpi_mul.rd[46] ),
    .X(_04128_));
 sky130_fd_sc_hd__nand3_1 _08781_ (.A(\genblk1.genblk1.pcpi_mul.rd[46] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[47] ),
    .C(net1090),
    .Y(_04129_));
 sky130_fd_sc_hd__a211o_1 _08782_ (.A1(_04128_),
    .A2(_04129_),
    .B1(_04123_),
    .C1(_04126_),
    .X(_04130_));
 sky130_fd_sc_hd__o211a_1 _08783_ (.A1(_04123_),
    .A2(_04126_),
    .B1(_04128_),
    .C1(_04129_),
    .X(_04131_));
 sky130_fd_sc_hd__inv_2 _08784_ (.A(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__a32o_1 _08785_ (.A1(net885),
    .A2(_04130_),
    .A3(_04132_),
    .B1(net2697),
    .B2(net1194),
    .X(_00130_));
 sky130_fd_sc_hd__nand3_1 _08786_ (.A(\genblk1.genblk1.pcpi_mul.rd[47] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[48] ),
    .C(net1094),
    .Y(_04133_));
 sky130_fd_sc_hd__a21o_1 _08787_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[48] ),
    .A2(net1095),
    .B1(\genblk1.genblk1.pcpi_mul.rd[47] ),
    .X(_04134_));
 sky130_fd_sc_hd__nand2_1 _08788_ (.A(_04133_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand2_1 _08789_ (.A(_04129_),
    .B(_04132_),
    .Y(_04136_));
 sky130_fd_sc_hd__xnor2_1 _08790_ (.A(_04135_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__a22o_1 _08791_ (.A1(net1196),
    .A2(net2913),
    .B1(net888),
    .B2(_04137_),
    .X(_00131_));
 sky130_fd_sc_hd__nand2_1 _08792_ (.A(\genblk1.genblk1.pcpi_mul.rd[48] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[48] ),
    .Y(_04138_));
 sky130_fd_sc_hd__inv_2 _08793_ (.A(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__or2_1 _08794_ (.A(\genblk1.genblk1.pcpi_mul.rd[48] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[48] ),
    .X(_04140_));
 sky130_fd_sc_hd__a22o_1 _08795_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[49] ),
    .A2(net1094),
    .B1(_04138_),
    .B2(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__and4_1 _08796_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[49] ),
    .B(net1094),
    .C(_04138_),
    .D(_04140_),
    .X(_04142_));
 sky130_fd_sc_hd__inv_2 _08797_ (.A(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__a32o_1 _08798_ (.A1(net889),
    .A2(_04141_),
    .A3(_04143_),
    .B1(net2576),
    .B2(net1195),
    .X(_00132_));
 sky130_fd_sc_hd__a21o_1 _08799_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[50] ),
    .A2(net1096),
    .B1(\genblk1.genblk1.pcpi_mul.rd[49] ),
    .X(_04144_));
 sky130_fd_sc_hd__and3_1 _08800_ (.A(\genblk1.genblk1.pcpi_mul.rd[49] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[50] ),
    .C(net1096),
    .X(_04145_));
 sky130_fd_sc_hd__nand3_1 _08801_ (.A(\genblk1.genblk1.pcpi_mul.rd[49] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[50] ),
    .C(net1096),
    .Y(_04146_));
 sky130_fd_sc_hd__a211o_1 _08802_ (.A1(_04144_),
    .A2(_04146_),
    .B1(_04139_),
    .C1(_04142_),
    .X(_04147_));
 sky130_fd_sc_hd__o211a_1 _08803_ (.A1(_04139_),
    .A2(_04142_),
    .B1(_04144_),
    .C1(_04146_),
    .X(_04148_));
 sky130_fd_sc_hd__inv_2 _08804_ (.A(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__a32o_1 _08805_ (.A1(net889),
    .A2(_04147_),
    .A3(_04149_),
    .B1(net2870),
    .B2(net1197),
    .X(_00133_));
 sky130_fd_sc_hd__a21o_1 _08806_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[51] ),
    .A2(net1096),
    .B1(\genblk1.genblk1.pcpi_mul.rd[50] ),
    .X(_04150_));
 sky130_fd_sc_hd__nand3_1 _08807_ (.A(\genblk1.genblk1.pcpi_mul.rd[50] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[51] ),
    .C(net1096),
    .Y(_04151_));
 sky130_fd_sc_hd__a211o_1 _08808_ (.A1(_04150_),
    .A2(_04151_),
    .B1(_04145_),
    .C1(_04148_),
    .X(_04152_));
 sky130_fd_sc_hd__o211a_1 _08809_ (.A1(_04145_),
    .A2(_04148_),
    .B1(_04150_),
    .C1(_04151_),
    .X(_04153_));
 sky130_fd_sc_hd__inv_2 _08810_ (.A(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__a32o_1 _08811_ (.A1(net892),
    .A2(_04152_),
    .A3(_04154_),
    .B1(net2652),
    .B2(net1195),
    .X(_00134_));
 sky130_fd_sc_hd__nand3_1 _08812_ (.A(\genblk1.genblk1.pcpi_mul.rd[51] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[52] ),
    .C(net1099),
    .Y(_04155_));
 sky130_fd_sc_hd__a21o_1 _08813_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[52] ),
    .A2(net1099),
    .B1(\genblk1.genblk1.pcpi_mul.rd[51] ),
    .X(_04156_));
 sky130_fd_sc_hd__nand2_1 _08814_ (.A(_04155_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand2_1 _08815_ (.A(_04151_),
    .B(_04154_),
    .Y(_04158_));
 sky130_fd_sc_hd__xnor2_1 _08816_ (.A(_04157_),
    .B(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__a22o_1 _08817_ (.A1(net1203),
    .A2(net2995),
    .B1(net895),
    .B2(_04159_),
    .X(_00135_));
 sky130_fd_sc_hd__nand2_1 _08818_ (.A(\genblk1.genblk1.pcpi_mul.rd[52] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[52] ),
    .Y(_04160_));
 sky130_fd_sc_hd__inv_2 _08819_ (.A(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__or2_1 _08820_ (.A(\genblk1.genblk1.pcpi_mul.rd[52] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[52] ),
    .X(_04162_));
 sky130_fd_sc_hd__a22o_1 _08821_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[53] ),
    .A2(net1102),
    .B1(_04160_),
    .B2(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__and4_1 _08822_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[53] ),
    .B(net1102),
    .C(_04160_),
    .D(_04162_),
    .X(_04164_));
 sky130_fd_sc_hd__inv_2 _08823_ (.A(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__a32o_1 _08824_ (.A1(net896),
    .A2(_04163_),
    .A3(_04165_),
    .B1(net2610),
    .B2(net1203),
    .X(_00136_));
 sky130_fd_sc_hd__a21o_1 _08825_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[54] ),
    .A2(net1102),
    .B1(\genblk1.genblk1.pcpi_mul.rd[53] ),
    .X(_04166_));
 sky130_fd_sc_hd__and3_1 _08826_ (.A(\genblk1.genblk1.pcpi_mul.rd[53] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[54] ),
    .C(net1102),
    .X(_04167_));
 sky130_fd_sc_hd__nand3_1 _08827_ (.A(\genblk1.genblk1.pcpi_mul.rd[53] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[54] ),
    .C(net1102),
    .Y(_04168_));
 sky130_fd_sc_hd__a211o_1 _08828_ (.A1(_04166_),
    .A2(_04168_),
    .B1(_04161_),
    .C1(_04164_),
    .X(_04169_));
 sky130_fd_sc_hd__o211a_1 _08829_ (.A1(_04161_),
    .A2(_04164_),
    .B1(_04166_),
    .C1(_04168_),
    .X(_04170_));
 sky130_fd_sc_hd__inv_2 _08830_ (.A(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__a32o_1 _08831_ (.A1(net900),
    .A2(_04169_),
    .A3(_04171_),
    .B1(net2884),
    .B2(net1203),
    .X(_00137_));
 sky130_fd_sc_hd__a21o_1 _08832_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[55] ),
    .A2(net1103),
    .B1(\genblk1.genblk1.pcpi_mul.rd[54] ),
    .X(_04172_));
 sky130_fd_sc_hd__nand3_1 _08833_ (.A(\genblk1.genblk1.pcpi_mul.rd[54] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[55] ),
    .C(net1103),
    .Y(_04173_));
 sky130_fd_sc_hd__a211o_1 _08834_ (.A1(_04172_),
    .A2(_04173_),
    .B1(_04167_),
    .C1(_04170_),
    .X(_04174_));
 sky130_fd_sc_hd__o211a_1 _08835_ (.A1(_04167_),
    .A2(_04170_),
    .B1(_04172_),
    .C1(_04173_),
    .X(_04175_));
 sky130_fd_sc_hd__inv_2 _08836_ (.A(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__a32o_1 _08837_ (.A1(net900),
    .A2(_04174_),
    .A3(_04176_),
    .B1(net2755),
    .B2(net1211),
    .X(_00138_));
 sky130_fd_sc_hd__nand3_1 _08838_ (.A(\genblk1.genblk1.pcpi_mul.rd[55] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[56] ),
    .C(net1103),
    .Y(_04177_));
 sky130_fd_sc_hd__a21o_1 _08839_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[56] ),
    .A2(net1104),
    .B1(\genblk1.genblk1.pcpi_mul.rd[55] ),
    .X(_04178_));
 sky130_fd_sc_hd__nand2_1 _08840_ (.A(_04177_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(_04173_),
    .B(_04176_),
    .Y(_04180_));
 sky130_fd_sc_hd__xnor2_1 _08842_ (.A(_04179_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__a22o_1 _08843_ (.A1(net1211),
    .A2(net2927),
    .B1(net900),
    .B2(_04181_),
    .X(_00139_));
 sky130_fd_sc_hd__nand2_1 _08844_ (.A(\genblk1.genblk1.pcpi_mul.rd[56] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[56] ),
    .Y(_04182_));
 sky130_fd_sc_hd__inv_2 _08845_ (.A(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__or2_1 _08846_ (.A(\genblk1.genblk1.pcpi_mul.rd[56] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[56] ),
    .X(_04184_));
 sky130_fd_sc_hd__a22o_1 _08847_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[57] ),
    .A2(net1103),
    .B1(_04182_),
    .B2(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__and4_1 _08848_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[57] ),
    .B(net1103),
    .C(_04182_),
    .D(_04184_),
    .X(_04186_));
 sky130_fd_sc_hd__inv_2 _08849_ (.A(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__a32o_1 _08850_ (.A1(net901),
    .A2(_04185_),
    .A3(_04187_),
    .B1(net2641),
    .B2(net1211),
    .X(_00140_));
 sky130_fd_sc_hd__a21o_1 _08851_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[58] ),
    .A2(net1105),
    .B1(\genblk1.genblk1.pcpi_mul.rd[57] ),
    .X(_04188_));
 sky130_fd_sc_hd__and3_1 _08852_ (.A(\genblk1.genblk1.pcpi_mul.rd[57] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[58] ),
    .C(net1105),
    .X(_04189_));
 sky130_fd_sc_hd__nand3_1 _08853_ (.A(\genblk1.genblk1.pcpi_mul.rd[57] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[58] ),
    .C(net1105),
    .Y(_04190_));
 sky130_fd_sc_hd__a211o_1 _08854_ (.A1(_04188_),
    .A2(_04190_),
    .B1(_04183_),
    .C1(_04186_),
    .X(_04191_));
 sky130_fd_sc_hd__o211a_1 _08855_ (.A1(_04183_),
    .A2(_04186_),
    .B1(_04188_),
    .C1(_04190_),
    .X(_04192_));
 sky130_fd_sc_hd__inv_2 _08856_ (.A(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__a32o_1 _08857_ (.A1(net901),
    .A2(_04191_),
    .A3(_04193_),
    .B1(net2878),
    .B2(net1213),
    .X(_00141_));
 sky130_fd_sc_hd__a21o_1 _08858_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[59] ),
    .A2(net1108),
    .B1(\genblk1.genblk1.pcpi_mul.rd[58] ),
    .X(_04194_));
 sky130_fd_sc_hd__nand3_1 _08859_ (.A(\genblk1.genblk1.pcpi_mul.rd[58] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[59] ),
    .C(net1108),
    .Y(_04195_));
 sky130_fd_sc_hd__a211o_1 _08860_ (.A1(_04194_),
    .A2(_04195_),
    .B1(_04189_),
    .C1(_04192_),
    .X(_04196_));
 sky130_fd_sc_hd__o211a_1 _08861_ (.A1(_04189_),
    .A2(_04192_),
    .B1(_04194_),
    .C1(_04195_),
    .X(_04197_));
 sky130_fd_sc_hd__inv_2 _08862_ (.A(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__a32o_1 _08863_ (.A1(net902),
    .A2(_04196_),
    .A3(_04198_),
    .B1(net2707),
    .B2(net1213),
    .X(_00142_));
 sky130_fd_sc_hd__nand3_1 _08864_ (.A(\genblk1.genblk1.pcpi_mul.rd[59] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[60] ),
    .C(net1108),
    .Y(_04199_));
 sky130_fd_sc_hd__a21o_1 _08865_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[60] ),
    .A2(net1105),
    .B1(\genblk1.genblk1.pcpi_mul.rd[59] ),
    .X(_04200_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_04199_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__nand2_1 _08867_ (.A(_04195_),
    .B(_04198_),
    .Y(_04202_));
 sky130_fd_sc_hd__xnor2_1 _08868_ (.A(_04201_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__a22o_1 _08869_ (.A1(net1213),
    .A2(net2917),
    .B1(net901),
    .B2(_04203_),
    .X(_00143_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(\genblk1.genblk1.pcpi_mul.rd[60] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[60] ),
    .Y(_04204_));
 sky130_fd_sc_hd__inv_2 _08871_ (.A(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__or2_1 _08872_ (.A(\genblk1.genblk1.pcpi_mul.rd[60] ),
    .B(\genblk1.genblk1.pcpi_mul.rdx[60] ),
    .X(_04206_));
 sky130_fd_sc_hd__a22o_1 _08873_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[61] ),
    .A2(net1106),
    .B1(_04204_),
    .B2(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__and4_1 _08874_ (.A(\genblk1.genblk1.pcpi_mul.next_rs2[61] ),
    .B(net1106),
    .C(_04204_),
    .D(_04206_),
    .X(_04208_));
 sky130_fd_sc_hd__nand2_1 _08875_ (.A(net904),
    .B(_04207_),
    .Y(_04209_));
 sky130_fd_sc_hd__a2bb2o_1 _08876_ (.A1_N(_04209_),
    .A2_N(_04208_),
    .B1(net2815),
    .B2(net1217),
    .X(_00144_));
 sky130_fd_sc_hd__a21o_1 _08877_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[62] ),
    .A2(net1106),
    .B1(\genblk1.genblk1.pcpi_mul.rd[61] ),
    .X(_04210_));
 sky130_fd_sc_hd__nand3_1 _08878_ (.A(\genblk1.genblk1.pcpi_mul.rd[61] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[62] ),
    .C(net1107),
    .Y(_04211_));
 sky130_fd_sc_hd__a211o_1 _08879_ (.A1(_04210_),
    .A2(_04211_),
    .B1(_04205_),
    .C1(_04208_),
    .X(_04212_));
 sky130_fd_sc_hd__o211a_1 _08880_ (.A1(_04205_),
    .A2(_04208_),
    .B1(_04210_),
    .C1(_04211_),
    .X(_04213_));
 sky130_fd_sc_hd__inv_2 _08881_ (.A(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__a32o_1 _08882_ (.A1(net904),
    .A2(_04212_),
    .A3(_04214_),
    .B1(net2721),
    .B2(net1217),
    .X(_00145_));
 sky130_fd_sc_hd__a21o_1 _08883_ (.A1(\genblk1.genblk1.pcpi_mul.next_rs2[63] ),
    .A2(net1107),
    .B1(\genblk1.genblk1.pcpi_mul.rd[62] ),
    .X(_04215_));
 sky130_fd_sc_hd__nand3_1 _08884_ (.A(\genblk1.genblk1.pcpi_mul.rd[62] ),
    .B(\genblk1.genblk1.pcpi_mul.next_rs2[63] ),
    .C(net1107),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_1 _08885_ (.A(_04215_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(_04211_),
    .B(_04214_),
    .Y(_04218_));
 sky130_fd_sc_hd__xnor2_1 _08887_ (.A(_04217_),
    .B(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__a22o_1 _08888_ (.A1(net1217),
    .A2(net2949),
    .B1(net904),
    .B2(_04219_),
    .X(_00146_));
 sky130_fd_sc_hd__a21bo_1 _08889_ (.A1(_04215_),
    .A2(_04218_),
    .B1_N(_04216_),
    .X(_04220_));
 sky130_fd_sc_hd__nand2_1 _08890_ (.A(net1107),
    .B(\genblk1.genblk1.pcpi_mul.rs2[63] ),
    .Y(_04221_));
 sky130_fd_sc_hd__xor2_1 _08891_ (.A(\genblk1.genblk1.pcpi_mul.rd[63] ),
    .B(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__xnor2_1 _08892_ (.A(_04220_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__a22o_1 _08893_ (.A1(net1217),
    .A2(net2941),
    .B1(net904),
    .B2(_04223_),
    .X(_00147_));
 sky130_fd_sc_hd__a21bo_1 _08894_ (.A1(_03892_),
    .A2(_03894_),
    .B1_N(_03891_),
    .X(_04224_));
 sky130_fd_sc_hd__a22o_1 _08895_ (.A1(net1200),
    .A2(net2674),
    .B1(net893),
    .B2(_04224_),
    .X(_00148_));
 sky130_fd_sc_hd__a21bo_1 _08896_ (.A1(_03914_),
    .A2(_03916_),
    .B1_N(_03913_),
    .X(_04225_));
 sky130_fd_sc_hd__a22o_1 _08897_ (.A1(net1195),
    .A2(net2646),
    .B1(net888),
    .B2(_04225_),
    .X(_00149_));
 sky130_fd_sc_hd__a21bo_1 _08898_ (.A1(_03936_),
    .A2(_03938_),
    .B1_N(_03935_),
    .X(_04226_));
 sky130_fd_sc_hd__a22o_1 _08899_ (.A1(net1192),
    .A2(net2649),
    .B1(net885),
    .B2(_04226_),
    .X(_00150_));
 sky130_fd_sc_hd__a21bo_1 _08900_ (.A1(_03958_),
    .A2(_03960_),
    .B1_N(_03957_),
    .X(_04227_));
 sky130_fd_sc_hd__a22o_1 _08901_ (.A1(net1196),
    .A2(net2712),
    .B1(net890),
    .B2(_04227_),
    .X(_00151_));
 sky130_fd_sc_hd__a21bo_1 _08902_ (.A1(_03980_),
    .A2(_03982_),
    .B1_N(_03979_),
    .X(_04228_));
 sky130_fd_sc_hd__a22o_1 _08903_ (.A1(net1202),
    .A2(net2621),
    .B1(net896),
    .B2(_04228_),
    .X(_00152_));
 sky130_fd_sc_hd__a21bo_1 _08904_ (.A1(_04002_),
    .A2(_04004_),
    .B1_N(_04001_),
    .X(_04229_));
 sky130_fd_sc_hd__a22o_1 _08905_ (.A1(net1210),
    .A2(net2706),
    .B1(net899),
    .B2(_04229_),
    .X(_00153_));
 sky130_fd_sc_hd__a21bo_1 _08906_ (.A1(_04024_),
    .A2(_04026_),
    .B1_N(_04023_),
    .X(_04230_));
 sky130_fd_sc_hd__a22o_1 _08907_ (.A1(net1212),
    .A2(net2625),
    .B1(net904),
    .B2(_04230_),
    .X(_00154_));
 sky130_fd_sc_hd__a21bo_1 _08908_ (.A1(_04046_),
    .A2(_04048_),
    .B1_N(_04045_),
    .X(_04231_));
 sky130_fd_sc_hd__a22o_1 _08909_ (.A1(net1210),
    .A2(net2780),
    .B1(net899),
    .B2(_04231_),
    .X(_00155_));
 sky130_fd_sc_hd__a21bo_1 _08910_ (.A1(_04068_),
    .A2(_04070_),
    .B1_N(_04067_),
    .X(_04232_));
 sky130_fd_sc_hd__a22o_1 _08911_ (.A1(net1200),
    .A2(net2662),
    .B1(net893),
    .B2(_04232_),
    .X(_00156_));
 sky130_fd_sc_hd__a21bo_1 _08912_ (.A1(_04090_),
    .A2(_04092_),
    .B1_N(_04089_),
    .X(_04233_));
 sky130_fd_sc_hd__a22o_1 _08913_ (.A1(net1195),
    .A2(net2711),
    .B1(net888),
    .B2(_04233_),
    .X(_00157_));
 sky130_fd_sc_hd__a21bo_1 _08914_ (.A1(_04112_),
    .A2(_04114_),
    .B1_N(_04111_),
    .X(_04234_));
 sky130_fd_sc_hd__a22o_1 _08915_ (.A1(net1194),
    .A2(net2679),
    .B1(net886),
    .B2(_04234_),
    .X(_00158_));
 sky130_fd_sc_hd__a21bo_1 _08916_ (.A1(_04134_),
    .A2(_04136_),
    .B1_N(_04133_),
    .X(_04235_));
 sky130_fd_sc_hd__a22o_1 _08917_ (.A1(net1196),
    .A2(net2640),
    .B1(net888),
    .B2(_04235_),
    .X(_00159_));
 sky130_fd_sc_hd__a21bo_1 _08918_ (.A1(_04156_),
    .A2(_04158_),
    .B1_N(_04155_),
    .X(_04236_));
 sky130_fd_sc_hd__a22o_1 _08919_ (.A1(net1203),
    .A2(net2708),
    .B1(net895),
    .B2(_04236_),
    .X(_00160_));
 sky130_fd_sc_hd__a21bo_1 _08920_ (.A1(_04178_),
    .A2(_04180_),
    .B1_N(_04177_),
    .X(_04237_));
 sky130_fd_sc_hd__a22o_1 _08921_ (.A1(net1211),
    .A2(net2670),
    .B1(net900),
    .B2(_04237_),
    .X(_00161_));
 sky130_fd_sc_hd__a21bo_1 _08922_ (.A1(_04200_),
    .A2(_04202_),
    .B1_N(_04199_),
    .X(_04238_));
 sky130_fd_sc_hd__a22o_1 _08923_ (.A1(net1213),
    .A2(net2665),
    .B1(net901),
    .B2(_04238_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _08924_ (.A0(\genblk1.genblk1.pcpi_mul.rd[0] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[32] ),
    .S(net956),
    .X(_04239_));
 sky130_fd_sc_hd__mux2_1 _08925_ (.A0(net1393),
    .A1(_04239_),
    .S(net945),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _08926_ (.A0(\genblk1.genblk1.pcpi_mul.rd[1] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[33] ),
    .S(net957),
    .X(_04240_));
 sky130_fd_sc_hd__mux2_1 _08927_ (.A0(net1467),
    .A1(_04240_),
    .S(net945),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _08928_ (.A0(\genblk1.genblk1.pcpi_mul.rd[2] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[34] ),
    .S(net955),
    .X(_04241_));
 sky130_fd_sc_hd__mux2_1 _08929_ (.A0(net1436),
    .A1(_04241_),
    .S(net944),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _08930_ (.A0(\genblk1.genblk1.pcpi_mul.rd[3] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[35] ),
    .S(net955),
    .X(_04242_));
 sky130_fd_sc_hd__mux2_1 _08931_ (.A0(net1633),
    .A1(_04242_),
    .S(net944),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _08932_ (.A0(\genblk1.genblk1.pcpi_mul.rd[4] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[36] ),
    .S(net955),
    .X(_04243_));
 sky130_fd_sc_hd__mux2_1 _08933_ (.A0(net2635),
    .A1(_04243_),
    .S(net944),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _08934_ (.A0(\genblk1.genblk1.pcpi_mul.rd[5] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[37] ),
    .S(net955),
    .X(_04244_));
 sky130_fd_sc_hd__mux2_1 _08935_ (.A0(net2539),
    .A1(_04244_),
    .S(net944),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _08936_ (.A0(\genblk1.genblk1.pcpi_mul.rd[6] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[38] ),
    .S(net955),
    .X(_04245_));
 sky130_fd_sc_hd__mux2_1 _08937_ (.A0(net2837),
    .A1(_04245_),
    .S(net944),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _08938_ (.A0(\genblk1.genblk1.pcpi_mul.rd[7] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[39] ),
    .S(net954),
    .X(_04246_));
 sky130_fd_sc_hd__mux2_1 _08939_ (.A0(net1861),
    .A1(_04246_),
    .S(net943),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _08940_ (.A0(\genblk1.genblk1.pcpi_mul.rd[8] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[40] ),
    .S(net954),
    .X(_04247_));
 sky130_fd_sc_hd__mux2_1 _08941_ (.A0(net1831),
    .A1(_04247_),
    .S(net943),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _08942_ (.A0(\genblk1.genblk1.pcpi_mul.rd[9] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[41] ),
    .S(net954),
    .X(_04248_));
 sky130_fd_sc_hd__mux2_1 _08943_ (.A0(net1374),
    .A1(_04248_),
    .S(net943),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _08944_ (.A0(\genblk1.genblk1.pcpi_mul.rd[10] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[42] ),
    .S(net954),
    .X(_04249_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(net2435),
    .A1(_04249_),
    .S(net943),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _08946_ (.A0(\genblk1.genblk1.pcpi_mul.rd[11] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[43] ),
    .S(net954),
    .X(_04250_));
 sky130_fd_sc_hd__mux2_1 _08947_ (.A0(net2739),
    .A1(_04250_),
    .S(net943),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _08948_ (.A0(\genblk1.genblk1.pcpi_mul.rd[12] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[44] ),
    .S(net954),
    .X(_04251_));
 sky130_fd_sc_hd__mux2_1 _08949_ (.A0(net2549),
    .A1(_04251_),
    .S(net943),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _08950_ (.A0(\genblk1.genblk1.pcpi_mul.rd[13] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[45] ),
    .S(net954),
    .X(_04252_));
 sky130_fd_sc_hd__mux2_1 _08951_ (.A0(net2430),
    .A1(_04252_),
    .S(net943),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _08952_ (.A0(\genblk1.genblk1.pcpi_mul.rd[14] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[46] ),
    .S(net954),
    .X(_04253_));
 sky130_fd_sc_hd__mux2_1 _08953_ (.A0(net2601),
    .A1(_04253_),
    .S(net943),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _08954_ (.A0(\genblk1.genblk1.pcpi_mul.rd[15] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[47] ),
    .S(net954),
    .X(_04254_));
 sky130_fd_sc_hd__mux2_1 _08955_ (.A0(net2568),
    .A1(_04254_),
    .S(net943),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _08956_ (.A0(\genblk1.genblk1.pcpi_mul.rd[16] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[48] ),
    .S(net954),
    .X(_04255_));
 sky130_fd_sc_hd__mux2_1 _08957_ (.A0(net2822),
    .A1(_04255_),
    .S(net943),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _08958_ (.A0(\genblk1.genblk1.pcpi_mul.rd[17] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[49] ),
    .S(net955),
    .X(_04256_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(net2091),
    .A1(_04256_),
    .S(net944),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _08960_ (.A0(\genblk1.genblk1.pcpi_mul.rd[18] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[50] ),
    .S(net955),
    .X(_04257_));
 sky130_fd_sc_hd__mux2_1 _08961_ (.A0(net2483),
    .A1(_04257_),
    .S(net944),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _08962_ (.A0(\genblk1.genblk1.pcpi_mul.rd[19] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[51] ),
    .S(net955),
    .X(_04258_));
 sky130_fd_sc_hd__mux2_1 _08963_ (.A0(net1676),
    .A1(_04258_),
    .S(net944),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _08964_ (.A0(\genblk1.genblk1.pcpi_mul.rd[20] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[52] ),
    .S(net955),
    .X(_04259_));
 sky130_fd_sc_hd__mux2_1 _08965_ (.A0(net2656),
    .A1(_04259_),
    .S(net945),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _08966_ (.A0(\genblk1.genblk1.pcpi_mul.rd[21] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[53] ),
    .S(net956),
    .X(_04260_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(net2300),
    .A1(_04260_),
    .S(net945),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _08968_ (.A0(\genblk1.genblk1.pcpi_mul.rd[22] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[54] ),
    .S(net956),
    .X(_04261_));
 sky130_fd_sc_hd__mux2_1 _08969_ (.A0(net1731),
    .A1(_04261_),
    .S(net945),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _08970_ (.A0(\genblk1.genblk1.pcpi_mul.rd[23] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[55] ),
    .S(net956),
    .X(_04262_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(net1460),
    .A1(_04262_),
    .S(net945),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _08972_ (.A0(\genblk1.genblk1.pcpi_mul.rd[24] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[56] ),
    .S(net956),
    .X(_04263_));
 sky130_fd_sc_hd__mux2_1 _08973_ (.A0(net1389),
    .A1(_04263_),
    .S(net945),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _08974_ (.A0(\genblk1.genblk1.pcpi_mul.rd[25] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[57] ),
    .S(net956),
    .X(_04264_));
 sky130_fd_sc_hd__mux2_1 _08975_ (.A0(net1424),
    .A1(_04264_),
    .S(net946),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _08976_ (.A0(\genblk1.genblk1.pcpi_mul.rd[26] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[58] ),
    .S(net957),
    .X(_04265_));
 sky130_fd_sc_hd__mux2_1 _08977_ (.A0(net1629),
    .A1(_04265_),
    .S(net945),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _08978_ (.A0(\genblk1.genblk1.pcpi_mul.rd[27] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[59] ),
    .S(net956),
    .X(_04266_));
 sky130_fd_sc_hd__mux2_1 _08979_ (.A0(net1382),
    .A1(_04266_),
    .S(net946),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _08980_ (.A0(\genblk1.genblk1.pcpi_mul.rd[28] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[60] ),
    .S(net957),
    .X(_04267_));
 sky130_fd_sc_hd__mux2_1 _08981_ (.A0(net1626),
    .A1(_04267_),
    .S(net946),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _08982_ (.A0(\genblk1.genblk1.pcpi_mul.rd[29] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[61] ),
    .S(net956),
    .X(_04268_));
 sky130_fd_sc_hd__mux2_1 _08983_ (.A0(net1504),
    .A1(_04268_),
    .S(net946),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _08984_ (.A0(\genblk1.genblk1.pcpi_mul.rd[30] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[62] ),
    .S(net957),
    .X(_04269_));
 sky130_fd_sc_hd__mux2_1 _08985_ (.A0(net1496),
    .A1(_04269_),
    .S(net946),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _08986_ (.A0(\genblk1.genblk1.pcpi_mul.rd[31] ),
    .A1(\genblk1.genblk1.pcpi_mul.rd[63] ),
    .S(net957),
    .X(_04270_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(net1748),
    .A1(_04270_),
    .S(net945),
    .X(_00194_));
 sky130_fd_sc_hd__and3b_1 _08988_ (.A_N(\genblk1.genblk1.pcpi_mul.pcpi_wait_q ),
    .B(net917),
    .C(net1315),
    .X(_04271_));
 sky130_fd_sc_hd__a21oi_1 _08989_ (.A1(_02414_),
    .A2(net907),
    .B1(_04271_),
    .Y(_00195_));
 sky130_fd_sc_hd__or3b_1 _08990_ (.A(\latched_rd[2] ),
    .B(\latched_rd[4] ),
    .C_N(\latched_rd[3] ),
    .X(_04272_));
 sky130_fd_sc_hd__or3_4 _08991_ (.A(\latched_rd[1] ),
    .B(\latched_rd[0] ),
    .C(_03743_),
    .X(_04273_));
 sky130_fd_sc_hd__or2_1 _08992_ (.A(_04272_),
    .B(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__mux2_1 _08993_ (.A0(net588),
    .A1(net1974),
    .S(net518),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _08994_ (.A0(net584),
    .A1(net1905),
    .S(net518),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _08995_ (.A0(net580),
    .A1(net1699),
    .S(net518),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _08996_ (.A0(net575),
    .A1(net1730),
    .S(net517),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _08997_ (.A0(net572),
    .A1(net1927),
    .S(net518),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _08998_ (.A0(net541),
    .A1(net2067),
    .S(net517),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _08999_ (.A0(net537),
    .A1(net1964),
    .S(net516),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _09000_ (.A0(net526),
    .A1(net1957),
    .S(net516),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _09001_ (.A0(net521),
    .A1(net1685),
    .S(net516),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _09002_ (.A0(net408),
    .A1(net2081),
    .S(net516),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _09003_ (.A0(net403),
    .A1(net1767),
    .S(net517),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _09004_ (.A0(net356),
    .A1(net1760),
    .S(net516),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _09005_ (.A0(net352),
    .A1(net1802),
    .S(net516),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _09006_ (.A0(net349),
    .A1(net1488),
    .S(net516),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _09007_ (.A0(net346),
    .A1(net1705),
    .S(net517),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _09008_ (.A0(net342),
    .A1(net2056),
    .S(net516),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _09009_ (.A0(net337),
    .A1(net2009),
    .S(net517),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _09010_ (.A0(net334),
    .A1(net1741),
    .S(net516),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _09011_ (.A0(net329),
    .A1(net1531),
    .S(net516),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _09012_ (.A0(net326),
    .A1(net2275),
    .S(net518),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _09013_ (.A0(net322),
    .A1(net2120),
    .S(net517),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _09014_ (.A0(net318),
    .A1(net1665),
    .S(net517),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _09015_ (.A0(net313),
    .A1(net2041),
    .S(net518),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _09016_ (.A0(net308),
    .A1(net1969),
    .S(net517),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _09017_ (.A0(net305),
    .A1(net1901),
    .S(net518),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _09018_ (.A0(net304),
    .A1(net2195),
    .S(net519),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _09019_ (.A0(net299),
    .A1(net2078),
    .S(net518),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _09020_ (.A0(net296),
    .A1(net2090),
    .S(net518),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _09021_ (.A0(net289),
    .A1(net1662),
    .S(net519),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _09022_ (.A0(net287),
    .A1(net1838),
    .S(net519),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _09023_ (.A0(net282),
    .A1(net2076),
    .S(net518),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _09024_ (.A0(net281),
    .A1(net2084),
    .S(net519),
    .X(_00227_));
 sky130_fd_sc_hd__or3b_4 _09025_ (.A(_03743_),
    .B(\latched_rd[1] ),
    .C_N(\latched_rd[0] ),
    .X(_04275_));
 sky130_fd_sc_hd__or2_1 _09026_ (.A(_03744_),
    .B(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__mux2_1 _09027_ (.A0(_03749_),
    .A1(net2326),
    .S(net514),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _09028_ (.A0(net585),
    .A1(net2327),
    .S(net514),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _09029_ (.A0(net580),
    .A1(net2524),
    .S(net514),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _09030_ (.A0(net576),
    .A1(net2485),
    .S(net513),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _09031_ (.A0(net571),
    .A1(net2254),
    .S(net513),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _09032_ (.A0(net541),
    .A1(net2482),
    .S(net513),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _09033_ (.A0(net537),
    .A1(net2297),
    .S(net512),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _09034_ (.A0(net527),
    .A1(net2221),
    .S(net512),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _09035_ (.A0(net521),
    .A1(net2143),
    .S(net513),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _09036_ (.A0(net408),
    .A1(net2513),
    .S(net513),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _09037_ (.A0(net403),
    .A1(net2266),
    .S(net513),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _09038_ (.A0(net356),
    .A1(net2312),
    .S(net512),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _09039_ (.A0(net353),
    .A1(net2298),
    .S(net512),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _09040_ (.A0(net349),
    .A1(net2351),
    .S(net512),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(net346),
    .A1(net2445),
    .S(net512),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _09042_ (.A0(net342),
    .A1(net2403),
    .S(net512),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _09043_ (.A0(net338),
    .A1(net2229),
    .S(net512),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _09044_ (.A0(net334),
    .A1(net2267),
    .S(net512),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(net330),
    .A1(net2426),
    .S(net512),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _09046_ (.A0(net326),
    .A1(net2411),
    .S(net515),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(net322),
    .A1(net2137),
    .S(net513),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _09048_ (.A0(net317),
    .A1(net2346),
    .S(net513),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _09049_ (.A0(net314),
    .A1(net2329),
    .S(net514),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _09050_ (.A0(net309),
    .A1(net2422),
    .S(net513),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _09051_ (.A0(net306),
    .A1(net2095),
    .S(net514),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _09052_ (.A0(net301),
    .A1(net2167),
    .S(net514),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _09053_ (.A0(net297),
    .A1(net2457),
    .S(net514),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _09054_ (.A0(net293),
    .A1(net2418),
    .S(net514),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _09055_ (.A0(net291),
    .A1(net2413),
    .S(net514),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _09056_ (.A0(net286),
    .A1(net2348),
    .S(net514),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _09057_ (.A0(net284),
    .A1(net2514),
    .S(net515),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _09058_ (.A0(net278),
    .A1(net2419),
    .S(net515),
    .X(_00259_));
 sky130_fd_sc_hd__nand3b_4 _09059_ (.A_N(\latched_rd[3] ),
    .B(\latched_rd[4] ),
    .C(\latched_rd[2] ),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_4 _09060_ (.A(_04273_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__mux2_1 _09061_ (.A0(net1572),
    .A1(net587),
    .S(net510),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _09062_ (.A0(net1950),
    .A1(net583),
    .S(net510),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _09063_ (.A0(net1404),
    .A1(net581),
    .S(net511),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _09064_ (.A0(net1434),
    .A1(net577),
    .S(net508),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _09065_ (.A0(net1386),
    .A1(net573),
    .S(net511),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _09066_ (.A0(net1361),
    .A1(net543),
    .S(net511),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _09067_ (.A0(net2129),
    .A1(net539),
    .S(net508),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _09068_ (.A0(net1507),
    .A1(net524),
    .S(net508),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _09069_ (.A0(net1607),
    .A1(net523),
    .S(net509),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _09070_ (.A0(net1930),
    .A1(net407),
    .S(net509),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _09071_ (.A0(net1534),
    .A1(net405),
    .S(net509),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _09072_ (.A0(net1728),
    .A1(net354),
    .S(net509),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _09073_ (.A0(net1552),
    .A1(net350),
    .S(net508),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _09074_ (.A0(net1745),
    .A1(net347),
    .S(net508),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _09075_ (.A0(net1850),
    .A1(net343),
    .S(net509),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _09076_ (.A0(net1599),
    .A1(net339),
    .S(net508),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _09077_ (.A0(net1852),
    .A1(net336),
    .S(net508),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _09078_ (.A0(net1514),
    .A1(net332),
    .S(net508),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _09079_ (.A0(net1471),
    .A1(net328),
    .S(net508),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _09080_ (.A0(net2103),
    .A1(net324),
    .S(net510),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _09081_ (.A0(net1598),
    .A1(net320),
    .S(net508),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _09082_ (.A0(net1704),
    .A1(net316),
    .S(net510),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _09083_ (.A0(net1395),
    .A1(net312),
    .S(net510),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _09084_ (.A0(net1538),
    .A1(net311),
    .S(net510),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _09085_ (.A0(net1666),
    .A1(net305),
    .S(net511),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(net1416),
    .A1(net302),
    .S(net511),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _09087_ (.A0(net1719),
    .A1(net298),
    .S(net511),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _09088_ (.A0(net1456),
    .A1(net294),
    .S(net510),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(net1608),
    .A1(net289),
    .S(net510),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _09090_ (.A0(net1545),
    .A1(net285),
    .S(net511),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _09091_ (.A0(net1498),
    .A1(net283),
    .S(net510),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _09092_ (.A0(net1995),
    .A1(net278),
    .S(net510),
    .X(_00291_));
 sky130_fd_sc_hd__nor2_4 _09093_ (.A(_04275_),
    .B(_04277_),
    .Y(_04279_));
 sky130_fd_sc_hd__mux2_1 _09094_ (.A0(net2250),
    .A1(net587),
    .S(net506),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _09095_ (.A0(net2538),
    .A1(net583),
    .S(net506),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _09096_ (.A0(net2047),
    .A1(net581),
    .S(net507),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _09097_ (.A0(net1889),
    .A1(net577),
    .S(net504),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _09098_ (.A0(net1918),
    .A1(net574),
    .S(net507),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _09099_ (.A0(net1650),
    .A1(net543),
    .S(net507),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _09100_ (.A0(net1792),
    .A1(net539),
    .S(net504),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _09101_ (.A0(net1501),
    .A1(net524),
    .S(net504),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _09102_ (.A0(net1668),
    .A1(net523),
    .S(net505),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _09103_ (.A0(net1773),
    .A1(net407),
    .S(net505),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _09104_ (.A0(net1568),
    .A1(net405),
    .S(net505),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _09105_ (.A0(net1840),
    .A1(net354),
    .S(net505),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _09106_ (.A0(net1744),
    .A1(net350),
    .S(net504),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _09107_ (.A0(net1887),
    .A1(net347),
    .S(net504),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _09108_ (.A0(net1933),
    .A1(net343),
    .S(net505),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _09109_ (.A0(net1475),
    .A1(net339),
    .S(net504),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _09110_ (.A0(net1912),
    .A1(net336),
    .S(net504),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _09111_ (.A0(net1725),
    .A1(net332),
    .S(net504),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _09112_ (.A0(net1835),
    .A1(net328),
    .S(net504),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _09113_ (.A0(net2291),
    .A1(net324),
    .S(net506),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _09114_ (.A0(net1502),
    .A1(net320),
    .S(net504),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _09115_ (.A0(net1653),
    .A1(net316),
    .S(net506),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(net1882),
    .A1(net312),
    .S(net506),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _09117_ (.A0(net2094),
    .A1(net310),
    .S(net506),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _09118_ (.A0(net1702),
    .A1(net305),
    .S(net507),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _09119_ (.A0(net1801),
    .A1(net302),
    .S(net507),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(net2219),
    .A1(net298),
    .S(net507),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _09121_ (.A0(net1959),
    .A1(net294),
    .S(net506),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(net2373),
    .A1(net289),
    .S(net506),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _09123_ (.A0(net1992),
    .A1(net285),
    .S(net507),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(net2244),
    .A1(net283),
    .S(net506),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _09125_ (.A0(net1865),
    .A1(net278),
    .S(net506),
    .X(_00323_));
 sky130_fd_sc_hd__nand2_1 _09126_ (.A(\latched_rd[4] ),
    .B(\latched_rd[3] ),
    .Y(_04280_));
 sky130_fd_sc_hd__nand3_2 _09127_ (.A(\latched_rd[2] ),
    .B(\latched_rd[4] ),
    .C(\latched_rd[3] ),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(\latched_rd[1] ),
    .B(\latched_rd[0] ),
    .Y(_04282_));
 sky130_fd_sc_hd__or2_2 _09129_ (.A(_03743_),
    .B(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__nor2_1 _09130_ (.A(_04281_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__mux2_1 _09131_ (.A0(net2071),
    .A1(net586),
    .S(net502),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _09132_ (.A0(net2225),
    .A1(net585),
    .S(net502),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _09133_ (.A0(net1474),
    .A1(net581),
    .S(net502),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(net1620),
    .A1(net578),
    .S(net501),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _09135_ (.A0(net1825),
    .A1(net573),
    .S(net501),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(net1750),
    .A1(net542),
    .S(net501),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _09137_ (.A0(net1616),
    .A1(net539),
    .S(net500),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _09138_ (.A0(net1603),
    .A1(net524),
    .S(net500),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _09139_ (.A0(net1600),
    .A1(net523),
    .S(net500),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _09140_ (.A0(net1867),
    .A1(net409),
    .S(net500),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _09141_ (.A0(net1564),
    .A1(net406),
    .S(net501),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _09142_ (.A0(net1652),
    .A1(net354),
    .S(net501),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _09143_ (.A0(net1683),
    .A1(net351),
    .S(net500),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _09144_ (.A0(net1422),
    .A1(net347),
    .S(net500),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _09145_ (.A0(net1758),
    .A1(net343),
    .S(net500),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _09146_ (.A0(net1656),
    .A1(net340),
    .S(net500),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _09147_ (.A0(net1764),
    .A1(net338),
    .S(net501),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _09148_ (.A0(net1763),
    .A1(net333),
    .S(net500),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _09149_ (.A0(net1687),
    .A1(net330),
    .S(net500),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _09150_ (.A0(net2073),
    .A1(net327),
    .S(net502),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _09151_ (.A0(net1875),
    .A1(net323),
    .S(net501),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _09152_ (.A0(net1509),
    .A1(net318),
    .S(net501),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _09153_ (.A0(net2020),
    .A1(net314),
    .S(net502),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(net1618),
    .A1(net310),
    .S(net502),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _09155_ (.A0(net1523),
    .A1(net307),
    .S(net502),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(net1935),
    .A1(net303),
    .S(net503),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(net2093),
    .A1(net299),
    .S(net503),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(net2098),
    .A1(net295),
    .S(net503),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(net1908),
    .A1(net291),
    .S(net502),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(net2124),
    .A1(net287),
    .S(net502),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(net1934),
    .A1(net284),
    .S(net502),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(net2061),
    .A1(net280),
    .S(net503),
    .X(_00355_));
 sky130_fd_sc_hd__or2_1 _09163_ (.A(_03744_),
    .B(_03745_),
    .X(_04285_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(net588),
    .A1(net1900),
    .S(net498),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _09165_ (.A0(net585),
    .A1(net2320),
    .S(net498),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(net580),
    .A1(net1774),
    .S(net499),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(net576),
    .A1(net2050),
    .S(net496),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(net571),
    .A1(net2341),
    .S(net496),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(net541),
    .A1(net2224),
    .S(net499),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(net537),
    .A1(net2208),
    .S(net496),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _09171_ (.A0(net526),
    .A1(net2387),
    .S(net496),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(net521),
    .A1(net1819),
    .S(net496),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _09173_ (.A0(net408),
    .A1(net1921),
    .S(net496),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(net403),
    .A1(net2021),
    .S(net496),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _09175_ (.A0(net356),
    .A1(net2140),
    .S(net496),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(net353),
    .A1(net2187),
    .S(net497),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _09177_ (.A0(net349),
    .A1(net1976),
    .S(net497),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(net346),
    .A1(net2385),
    .S(net496),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _09179_ (.A0(net342),
    .A1(net2037),
    .S(net497),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(_03810_),
    .A1(net1808),
    .S(net497),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _09181_ (.A0(net335),
    .A1(net2151),
    .S(net497),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(net330),
    .A1(net1729),
    .S(net497),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _09183_ (.A0(net326),
    .A1(net1783),
    .S(net497),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(net322),
    .A1(net2014),
    .S(net497),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _09185_ (.A0(net317),
    .A1(net2112),
    .S(net497),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(net315),
    .A1(net1987),
    .S(net498),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(net309),
    .A1(net2241),
    .S(net496),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _09188_ (.A0(net307),
    .A1(net1570),
    .S(net498),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _09189_ (.A0(net301),
    .A1(net1765),
    .S(net498),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(net297),
    .A1(net1945),
    .S(net498),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _09191_ (.A0(net293),
    .A1(net2051),
    .S(net498),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(net291),
    .A1(net1949),
    .S(net498),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _09193_ (.A0(net286),
    .A1(net2125),
    .S(net499),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(net284),
    .A1(net2054),
    .S(net498),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _09195_ (.A0(net278),
    .A1(net2285),
    .S(net498),
    .X(_00387_));
 sky130_fd_sc_hd__nor2_2 _09196_ (.A(_04275_),
    .B(_04281_),
    .Y(_04286_));
 sky130_fd_sc_hd__mux2_1 _09197_ (.A0(net1539),
    .A1(net586),
    .S(net494),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(net2199),
    .A1(net585),
    .S(net494),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(net2007),
    .A1(net582),
    .S(net494),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(net1609),
    .A1(net577),
    .S(net493),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(net1916),
    .A1(net573),
    .S(net494),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(net1536),
    .A1(net542),
    .S(net493),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(net1587),
    .A1(net539),
    .S(net492),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(net1897),
    .A1(net525),
    .S(net492),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(net1851),
    .A1(net522),
    .S(net492),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(net1766),
    .A1(net409),
    .S(net492),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(net1430),
    .A1(net405),
    .S(net493),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(net1648),
    .A1(net354),
    .S(net493),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(net1427),
    .A1(net350),
    .S(net492),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(net1453),
    .A1(net347),
    .S(net492),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(net1841),
    .A1(net343),
    .S(net492),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(net1697),
    .A1(net340),
    .S(net492),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _09213_ (.A0(net1734),
    .A1(net338),
    .S(net493),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(net1714),
    .A1(net333),
    .S(net492),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(net1713),
    .A1(net330),
    .S(net492),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _09216_ (.A0(net2190),
    .A1(net326),
    .S(net494),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _09217_ (.A0(net1606),
    .A1(net322),
    .S(net493),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _09218_ (.A0(net1511),
    .A1(net319),
    .S(net493),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _09219_ (.A0(net1592),
    .A1(net314),
    .S(net494),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _09220_ (.A0(net1993),
    .A1(net310),
    .S(net494),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(net1997),
    .A1(net307),
    .S(net494),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _09222_ (.A0(net1820),
    .A1(net303),
    .S(net495),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _09223_ (.A0(net1932),
    .A1(net299),
    .S(net495),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _09224_ (.A0(net1654),
    .A1(net295),
    .S(net494),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _09225_ (.A0(net1772),
    .A1(net292),
    .S(net494),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _09226_ (.A0(net1829),
    .A1(net287),
    .S(net495),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _09227_ (.A0(net1674),
    .A1(net284),
    .S(net495),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _09228_ (.A0(net1751),
    .A1(net280),
    .S(net495),
    .X(_00419_));
 sky130_fd_sc_hd__nor2_4 _09229_ (.A(_03745_),
    .B(_04277_),
    .Y(_04287_));
 sky130_fd_sc_hd__mux2_1 _09230_ (.A0(net1555),
    .A1(net587),
    .S(net490),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _09231_ (.A0(net1490),
    .A1(net583),
    .S(net490),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _09232_ (.A0(net1360),
    .A1(net581),
    .S(net491),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _09233_ (.A0(net1845),
    .A1(net577),
    .S(net489),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _09234_ (.A0(net1658),
    .A1(net574),
    .S(net491),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _09235_ (.A0(net1715),
    .A1(net543),
    .S(net491),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _09236_ (.A0(net1637),
    .A1(net539),
    .S(net488),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _09237_ (.A0(net1958),
    .A1(net524),
    .S(net488),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _09238_ (.A0(net1529),
    .A1(net520),
    .S(net488),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _09239_ (.A0(net1469),
    .A1(net408),
    .S(net489),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(net1749),
    .A1(net405),
    .S(net489),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _09241_ (.A0(net1548),
    .A1(net354),
    .S(net489),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _09242_ (.A0(net1689),
    .A1(net350),
    .S(net488),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _09243_ (.A0(net1892),
    .A1(net347),
    .S(net488),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _09244_ (.A0(net1392),
    .A1(net343),
    .S(net489),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _09245_ (.A0(net1667),
    .A1(net339),
    .S(net488),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _09246_ (.A0(net1528),
    .A1(net336),
    .S(net488),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _09247_ (.A0(net1701),
    .A1(net332),
    .S(net488),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _09248_ (.A0(net1810),
    .A1(net328),
    .S(net488),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(net1440),
    .A1(net324),
    .S(net490),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _09250_ (.A0(net1385),
    .A1(net320),
    .S(net488),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _09251_ (.A0(net1591),
    .A1(net316),
    .S(net490),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _09252_ (.A0(net1481),
    .A1(net312),
    .S(net490),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _09253_ (.A0(net1602),
    .A1(net308),
    .S(net490),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _09254_ (.A0(net1660),
    .A1(_03844_),
    .S(net491),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(net1619),
    .A1(net302),
    .S(net491),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _09256_ (.A0(net1421),
    .A1(net298),
    .S(net491),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(net1679),
    .A1(net294),
    .S(net490),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _09258_ (.A0(net1780),
    .A1(net289),
    .S(net490),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(net1513),
    .A1(net285),
    .S(net491),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _09260_ (.A0(net2002),
    .A1(net283),
    .S(net490),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _09261_ (.A0(net1768),
    .A1(net278),
    .S(net490),
    .X(_00451_));
 sky130_fd_sc_hd__nor2_4 _09262_ (.A(_04277_),
    .B(_04283_),
    .Y(_04288_));
 sky130_fd_sc_hd__mux2_1 _09263_ (.A0(net2191),
    .A1(net587),
    .S(net486),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _09264_ (.A0(net2322),
    .A1(net583),
    .S(net486),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _09265_ (.A0(net1830),
    .A1(net581),
    .S(net487),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _09266_ (.A0(net1651),
    .A1(net577),
    .S(net485),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _09267_ (.A0(net1517),
    .A1(net574),
    .S(net487),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _09268_ (.A0(net2087),
    .A1(net543),
    .S(net487),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(net1643),
    .A1(net539),
    .S(net484),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _09270_ (.A0(net1948),
    .A1(net524),
    .S(net484),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _09271_ (.A0(net2012),
    .A1(net520),
    .S(net484),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _09272_ (.A0(net1703),
    .A1(net408),
    .S(net485),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _09273_ (.A0(net1804),
    .A1(net405),
    .S(net485),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _09274_ (.A0(net1880),
    .A1(net354),
    .S(net485),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _09275_ (.A0(net1691),
    .A1(net350),
    .S(net484),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _09276_ (.A0(net1611),
    .A1(net347),
    .S(net484),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _09277_ (.A0(net1577),
    .A1(net343),
    .S(net485),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _09278_ (.A0(net1454),
    .A1(net339),
    .S(net484),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _09279_ (.A0(net1525),
    .A1(net336),
    .S(net484),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _09280_ (.A0(net1869),
    .A1(net332),
    .S(net484),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _09281_ (.A0(net1573),
    .A1(net328),
    .S(net484),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _09282_ (.A0(net1822),
    .A1(net324),
    .S(net486),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _09283_ (.A0(net2201),
    .A1(net320),
    .S(net484),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _09284_ (.A0(net1500),
    .A1(net316),
    .S(net486),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _09285_ (.A0(net2177),
    .A1(net312),
    .S(net486),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _09286_ (.A0(net1612),
    .A1(net308),
    .S(net486),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _09287_ (.A0(net1970),
    .A1(_03844_),
    .S(net487),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _09288_ (.A0(net1721),
    .A1(net302),
    .S(net487),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(net2082),
    .A1(net298),
    .S(net487),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _09290_ (.A0(net1818),
    .A1(net294),
    .S(net486),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _09291_ (.A0(net2355),
    .A1(net289),
    .S(net486),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _09292_ (.A0(net1799),
    .A1(net285),
    .S(net487),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _09293_ (.A0(net2499),
    .A1(net283),
    .S(net486),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(net2077),
    .A1(net278),
    .S(net486),
    .X(_00483_));
 sky130_fd_sc_hd__or3_1 _09295_ (.A(\latched_rd[2] ),
    .B(_03743_),
    .C(_04280_),
    .X(_04289_));
 sky130_fd_sc_hd__inv_2 _09296_ (.A(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__nor3_2 _09297_ (.A(\latched_rd[1] ),
    .B(\latched_rd[0] ),
    .C(_04289_),
    .Y(_04291_));
 sky130_fd_sc_hd__mux2_1 _09298_ (.A0(net1894),
    .A1(net586),
    .S(net481),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(net1746),
    .A1(net584),
    .S(net481),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _09300_ (.A0(net1380),
    .A1(net581),
    .S(net482),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(net1503),
    .A1(net578),
    .S(net480),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _09302_ (.A0(net1449),
    .A1(net573),
    .S(net482),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(net1455),
    .A1(net542),
    .S(net480),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(net1478),
    .A1(net540),
    .S(net479),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _09305_ (.A0(net1349),
    .A1(net525),
    .S(net480),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(net1530),
    .A1(net522),
    .S(net480),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(net1357),
    .A1(_03782_),
    .S(net480),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _09308_ (.A0(net1369),
    .A1(net406),
    .S(net480),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(net1351),
    .A1(net354),
    .S(net480),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(net1505),
    .A1(net350),
    .S(net479),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(net1350),
    .A1(net348),
    .S(net479),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _09312_ (.A0(net1379),
    .A1(net344),
    .S(net479),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(net1754),
    .A1(net339),
    .S(net479),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _09314_ (.A0(net1435),
    .A1(net337),
    .S(net479),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(net1368),
    .A1(net332),
    .S(net479),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _09316_ (.A0(net1864),
    .A1(net330),
    .S(net479),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(net2271),
    .A1(net325),
    .S(net481),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(net1390),
    .A1(net321),
    .S(net479),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(net1401),
    .A1(net319),
    .S(net479),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(net1400),
    .A1(net313),
    .S(net481),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(net1931),
    .A1(net310),
    .S(net481),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _09322_ (.A0(net1624),
    .A1(net307),
    .S(net481),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(net1410),
    .A1(net303),
    .S(net482),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(net1569),
    .A1(net299),
    .S(net482),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _09325_ (.A0(net1788),
    .A1(net295),
    .S(net481),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _09326_ (.A0(net1553),
    .A1(net291),
    .S(net481),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(net1743),
    .A1(net288),
    .S(net482),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _09328_ (.A0(net1605),
    .A1(net282),
    .S(net481),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(net1659),
    .A1(net280),
    .S(net481),
    .X(_00515_));
 sky130_fd_sc_hd__nor2_2 _09330_ (.A(_04273_),
    .B(_04281_),
    .Y(_04292_));
 sky130_fd_sc_hd__mux2_1 _09331_ (.A0(net1537),
    .A1(net586),
    .S(net477),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _09332_ (.A0(net1402),
    .A1(net585),
    .S(net477),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _09333_ (.A0(net1451),
    .A1(net582),
    .S(net477),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _09334_ (.A0(net1706),
    .A1(net577),
    .S(net476),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(net1359),
    .A1(net573),
    .S(net477),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _09336_ (.A0(net1394),
    .A1(net542),
    .S(net476),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(net1617),
    .A1(net539),
    .S(net475),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _09338_ (.A0(net1847),
    .A1(net525),
    .S(net475),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _09339_ (.A0(net1805),
    .A1(net522),
    .S(net475),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _09340_ (.A0(net1798),
    .A1(_03782_),
    .S(net475),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(net1790),
    .A1(net405),
    .S(net476),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(net1692),
    .A1(net354),
    .S(net476),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(net1557),
    .A1(net350),
    .S(net475),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(net1565),
    .A1(net347),
    .S(net475),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _09345_ (.A0(net1486),
    .A1(net343),
    .S(net475),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(net1580),
    .A1(net340),
    .S(net475),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _09347_ (.A0(net1784),
    .A1(net338),
    .S(net476),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(net1955),
    .A1(net333),
    .S(net475),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _09349_ (.A0(net1655),
    .A1(net330),
    .S(net475),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(net1797),
    .A1(net326),
    .S(net477),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _09351_ (.A0(net1630),
    .A1(net322),
    .S(net476),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(net1438),
    .A1(net319),
    .S(net476),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _09353_ (.A0(net1675),
    .A1(net314),
    .S(net477),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(net1378),
    .A1(net310),
    .S(net477),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(net1358),
    .A1(net307),
    .S(net477),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _09356_ (.A0(net1356),
    .A1(net303),
    .S(net478),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(net1562),
    .A1(net299),
    .S(net478),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _09358_ (.A0(net1584),
    .A1(net296),
    .S(net477),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _09359_ (.A0(net1417),
    .A1(net292),
    .S(net477),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(net1384),
    .A1(net287),
    .S(net478),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(net1786),
    .A1(_03870_),
    .S(net478),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _09362_ (.A0(net1903),
    .A1(net280),
    .S(net478),
    .X(_00547_));
 sky130_fd_sc_hd__and3b_4 _09363_ (.A_N(\latched_rd[1] ),
    .B(\latched_rd[0] ),
    .C(_04290_),
    .X(_04293_));
 sky130_fd_sc_hd__mux2_1 _09364_ (.A0(net2150),
    .A1(net586),
    .S(net401),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _09365_ (.A0(net2262),
    .A1(net584),
    .S(net401),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _09366_ (.A0(net1737),
    .A1(net581),
    .S(net402),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _09367_ (.A0(net1898),
    .A1(net577),
    .S(net400),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _09368_ (.A0(net1941),
    .A1(net573),
    .S(net402),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _09369_ (.A0(net1778),
    .A1(net542),
    .S(net400),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(net2092),
    .A1(net540),
    .S(net400),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _09371_ (.A0(net1823),
    .A1(net524),
    .S(net399),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _09372_ (.A0(net1928),
    .A1(net522),
    .S(net400),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _09373_ (.A0(net2115),
    .A1(net409),
    .S(net400),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _09374_ (.A0(net1920),
    .A1(net406),
    .S(net400),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _09375_ (.A0(net1899),
    .A1(net355),
    .S(net400),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _09376_ (.A0(net1684),
    .A1(net351),
    .S(net399),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _09377_ (.A0(net1762),
    .A1(net348),
    .S(net399),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _09378_ (.A0(net1843),
    .A1(net344),
    .S(net399),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(net1813),
    .A1(net339),
    .S(net399),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _09380_ (.A0(net1886),
    .A1(net337),
    .S(net399),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(net2004),
    .A1(net333),
    .S(net399),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(net1811),
    .A1(net330),
    .S(net399),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _09383_ (.A0(net2226),
    .A1(net325),
    .S(net401),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(net1803),
    .A1(net322),
    .S(net399),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(net1837),
    .A1(net316),
    .S(net399),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(net2085),
    .A1(net314),
    .S(net401),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(net2017),
    .A1(net311),
    .S(net401),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _09388_ (.A0(net2018),
    .A1(net307),
    .S(net401),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(net2332),
    .A1(net304),
    .S(net402),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(net2136),
    .A1(net300),
    .S(net402),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _09391_ (.A0(net1963),
    .A1(net295),
    .S(net401),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(net1989),
    .A1(net292),
    .S(net401),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(net2145),
    .A1(net288),
    .S(net402),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _09394_ (.A0(net2263),
    .A1(net282),
    .S(net401),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(net2361),
    .A1(net280),
    .S(net401),
    .X(_00579_));
 sky130_fd_sc_hd__or4bb_1 _09396_ (.A(net196),
    .B(net193),
    .C_N(net197),
    .D_N(net198),
    .X(_04294_));
 sky130_fd_sc_hd__nand4_1 _09397_ (.A(net267),
    .B(net1234),
    .C(net171),
    .D(net182),
    .Y(_04295_));
 sky130_fd_sc_hd__or4_1 _09398_ (.A(net190),
    .B(net194),
    .C(net192),
    .D(net195),
    .X(_04296_));
 sky130_fd_sc_hd__or4b_1 _09399_ (.A(net199),
    .B(net189),
    .C(net191),
    .D_N(net188),
    .X(_04297_));
 sky130_fd_sc_hd__or4_4 _09400_ (.A(_04294_),
    .B(_04295_),
    .C(_04296_),
    .D(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__nor3b_1 _09401_ (.A(_04298_),
    .B(net1113),
    .C_N(net176),
    .Y(_04299_));
 sky130_fd_sc_hd__and3_1 _09402_ (.A(net175),
    .B(net174),
    .C(_04299_),
    .X(_00580_));
 sky130_fd_sc_hd__and3_1 _09403_ (.A(net267),
    .B(net1233),
    .C(_02437_),
    .X(_04300_));
 sky130_fd_sc_hd__a31o_1 _09404_ (.A1(net1233),
    .A2(_02439_),
    .A3(_02440_),
    .B1(_04300_),
    .X(_00581_));
 sky130_fd_sc_hd__a21o_1 _09405_ (.A1(net1089),
    .A2(net1186),
    .B1(\count_instr[0] ),
    .X(_04301_));
 sky130_fd_sc_hd__and3_1 _09406_ (.A(net1089),
    .B(\count_instr[0] ),
    .C(net1184),
    .X(_04302_));
 sky130_fd_sc_hd__and3b_1 _09407_ (.A_N(_04302_),
    .B(net1231),
    .C(_04301_),
    .X(_00583_));
 sky130_fd_sc_hd__and4_1 _09408_ (.A(\cpu_state[1] ),
    .B(\count_instr[1] ),
    .C(\count_instr[0] ),
    .D(net1186),
    .X(_04303_));
 sky130_fd_sc_hd__nor2_1 _09409_ (.A(net1206),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__o21a_1 _09410_ (.A1(net2558),
    .A2(_04302_),
    .B1(_04304_),
    .X(_00584_));
 sky130_fd_sc_hd__and2_1 _09411_ (.A(\count_instr[2] ),
    .B(_04303_),
    .X(_04305_));
 sky130_fd_sc_hd__o21ai_1 _09412_ (.A1(net3028),
    .A2(_04303_),
    .B1(net1231),
    .Y(_04306_));
 sky130_fd_sc_hd__nor2_1 _09413_ (.A(_04305_),
    .B(_04306_),
    .Y(_00585_));
 sky130_fd_sc_hd__and3_1 _09414_ (.A(\count_instr[3] ),
    .B(\count_instr[2] ),
    .C(_04303_),
    .X(_04307_));
 sky130_fd_sc_hd__o21ai_1 _09415_ (.A1(net2982),
    .A2(_04305_),
    .B1(net1231),
    .Y(_04308_));
 sky130_fd_sc_hd__nor2_1 _09416_ (.A(_04307_),
    .B(_04308_),
    .Y(_00586_));
 sky130_fd_sc_hd__or2_1 _09417_ (.A(\count_instr[4] ),
    .B(_04307_),
    .X(_04309_));
 sky130_fd_sc_hd__and2_1 _09418_ (.A(\count_instr[4] ),
    .B(_04307_),
    .X(_04310_));
 sky130_fd_sc_hd__and3b_1 _09419_ (.A_N(_04310_),
    .B(net1231),
    .C(_04309_),
    .X(_00587_));
 sky130_fd_sc_hd__or2_1 _09420_ (.A(\count_instr[5] ),
    .B(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__and2_1 _09421_ (.A(\count_instr[5] ),
    .B(\count_instr[4] ),
    .X(_04312_));
 sky130_fd_sc_hd__and4_1 _09422_ (.A(\count_instr[3] ),
    .B(\count_instr[2] ),
    .C(_04303_),
    .D(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__and3b_1 _09423_ (.A_N(_04313_),
    .B(net1231),
    .C(_04311_),
    .X(_00588_));
 sky130_fd_sc_hd__and2_1 _09424_ (.A(\count_instr[6] ),
    .B(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__o21ai_1 _09425_ (.A1(net3053),
    .A2(_04313_),
    .B1(net1225),
    .Y(_04315_));
 sky130_fd_sc_hd__nor2_1 _09426_ (.A(_04314_),
    .B(_04315_),
    .Y(_00589_));
 sky130_fd_sc_hd__and3_1 _09427_ (.A(\count_instr[7] ),
    .B(\count_instr[6] ),
    .C(_04313_),
    .X(_04316_));
 sky130_fd_sc_hd__o21ai_1 _09428_ (.A1(net2973),
    .A2(_04314_),
    .B1(net1225),
    .Y(_04317_));
 sky130_fd_sc_hd__nor2_1 _09429_ (.A(_04316_),
    .B(_04317_),
    .Y(_00590_));
 sky130_fd_sc_hd__and4_1 _09430_ (.A(\count_instr[8] ),
    .B(\count_instr[7] ),
    .C(\count_instr[6] ),
    .D(_04313_),
    .X(_04318_));
 sky130_fd_sc_hd__o21ai_1 _09431_ (.A1(net2831),
    .A2(_04316_),
    .B1(net1225),
    .Y(_04319_));
 sky130_fd_sc_hd__nor2_1 _09432_ (.A(_04318_),
    .B(_04319_),
    .Y(_00591_));
 sky130_fd_sc_hd__and2_1 _09433_ (.A(\count_instr[9] ),
    .B(_04318_),
    .X(_04320_));
 sky130_fd_sc_hd__o21ai_1 _09434_ (.A1(\count_instr[9] ),
    .A2(_04318_),
    .B1(net1225),
    .Y(_04321_));
 sky130_fd_sc_hd__nor2_1 _09435_ (.A(_04320_),
    .B(_04321_),
    .Y(_00592_));
 sky130_fd_sc_hd__or2_1 _09436_ (.A(\count_instr[10] ),
    .B(_04320_),
    .X(_04322_));
 sky130_fd_sc_hd__and3_1 _09437_ (.A(\count_instr[10] ),
    .B(\count_instr[9] ),
    .C(_04318_),
    .X(_04323_));
 sky130_fd_sc_hd__and3b_1 _09438_ (.A_N(_04323_),
    .B(net1226),
    .C(_04322_),
    .X(_00593_));
 sky130_fd_sc_hd__or2_1 _09439_ (.A(\count_instr[11] ),
    .B(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__and4_1 _09440_ (.A(\count_instr[11] ),
    .B(\count_instr[10] ),
    .C(\count_instr[9] ),
    .D(_04318_),
    .X(_04325_));
 sky130_fd_sc_hd__and3b_1 _09441_ (.A_N(_04325_),
    .B(net1226),
    .C(_04324_),
    .X(_00594_));
 sky130_fd_sc_hd__and2_1 _09442_ (.A(\count_instr[12] ),
    .B(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__o21ai_1 _09443_ (.A1(net3065),
    .A2(_04325_),
    .B1(net1226),
    .Y(_04327_));
 sky130_fd_sc_hd__nor2_1 _09444_ (.A(_04326_),
    .B(_04327_),
    .Y(_00595_));
 sky130_fd_sc_hd__and3_1 _09445_ (.A(\count_instr[13] ),
    .B(\count_instr[12] ),
    .C(_04325_),
    .X(_04328_));
 sky130_fd_sc_hd__o21ai_1 _09446_ (.A1(net2974),
    .A2(_04326_),
    .B1(net1228),
    .Y(_04329_));
 sky130_fd_sc_hd__nor2_1 _09447_ (.A(_04328_),
    .B(_04329_),
    .Y(_00596_));
 sky130_fd_sc_hd__and4_1 _09448_ (.A(\count_instr[14] ),
    .B(\count_instr[13] ),
    .C(\count_instr[12] ),
    .D(_04325_),
    .X(_04330_));
 sky130_fd_sc_hd__o21ai_1 _09449_ (.A1(net2779),
    .A2(_04328_),
    .B1(net1228),
    .Y(_04331_));
 sky130_fd_sc_hd__nor2_1 _09450_ (.A(_04330_),
    .B(_04331_),
    .Y(_00597_));
 sky130_fd_sc_hd__and2_1 _09451_ (.A(\count_instr[15] ),
    .B(_04330_),
    .X(_04332_));
 sky130_fd_sc_hd__o21ai_1 _09452_ (.A1(net3042),
    .A2(_04330_),
    .B1(net1228),
    .Y(_04333_));
 sky130_fd_sc_hd__nor2_1 _09453_ (.A(_04332_),
    .B(_04333_),
    .Y(_00598_));
 sky130_fd_sc_hd__or2_1 _09454_ (.A(\count_instr[16] ),
    .B(_04332_),
    .X(_04334_));
 sky130_fd_sc_hd__nand2_1 _09455_ (.A(\count_instr[16] ),
    .B(_04332_),
    .Y(_04335_));
 sky130_fd_sc_hd__and3_1 _09456_ (.A(net1228),
    .B(_04334_),
    .C(_04335_),
    .X(_00599_));
 sky130_fd_sc_hd__and2_1 _09457_ (.A(\count_instr[17] ),
    .B(\count_instr[16] ),
    .X(_04336_));
 sky130_fd_sc_hd__and3_1 _09458_ (.A(\count_instr[15] ),
    .B(_04330_),
    .C(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__a211oi_1 _09459_ (.A1(_02376_),
    .A2(_04335_),
    .B1(_04337_),
    .C1(net1206),
    .Y(_00600_));
 sky130_fd_sc_hd__and4_1 _09460_ (.A(\count_instr[18] ),
    .B(\count_instr[15] ),
    .C(_04330_),
    .D(_04336_),
    .X(_04338_));
 sky130_fd_sc_hd__o21ai_1 _09461_ (.A1(net2774),
    .A2(_04337_),
    .B1(net1229),
    .Y(_04339_));
 sky130_fd_sc_hd__nor2_1 _09462_ (.A(_04338_),
    .B(_04339_),
    .Y(_00601_));
 sky130_fd_sc_hd__and2_1 _09463_ (.A(\count_instr[19] ),
    .B(_04338_),
    .X(_04340_));
 sky130_fd_sc_hd__o21ai_1 _09464_ (.A1(net3040),
    .A2(_04338_),
    .B1(net1229),
    .Y(_04341_));
 sky130_fd_sc_hd__nor2_1 _09465_ (.A(_04340_),
    .B(_04341_),
    .Y(_00602_));
 sky130_fd_sc_hd__and3_1 _09466_ (.A(\count_instr[20] ),
    .B(\count_instr[19] ),
    .C(_04338_),
    .X(_04342_));
 sky130_fd_sc_hd__o21ai_1 _09467_ (.A1(net2997),
    .A2(_04340_),
    .B1(net1229),
    .Y(_04343_));
 sky130_fd_sc_hd__nor2_1 _09468_ (.A(_04342_),
    .B(_04343_),
    .Y(_00603_));
 sky130_fd_sc_hd__and4_1 _09469_ (.A(\count_instr[21] ),
    .B(\count_instr[20] ),
    .C(\count_instr[19] ),
    .D(_04338_),
    .X(_04344_));
 sky130_fd_sc_hd__o21ai_1 _09470_ (.A1(net2825),
    .A2(_04342_),
    .B1(net1235),
    .Y(_04345_));
 sky130_fd_sc_hd__nor2_1 _09471_ (.A(_04344_),
    .B(_04345_),
    .Y(_00604_));
 sky130_fd_sc_hd__or2_1 _09472_ (.A(\count_instr[22] ),
    .B(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _09473_ (.A(\count_instr[22] ),
    .B(_04344_),
    .Y(_04347_));
 sky130_fd_sc_hd__and3_1 _09474_ (.A(net1235),
    .B(_04346_),
    .C(_04347_),
    .X(_00605_));
 sky130_fd_sc_hd__and2_1 _09475_ (.A(\count_instr[23] ),
    .B(\count_instr[22] ),
    .X(_04348_));
 sky130_fd_sc_hd__and2_1 _09476_ (.A(_04344_),
    .B(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__a211oi_1 _09477_ (.A1(_02375_),
    .A2(_04347_),
    .B1(_04349_),
    .C1(net1215),
    .Y(_00606_));
 sky130_fd_sc_hd__and3_1 _09478_ (.A(\count_instr[24] ),
    .B(_04344_),
    .C(_04348_),
    .X(_04350_));
 sky130_fd_sc_hd__o21ai_1 _09479_ (.A1(net2998),
    .A2(_04349_),
    .B1(net1239),
    .Y(_04351_));
 sky130_fd_sc_hd__nor2_1 _09480_ (.A(_04350_),
    .B(_04351_),
    .Y(_00607_));
 sky130_fd_sc_hd__and4_1 _09481_ (.A(\count_instr[25] ),
    .B(\count_instr[24] ),
    .C(_04344_),
    .D(_04348_),
    .X(_04352_));
 sky130_fd_sc_hd__o21ai_1 _09482_ (.A1(net2935),
    .A2(_04350_),
    .B1(net1239),
    .Y(_04353_));
 sky130_fd_sc_hd__nor2_1 _09483_ (.A(_04352_),
    .B(_04353_),
    .Y(_00608_));
 sky130_fd_sc_hd__and2_1 _09484_ (.A(\count_instr[26] ),
    .B(_04352_),
    .X(_04354_));
 sky130_fd_sc_hd__o21ai_1 _09485_ (.A1(net3066),
    .A2(_04352_),
    .B1(net1239),
    .Y(_04355_));
 sky130_fd_sc_hd__nor2_1 _09486_ (.A(_04354_),
    .B(_04355_),
    .Y(_00609_));
 sky130_fd_sc_hd__and3_1 _09487_ (.A(\count_instr[27] ),
    .B(\count_instr[26] ),
    .C(_04352_),
    .X(_04356_));
 sky130_fd_sc_hd__o21ai_1 _09488_ (.A1(net2976),
    .A2(_04354_),
    .B1(net1239),
    .Y(_04357_));
 sky130_fd_sc_hd__nor2_1 _09489_ (.A(_04356_),
    .B(_04357_),
    .Y(_00610_));
 sky130_fd_sc_hd__and4_1 _09490_ (.A(\count_instr[28] ),
    .B(\count_instr[27] ),
    .C(\count_instr[26] ),
    .D(_04352_),
    .X(_04358_));
 sky130_fd_sc_hd__o21ai_1 _09491_ (.A1(net2892),
    .A2(_04356_),
    .B1(net1239),
    .Y(_04359_));
 sky130_fd_sc_hd__nor2_1 _09492_ (.A(_04358_),
    .B(_04359_),
    .Y(_00611_));
 sky130_fd_sc_hd__a21oi_1 _09493_ (.A1(\count_instr[29] ),
    .A2(_04358_),
    .B1(net1209),
    .Y(_04360_));
 sky130_fd_sc_hd__o21a_1 _09494_ (.A1(net3047),
    .A2(_04358_),
    .B1(_04360_),
    .X(_00612_));
 sky130_fd_sc_hd__a21o_1 _09495_ (.A1(\count_instr[29] ),
    .A2(_04358_),
    .B1(\count_instr[30] ),
    .X(_04361_));
 sky130_fd_sc_hd__and3_1 _09496_ (.A(\count_instr[30] ),
    .B(\count_instr[29] ),
    .C(_04358_),
    .X(_04362_));
 sky130_fd_sc_hd__and3b_1 _09497_ (.A_N(_04362_),
    .B(net1239),
    .C(_04361_),
    .X(_00613_));
 sky130_fd_sc_hd__and4_2 _09498_ (.A(\count_instr[31] ),
    .B(\count_instr[30] ),
    .C(\count_instr[29] ),
    .D(_04358_),
    .X(_04363_));
 sky130_fd_sc_hd__o21ai_1 _09499_ (.A1(net2805),
    .A2(_04362_),
    .B1(net1239),
    .Y(_04364_));
 sky130_fd_sc_hd__nor2_1 _09500_ (.A(_04363_),
    .B(_04364_),
    .Y(_00614_));
 sky130_fd_sc_hd__a21oi_1 _09501_ (.A1(\count_instr[32] ),
    .A2(_04363_),
    .B1(net1207),
    .Y(_04365_));
 sky130_fd_sc_hd__o21a_1 _09502_ (.A1(\count_instr[32] ),
    .A2(_04363_),
    .B1(_04365_),
    .X(_00615_));
 sky130_fd_sc_hd__a21o_1 _09503_ (.A1(\count_instr[32] ),
    .A2(_04363_),
    .B1(\count_instr[33] ),
    .X(_04366_));
 sky130_fd_sc_hd__nand3_1 _09504_ (.A(\count_instr[33] ),
    .B(\count_instr[32] ),
    .C(_04363_),
    .Y(_04367_));
 sky130_fd_sc_hd__and3_1 _09505_ (.A(net1226),
    .B(_04366_),
    .C(_04367_),
    .X(_00616_));
 sky130_fd_sc_hd__and3_1 _09506_ (.A(\count_instr[34] ),
    .B(\count_instr[33] ),
    .C(\count_instr[32] ),
    .X(_04368_));
 sky130_fd_sc_hd__and2_1 _09507_ (.A(_04363_),
    .B(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__a211oi_1 _09508_ (.A1(_02374_),
    .A2(_04367_),
    .B1(_04369_),
    .C1(net1206),
    .Y(_00617_));
 sky130_fd_sc_hd__and3_1 _09509_ (.A(\count_instr[35] ),
    .B(_04363_),
    .C(_04368_),
    .X(_04370_));
 sky130_fd_sc_hd__o21ai_1 _09510_ (.A1(net2992),
    .A2(_04369_),
    .B1(net1226),
    .Y(_04371_));
 sky130_fd_sc_hd__nor2_1 _09511_ (.A(_04370_),
    .B(_04371_),
    .Y(_00618_));
 sky130_fd_sc_hd__and4_1 _09512_ (.A(\count_instr[36] ),
    .B(\count_instr[35] ),
    .C(_04363_),
    .D(_04368_),
    .X(_04372_));
 sky130_fd_sc_hd__o21ai_1 _09513_ (.A1(net2799),
    .A2(_04370_),
    .B1(net1226),
    .Y(_04373_));
 sky130_fd_sc_hd__nor2_1 _09514_ (.A(_04372_),
    .B(_04373_),
    .Y(_00619_));
 sky130_fd_sc_hd__a21oi_1 _09515_ (.A1(\count_instr[37] ),
    .A2(_04372_),
    .B1(net1206),
    .Y(_04374_));
 sky130_fd_sc_hd__o21a_1 _09516_ (.A1(net3060),
    .A2(_04372_),
    .B1(_04374_),
    .X(_00620_));
 sky130_fd_sc_hd__a21o_1 _09517_ (.A1(\count_instr[37] ),
    .A2(_04372_),
    .B1(\count_instr[38] ),
    .X(_04375_));
 sky130_fd_sc_hd__and3_1 _09518_ (.A(\count_instr[38] ),
    .B(\count_instr[37] ),
    .C(_04372_),
    .X(_04376_));
 sky130_fd_sc_hd__and3b_1 _09519_ (.A_N(_04376_),
    .B(net1226),
    .C(_04375_),
    .X(_00621_));
 sky130_fd_sc_hd__and4_1 _09520_ (.A(\count_instr[39] ),
    .B(\count_instr[38] ),
    .C(\count_instr[37] ),
    .D(_04372_),
    .X(_04377_));
 sky130_fd_sc_hd__o21ai_1 _09521_ (.A1(net2796),
    .A2(_04376_),
    .B1(net1226),
    .Y(_04378_));
 sky130_fd_sc_hd__nor2_1 _09522_ (.A(_04377_),
    .B(_04378_),
    .Y(_00622_));
 sky130_fd_sc_hd__a21oi_1 _09523_ (.A1(\count_instr[40] ),
    .A2(_04377_),
    .B1(net1214),
    .Y(_04379_));
 sky130_fd_sc_hd__o21a_1 _09524_ (.A1(\count_instr[40] ),
    .A2(_04377_),
    .B1(_04379_),
    .X(_00623_));
 sky130_fd_sc_hd__a21o_1 _09525_ (.A1(\count_instr[40] ),
    .A2(_04377_),
    .B1(\count_instr[41] ),
    .X(_04380_));
 sky130_fd_sc_hd__and3_1 _09526_ (.A(\count_instr[41] ),
    .B(\count_instr[40] ),
    .C(_04377_),
    .X(_04381_));
 sky130_fd_sc_hd__and3b_1 _09527_ (.A_N(_04381_),
    .B(net1227),
    .C(_04380_),
    .X(_00624_));
 sky130_fd_sc_hd__and4_1 _09528_ (.A(\count_instr[42] ),
    .B(\count_instr[41] ),
    .C(\count_instr[40] ),
    .D(_04377_),
    .X(_04382_));
 sky130_fd_sc_hd__o21ai_1 _09529_ (.A1(net2836),
    .A2(_04381_),
    .B1(net1227),
    .Y(_04383_));
 sky130_fd_sc_hd__nor2_1 _09530_ (.A(_04382_),
    .B(_04383_),
    .Y(_00625_));
 sky130_fd_sc_hd__a21oi_1 _09531_ (.A1(\count_instr[43] ),
    .A2(_04382_),
    .B1(net1214),
    .Y(_04384_));
 sky130_fd_sc_hd__o21a_1 _09532_ (.A1(\count_instr[43] ),
    .A2(_04382_),
    .B1(_04384_),
    .X(_00626_));
 sky130_fd_sc_hd__a21o_1 _09533_ (.A1(\count_instr[43] ),
    .A2(_04382_),
    .B1(\count_instr[44] ),
    .X(_04385_));
 sky130_fd_sc_hd__and3_1 _09534_ (.A(\count_instr[44] ),
    .B(\count_instr[43] ),
    .C(_04382_),
    .X(_04386_));
 sky130_fd_sc_hd__and3b_1 _09535_ (.A_N(_04386_),
    .B(net1227),
    .C(_04385_),
    .X(_00627_));
 sky130_fd_sc_hd__and4_1 _09536_ (.A(\count_instr[45] ),
    .B(\count_instr[44] ),
    .C(\count_instr[43] ),
    .D(_04382_),
    .X(_04387_));
 sky130_fd_sc_hd__o21ai_1 _09537_ (.A1(net2832),
    .A2(_04386_),
    .B1(net1227),
    .Y(_04388_));
 sky130_fd_sc_hd__nor2_1 _09538_ (.A(_04387_),
    .B(_04388_),
    .Y(_00628_));
 sky130_fd_sc_hd__a21oi_1 _09539_ (.A1(\count_instr[46] ),
    .A2(_04387_),
    .B1(net1214),
    .Y(_04389_));
 sky130_fd_sc_hd__o21a_1 _09540_ (.A1(\count_instr[46] ),
    .A2(_04387_),
    .B1(_04389_),
    .X(_00629_));
 sky130_fd_sc_hd__a21o_1 _09541_ (.A1(\count_instr[46] ),
    .A2(_04387_),
    .B1(\count_instr[47] ),
    .X(_04390_));
 sky130_fd_sc_hd__and3_1 _09542_ (.A(\count_instr[47] ),
    .B(\count_instr[46] ),
    .C(_04387_),
    .X(_04391_));
 sky130_fd_sc_hd__and3b_1 _09543_ (.A_N(_04391_),
    .B(net1230),
    .C(_04390_),
    .X(_00630_));
 sky130_fd_sc_hd__or2_1 _09544_ (.A(\count_instr[48] ),
    .B(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(\count_instr[48] ),
    .B(_04391_),
    .Y(_04393_));
 sky130_fd_sc_hd__and3_1 _09546_ (.A(net1230),
    .B(_04392_),
    .C(_04393_),
    .X(_00631_));
 sky130_fd_sc_hd__and2_1 _09547_ (.A(\count_instr[49] ),
    .B(\count_instr[48] ),
    .X(_04394_));
 sky130_fd_sc_hd__and4_1 _09548_ (.A(\count_instr[47] ),
    .B(\count_instr[46] ),
    .C(_04387_),
    .D(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__a211oi_1 _09549_ (.A1(_02373_),
    .A2(_04393_),
    .B1(_04395_),
    .C1(net1214),
    .Y(_00632_));
 sky130_fd_sc_hd__and2_1 _09550_ (.A(\count_instr[50] ),
    .B(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__o21ai_1 _09551_ (.A1(net3051),
    .A2(_04395_),
    .B1(net1230),
    .Y(_04397_));
 sky130_fd_sc_hd__nor2_1 _09552_ (.A(_04396_),
    .B(_04397_),
    .Y(_00633_));
 sky130_fd_sc_hd__and3_1 _09553_ (.A(\count_instr[51] ),
    .B(\count_instr[50] ),
    .C(_04395_),
    .X(_04398_));
 sky130_fd_sc_hd__o21ai_1 _09554_ (.A1(net2954),
    .A2(_04396_),
    .B1(net1230),
    .Y(_04399_));
 sky130_fd_sc_hd__nor2_1 _09555_ (.A(_04398_),
    .B(_04399_),
    .Y(_00634_));
 sky130_fd_sc_hd__or2_1 _09556_ (.A(\count_instr[52] ),
    .B(_04398_),
    .X(_04400_));
 sky130_fd_sc_hd__nand2_1 _09557_ (.A(\count_instr[52] ),
    .B(_04398_),
    .Y(_04401_));
 sky130_fd_sc_hd__and3_1 _09558_ (.A(net1237),
    .B(_04400_),
    .C(_04401_),
    .X(_00635_));
 sky130_fd_sc_hd__and2_1 _09559_ (.A(\count_instr[53] ),
    .B(\count_instr[52] ),
    .X(_04402_));
 sky130_fd_sc_hd__and4_1 _09560_ (.A(\count_instr[51] ),
    .B(\count_instr[50] ),
    .C(_04395_),
    .D(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__a211oi_1 _09561_ (.A1(_02372_),
    .A2(_04401_),
    .B1(_04403_),
    .C1(net1216),
    .Y(_00636_));
 sky130_fd_sc_hd__and2_1 _09562_ (.A(\count_instr[54] ),
    .B(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__o21ai_1 _09563_ (.A1(net3034),
    .A2(_04403_),
    .B1(net1240),
    .Y(_04405_));
 sky130_fd_sc_hd__nor2_1 _09564_ (.A(_04404_),
    .B(_04405_),
    .Y(_00637_));
 sky130_fd_sc_hd__and3_1 _09565_ (.A(\count_instr[55] ),
    .B(\count_instr[54] ),
    .C(_04403_),
    .X(_04406_));
 sky130_fd_sc_hd__o21ai_1 _09566_ (.A1(net3013),
    .A2(_04404_),
    .B1(net1240),
    .Y(_04407_));
 sky130_fd_sc_hd__nor2_1 _09567_ (.A(_04406_),
    .B(_04407_),
    .Y(_00638_));
 sky130_fd_sc_hd__and4_1 _09568_ (.A(\count_instr[56] ),
    .B(\count_instr[55] ),
    .C(\count_instr[54] ),
    .D(_04403_),
    .X(_04408_));
 sky130_fd_sc_hd__o21ai_1 _09569_ (.A1(net2889),
    .A2(_04406_),
    .B1(net1240),
    .Y(_04409_));
 sky130_fd_sc_hd__nor2_1 _09570_ (.A(_04408_),
    .B(_04409_),
    .Y(_00639_));
 sky130_fd_sc_hd__a21oi_1 _09571_ (.A1(\count_instr[57] ),
    .A2(_04408_),
    .B1(net1215),
    .Y(_04410_));
 sky130_fd_sc_hd__o21a_1 _09572_ (.A1(\count_instr[57] ),
    .A2(_04408_),
    .B1(_04410_),
    .X(_00640_));
 sky130_fd_sc_hd__a21o_1 _09573_ (.A1(\count_instr[57] ),
    .A2(_04408_),
    .B1(\count_instr[58] ),
    .X(_04411_));
 sky130_fd_sc_hd__and3_1 _09574_ (.A(\count_instr[58] ),
    .B(\count_instr[57] ),
    .C(_04408_),
    .X(_04412_));
 sky130_fd_sc_hd__and3b_1 _09575_ (.A_N(_04412_),
    .B(net1238),
    .C(_04411_),
    .X(_00641_));
 sky130_fd_sc_hd__and4_1 _09576_ (.A(\count_instr[59] ),
    .B(\count_instr[58] ),
    .C(\count_instr[57] ),
    .D(_04408_),
    .X(_04413_));
 sky130_fd_sc_hd__o21ai_1 _09577_ (.A1(net2855),
    .A2(_04412_),
    .B1(net1238),
    .Y(_04414_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(_04413_),
    .B(_04414_),
    .Y(_00642_));
 sky130_fd_sc_hd__a21oi_1 _09579_ (.A1(\count_instr[60] ),
    .A2(_04413_),
    .B1(net1209),
    .Y(_04415_));
 sky130_fd_sc_hd__o21a_1 _09580_ (.A1(\count_instr[60] ),
    .A2(_04413_),
    .B1(_04415_),
    .X(_00643_));
 sky130_fd_sc_hd__a21o_1 _09581_ (.A1(\count_instr[60] ),
    .A2(_04413_),
    .B1(\count_instr[61] ),
    .X(_04416_));
 sky130_fd_sc_hd__and3_1 _09582_ (.A(\count_instr[61] ),
    .B(\count_instr[60] ),
    .C(_04413_),
    .X(_04417_));
 sky130_fd_sc_hd__and3b_1 _09583_ (.A_N(_04417_),
    .B(net1238),
    .C(_04416_),
    .X(_00644_));
 sky130_fd_sc_hd__and4_1 _09584_ (.A(\count_instr[62] ),
    .B(\count_instr[61] ),
    .C(\count_instr[60] ),
    .D(_04413_),
    .X(_04418_));
 sky130_fd_sc_hd__o21ai_1 _09585_ (.A1(net2865),
    .A2(_04417_),
    .B1(net1238),
    .Y(_04419_));
 sky130_fd_sc_hd__nor2_1 _09586_ (.A(_04418_),
    .B(_04419_),
    .Y(_00645_));
 sky130_fd_sc_hd__o21ai_1 _09587_ (.A1(net1940),
    .A2(_04418_),
    .B1(net1238),
    .Y(_04420_));
 sky130_fd_sc_hd__a21oi_1 _09588_ (.A1(net1940),
    .A2(_04418_),
    .B1(_04420_),
    .Y(_00646_));
 sky130_fd_sc_hd__nor2_1 _09589_ (.A(net1089),
    .B(net1207),
    .Y(_04421_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(_03750_),
    .A1(\reg_next_pc[1] ),
    .S(net922),
    .X(_04422_));
 sky130_fd_sc_hd__a22o_1 _09591_ (.A1(\reg_pc[1] ),
    .A2(net878),
    .B1(_04422_),
    .B2(net848),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_2 _09592_ (.A0(_03752_),
    .A1(\reg_next_pc[2] ),
    .S(net923),
    .X(_04423_));
 sky130_fd_sc_hd__a22o_1 _09593_ (.A1(\reg_pc[2] ),
    .A2(net878),
    .B1(_04423_),
    .B2(net848),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_2 _09594_ (.A0(_03754_),
    .A1(\reg_next_pc[3] ),
    .S(net923),
    .X(_04424_));
 sky130_fd_sc_hd__a22o_1 _09595_ (.A1(\reg_pc[3] ),
    .A2(net878),
    .B1(_04424_),
    .B2(net848),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_2 _09596_ (.A0(_03757_),
    .A1(\reg_next_pc[4] ),
    .S(net923),
    .X(_04425_));
 sky130_fd_sc_hd__a22o_1 _09597_ (.A1(\reg_pc[4] ),
    .A2(net878),
    .B1(_04425_),
    .B2(net848),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _09598_ (.A0(_03762_),
    .A1(\reg_next_pc[5] ),
    .S(net923),
    .X(_04426_));
 sky130_fd_sc_hd__a22o_1 _09599_ (.A1(\reg_pc[5] ),
    .A2(net877),
    .B1(_04426_),
    .B2(net847),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_4 _09600_ (.A0(_03767_),
    .A1(\reg_next_pc[6] ),
    .S(net921),
    .X(_04427_));
 sky130_fd_sc_hd__a22o_1 _09601_ (.A1(\reg_pc[6] ),
    .A2(net876),
    .B1(_04427_),
    .B2(net846),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_2 _09602_ (.A0(_03770_),
    .A1(\reg_next_pc[7] ),
    .S(net921),
    .X(_04428_));
 sky130_fd_sc_hd__a22o_1 _09603_ (.A1(\reg_pc[7] ),
    .A2(net882),
    .B1(_04428_),
    .B2(net846),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_2 _09604_ (.A0(_03775_),
    .A1(\reg_next_pc[8] ),
    .S(net921),
    .X(_04429_));
 sky130_fd_sc_hd__a22o_1 _09605_ (.A1(\reg_pc[8] ),
    .A2(net876),
    .B1(_04429_),
    .B2(net846),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_2 _09606_ (.A0(_03778_),
    .A1(\reg_next_pc[9] ),
    .S(net927),
    .X(_04430_));
 sky130_fd_sc_hd__a22o_1 _09607_ (.A1(\reg_pc[9] ),
    .A2(net876),
    .B1(_04430_),
    .B2(net845),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_2 _09608_ (.A0(_03783_),
    .A1(\reg_next_pc[10] ),
    .S(net920),
    .X(_04431_));
 sky130_fd_sc_hd__a22o_1 _09609_ (.A1(\reg_pc[10] ),
    .A2(net876),
    .B1(_04431_),
    .B2(net845),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_2 _09610_ (.A0(_03786_),
    .A1(\reg_next_pc[11] ),
    .S(net920),
    .X(_04432_));
 sky130_fd_sc_hd__a22o_1 _09611_ (.A1(\reg_pc[11] ),
    .A2(net875),
    .B1(_04432_),
    .B2(net845),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_2 _09612_ (.A0(_03792_),
    .A1(\reg_next_pc[12] ),
    .S(net920),
    .X(_04433_));
 sky130_fd_sc_hd__a22o_1 _09613_ (.A1(\reg_pc[12] ),
    .A2(net875),
    .B1(_04433_),
    .B2(net845),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_2 _09614_ (.A0(_03795_),
    .A1(\reg_next_pc[13] ),
    .S(net920),
    .X(_04434_));
 sky130_fd_sc_hd__a22o_1 _09615_ (.A1(\reg_pc[13] ),
    .A2(net875),
    .B1(_04434_),
    .B2(net845),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_2 _09616_ (.A0(_03800_),
    .A1(\reg_next_pc[14] ),
    .S(net920),
    .X(_04435_));
 sky130_fd_sc_hd__a22o_1 _09617_ (.A1(\reg_pc[14] ),
    .A2(net875),
    .B1(_04435_),
    .B2(net845),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(_03803_),
    .A1(\reg_next_pc[15] ),
    .S(net920),
    .X(_04436_));
 sky130_fd_sc_hd__a22o_1 _09619_ (.A1(\reg_pc[15] ),
    .A2(net876),
    .B1(_04436_),
    .B2(net846),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _09620_ (.A0(_03808_),
    .A1(\reg_next_pc[16] ),
    .S(net922),
    .X(_04437_));
 sky130_fd_sc_hd__a22o_1 _09621_ (.A1(net3061),
    .A2(net877),
    .B1(_04437_),
    .B2(net847),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_4 _09622_ (.A0(_03811_),
    .A1(\reg_next_pc[17] ),
    .S(net922),
    .X(_04438_));
 sky130_fd_sc_hd__a22o_1 _09623_ (.A1(\reg_pc[17] ),
    .A2(net877),
    .B1(_04438_),
    .B2(net847),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_2 _09624_ (.A0(_03816_),
    .A1(\reg_next_pc[18] ),
    .S(net922),
    .X(_04439_));
 sky130_fd_sc_hd__a22o_1 _09625_ (.A1(\reg_pc[18] ),
    .A2(net877),
    .B1(_04439_),
    .B2(net847),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_2 _09626_ (.A0(_03819_),
    .A1(\reg_next_pc[19] ),
    .S(net922),
    .X(_04440_));
 sky130_fd_sc_hd__a22o_1 _09627_ (.A1(net3037),
    .A2(net877),
    .B1(_04440_),
    .B2(net847),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_2 _09628_ (.A0(_03824_),
    .A1(\reg_next_pc[20] ),
    .S(net926),
    .X(_04441_));
 sky130_fd_sc_hd__a22o_1 _09629_ (.A1(\reg_pc[20] ),
    .A2(net877),
    .B1(_04441_),
    .B2(net847),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_2 _09630_ (.A0(_03827_),
    .A1(\reg_next_pc[21] ),
    .S(net926),
    .X(_04442_));
 sky130_fd_sc_hd__a22o_1 _09631_ (.A1(\reg_pc[21] ),
    .A2(net881),
    .B1(_04442_),
    .B2(net851),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_2 _09632_ (.A0(_03832_),
    .A1(\reg_next_pc[22] ),
    .S(net926),
    .X(_04443_));
 sky130_fd_sc_hd__a22o_1 _09633_ (.A1(\reg_pc[22] ),
    .A2(net881),
    .B1(_04443_),
    .B2(net851),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_2 _09634_ (.A0(_03837_),
    .A1(\reg_next_pc[23] ),
    .S(net926),
    .X(_04444_));
 sky130_fd_sc_hd__a22o_1 _09635_ (.A1(net3059),
    .A2(net881),
    .B1(_04444_),
    .B2(net851),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_2 _09636_ (.A0(_03840_),
    .A1(\reg_next_pc[24] ),
    .S(net926),
    .X(_04445_));
 sky130_fd_sc_hd__a22o_1 _09637_ (.A1(\reg_pc[24] ),
    .A2(net881),
    .B1(_04445_),
    .B2(net851),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_2 _09638_ (.A0(_03845_),
    .A1(\reg_next_pc[25] ),
    .S(net924),
    .X(_04446_));
 sky130_fd_sc_hd__a22o_1 _09639_ (.A1(\reg_pc[25] ),
    .A2(net879),
    .B1(_04446_),
    .B2(net849),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_2 _09640_ (.A0(_03850_),
    .A1(\reg_next_pc[26] ),
    .S(net924),
    .X(_04447_));
 sky130_fd_sc_hd__a22o_1 _09641_ (.A1(\reg_pc[26] ),
    .A2(net879),
    .B1(_04447_),
    .B2(net849),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_2 _09642_ (.A0(_03853_),
    .A1(\reg_next_pc[27] ),
    .S(net925),
    .X(_04448_));
 sky130_fd_sc_hd__a22o_1 _09643_ (.A1(\reg_pc[27] ),
    .A2(net879),
    .B1(_04448_),
    .B2(net849),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_2 _09644_ (.A0(_03858_),
    .A1(\reg_next_pc[28] ),
    .S(net924),
    .X(_04449_));
 sky130_fd_sc_hd__a22o_1 _09645_ (.A1(\reg_pc[28] ),
    .A2(net880),
    .B1(_04449_),
    .B2(net850),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_2 _09646_ (.A0(_03861_),
    .A1(\reg_next_pc[29] ),
    .S(net924),
    .X(_04450_));
 sky130_fd_sc_hd__a22o_1 _09647_ (.A1(\reg_pc[29] ),
    .A2(net880),
    .B1(_04450_),
    .B2(net850),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _09648_ (.A0(_03866_),
    .A1(\reg_next_pc[30] ),
    .S(net924),
    .X(_04451_));
 sky130_fd_sc_hd__a22o_1 _09649_ (.A1(\reg_pc[30] ),
    .A2(net880),
    .B1(_04451_),
    .B2(net850),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _09650_ (.A0(_03871_),
    .A1(\reg_next_pc[31] ),
    .S(net924),
    .X(_04452_));
 sky130_fd_sc_hd__a22o_1 _09651_ (.A1(\reg_pc[31] ),
    .A2(net879),
    .B1(_04452_),
    .B2(net849),
    .X(_00677_));
 sky130_fd_sc_hd__and3_1 _09652_ (.A(net1182),
    .B(net1148),
    .C(\decoded_imm_j[1] ),
    .X(_04453_));
 sky130_fd_sc_hd__nand2_1 _09653_ (.A(_04422_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__or2_1 _09654_ (.A(_04422_),
    .B(_04453_),
    .X(_04455_));
 sky130_fd_sc_hd__a32o_1 _09655_ (.A1(net848),
    .A2(_04454_),
    .A3(_04455_),
    .B1(net878),
    .B2(net1330),
    .X(_00678_));
 sky130_fd_sc_hd__and2_1 _09656_ (.A(\decoded_imm_j[2] ),
    .B(_04423_),
    .X(_04456_));
 sky130_fd_sc_hd__xor2_1 _09657_ (.A(\decoded_imm_j[2] ),
    .B(_04423_),
    .X(_04457_));
 sky130_fd_sc_hd__a21o_1 _09658_ (.A1(\decoded_imm_j[1] ),
    .A2(_04422_),
    .B1(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__nand3_1 _09659_ (.A(\decoded_imm_j[1] ),
    .B(_04422_),
    .C(_04457_),
    .Y(_04459_));
 sky130_fd_sc_hd__nor2_1 _09660_ (.A(net1148),
    .B(_04423_),
    .Y(_04460_));
 sky130_fd_sc_hd__a311o_1 _09661_ (.A1(net1148),
    .A2(_04458_),
    .A3(_04459_),
    .B1(_04460_),
    .C1(_02380_),
    .X(_04461_));
 sky130_fd_sc_hd__or2_1 _09662_ (.A(net1187),
    .B(_04423_),
    .X(_04462_));
 sky130_fd_sc_hd__a32o_1 _09663_ (.A1(net848),
    .A2(_04461_),
    .A3(_04462_),
    .B1(net878),
    .B2(net2630),
    .X(_00679_));
 sky130_fd_sc_hd__nand2_1 _09664_ (.A(\decoded_imm_j[3] ),
    .B(_04424_),
    .Y(_04463_));
 sky130_fd_sc_hd__or2_1 _09665_ (.A(\decoded_imm_j[3] ),
    .B(_04424_),
    .X(_04464_));
 sky130_fd_sc_hd__and2_1 _09666_ (.A(_04463_),
    .B(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__a31o_1 _09667_ (.A1(\decoded_imm_j[1] ),
    .A2(_04422_),
    .A3(_04457_),
    .B1(_04456_),
    .X(_04466_));
 sky130_fd_sc_hd__nand2_1 _09668_ (.A(_04465_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__or2_1 _09669_ (.A(_04465_),
    .B(_04466_),
    .X(_04468_));
 sky130_fd_sc_hd__and2_1 _09670_ (.A(_04467_),
    .B(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__a2bb2o_1 _09671_ (.A1_N(_04460_),
    .A2_N(_02479_),
    .B1(net848),
    .B2(_04424_),
    .X(_04470_));
 sky130_fd_sc_hd__nand2_1 _09672_ (.A(_04423_),
    .B(_04424_),
    .Y(_04471_));
 sky130_fd_sc_hd__o221a_1 _09673_ (.A1(_02481_),
    .A2(_04469_),
    .B1(_04471_),
    .B2(_02489_),
    .C1(_04470_),
    .X(_04472_));
 sky130_fd_sc_hd__a21o_1 _09674_ (.A1(net2651),
    .A2(net878),
    .B1(_04472_),
    .X(_00680_));
 sky130_fd_sc_hd__nand2_1 _09675_ (.A(_04463_),
    .B(_04467_),
    .Y(_04473_));
 sky130_fd_sc_hd__or2_1 _09676_ (.A(\decoded_imm_j[4] ),
    .B(_04425_),
    .X(_04474_));
 sky130_fd_sc_hd__and2_1 _09677_ (.A(\decoded_imm_j[4] ),
    .B(_04425_),
    .X(_04475_));
 sky130_fd_sc_hd__inv_2 _09678_ (.A(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__and3_1 _09679_ (.A(_04473_),
    .B(_04474_),
    .C(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__a21oi_1 _09680_ (.A1(_04474_),
    .A2(_04476_),
    .B1(_04473_),
    .Y(_04478_));
 sky130_fd_sc_hd__o21ai_1 _09681_ (.A1(_04477_),
    .A2(_04478_),
    .B1(_02480_),
    .Y(_04479_));
 sky130_fd_sc_hd__xnor2_1 _09682_ (.A(_04425_),
    .B(_04471_),
    .Y(_04480_));
 sky130_fd_sc_hd__o221a_1 _09683_ (.A1(net1187),
    .A2(_04425_),
    .B1(_04480_),
    .B2(_02489_),
    .C1(net848),
    .X(_04481_));
 sky130_fd_sc_hd__a22o_1 _09684_ (.A1(net2740),
    .A2(net878),
    .B1(_04479_),
    .B2(_04481_),
    .X(_00681_));
 sky130_fd_sc_hd__nor2_1 _09685_ (.A(\decoded_imm_j[5] ),
    .B(_04426_),
    .Y(_04482_));
 sky130_fd_sc_hd__and2_1 _09686_ (.A(\decoded_imm_j[5] ),
    .B(_04426_),
    .X(_04483_));
 sky130_fd_sc_hd__nor2_1 _09687_ (.A(_04482_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__nand3_1 _09688_ (.A(_04463_),
    .B(_04467_),
    .C(_04476_),
    .Y(_04485_));
 sky130_fd_sc_hd__a21oi_1 _09689_ (.A1(_04474_),
    .A2(_04485_),
    .B1(_04484_),
    .Y(_04486_));
 sky130_fd_sc_hd__a31o_1 _09690_ (.A1(_04474_),
    .A2(_04484_),
    .A3(_04485_),
    .B1(net984),
    .X(_04487_));
 sky130_fd_sc_hd__and4_2 _09691_ (.A(_04423_),
    .B(_04424_),
    .C(_04425_),
    .D(_04426_),
    .X(_04488_));
 sky130_fd_sc_hd__a31o_1 _09692_ (.A1(_04423_),
    .A2(_04424_),
    .A3(_04425_),
    .B1(_04426_),
    .X(_04489_));
 sky130_fd_sc_hd__or3b_1 _09693_ (.A(net1149),
    .B(_04488_),
    .C_N(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__o211a_1 _09694_ (.A1(_04486_),
    .A2(_04487_),
    .B1(_04490_),
    .C1(net1182),
    .X(_04491_));
 sky130_fd_sc_hd__o21ai_1 _09695_ (.A1(net1182),
    .A2(_04426_),
    .B1(net848),
    .Y(_04492_));
 sky130_fd_sc_hd__a2bb2o_1 _09696_ (.A1_N(_04491_),
    .A2_N(_04492_),
    .B1(net2821),
    .B2(net878),
    .X(_00682_));
 sky130_fd_sc_hd__or2_1 _09697_ (.A(\decoded_imm_j[6] ),
    .B(_04427_),
    .X(_04493_));
 sky130_fd_sc_hd__and2_1 _09698_ (.A(\decoded_imm_j[6] ),
    .B(_04427_),
    .X(_04494_));
 sky130_fd_sc_hd__nand2_1 _09699_ (.A(\decoded_imm_j[6] ),
    .B(_04427_),
    .Y(_04495_));
 sky130_fd_sc_hd__nand2_1 _09700_ (.A(_04493_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__a31o_1 _09701_ (.A1(_04474_),
    .A2(_04484_),
    .A3(_04485_),
    .B1(_04483_),
    .X(_04497_));
 sky130_fd_sc_hd__a21oi_1 _09702_ (.A1(_04496_),
    .A2(_04497_),
    .B1(_02481_),
    .Y(_04498_));
 sky130_fd_sc_hd__o21a_1 _09703_ (.A1(_04496_),
    .A2(_04497_),
    .B1(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__xor2_1 _09704_ (.A(_04427_),
    .B(_04488_),
    .X(_04500_));
 sky130_fd_sc_hd__o221ai_1 _09705_ (.A1(net1183),
    .A2(_04427_),
    .B1(_04500_),
    .B2(_02489_),
    .C1(net846),
    .Y(_04501_));
 sky130_fd_sc_hd__a2bb2o_1 _09706_ (.A1_N(_04499_),
    .A2_N(_04501_),
    .B1(net2593),
    .B2(net876),
    .X(_00683_));
 sky130_fd_sc_hd__and2_1 _09707_ (.A(\decoded_imm_j[7] ),
    .B(_04428_),
    .X(_04502_));
 sky130_fd_sc_hd__or2_1 _09708_ (.A(\decoded_imm_j[7] ),
    .B(_04428_),
    .X(_04503_));
 sky130_fd_sc_hd__nand2b_1 _09709_ (.A_N(_04502_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__o21a_1 _09710_ (.A1(_04494_),
    .A2(_04497_),
    .B1(_04493_),
    .X(_04505_));
 sky130_fd_sc_hd__xnor2_1 _09711_ (.A(_04504_),
    .B(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__a21oi_1 _09712_ (.A1(_04427_),
    .A2(_04488_),
    .B1(_04428_),
    .Y(_04507_));
 sky130_fd_sc_hd__a31o_1 _09713_ (.A1(_04427_),
    .A2(_04428_),
    .A3(_04488_),
    .B1(net1149),
    .X(_04508_));
 sky130_fd_sc_hd__a2bb2o_1 _09714_ (.A1_N(_04507_),
    .A2_N(_04508_),
    .B1(net1149),
    .B2(_04506_),
    .X(_04509_));
 sky130_fd_sc_hd__mux2_1 _09715_ (.A0(_04428_),
    .A1(_04509_),
    .S(net1183),
    .X(_04510_));
 sky130_fd_sc_hd__a22o_1 _09716_ (.A1(net2560),
    .A2(net876),
    .B1(_04510_),
    .B2(net852),
    .X(_00684_));
 sky130_fd_sc_hd__and2_1 _09717_ (.A(\decoded_imm_j[8] ),
    .B(_04429_),
    .X(_04511_));
 sky130_fd_sc_hd__or2_1 _09718_ (.A(\decoded_imm_j[8] ),
    .B(_04429_),
    .X(_04512_));
 sky130_fd_sc_hd__and2b_1 _09719_ (.A_N(_04511_),
    .B(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__a21oi_1 _09720_ (.A1(_04503_),
    .A2(_04505_),
    .B1(_04502_),
    .Y(_04514_));
 sky130_fd_sc_hd__xnor2_1 _09721_ (.A(_04513_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__nand4_2 _09722_ (.A(_04427_),
    .B(_04428_),
    .C(_04429_),
    .D(_04488_),
    .Y(_04516_));
 sky130_fd_sc_hd__a31o_1 _09723_ (.A1(_04427_),
    .A2(_04428_),
    .A3(_04488_),
    .B1(_04429_),
    .X(_04517_));
 sky130_fd_sc_hd__a31o_1 _09724_ (.A1(net984),
    .A2(_04516_),
    .A3(_04517_),
    .B1(_02380_),
    .X(_04518_));
 sky130_fd_sc_hd__a21o_1 _09725_ (.A1(net1149),
    .A2(_04515_),
    .B1(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__or2_1 _09726_ (.A(net1183),
    .B(_04429_),
    .X(_04520_));
 sky130_fd_sc_hd__a32o_1 _09727_ (.A1(net846),
    .A2(_04519_),
    .A3(_04520_),
    .B1(net876),
    .B2(net2256),
    .X(_00685_));
 sky130_fd_sc_hd__or2_1 _09728_ (.A(_04503_),
    .B(_04511_),
    .X(_04521_));
 sky130_fd_sc_hd__o311a_1 _09729_ (.A1(_04502_),
    .A2(_04505_),
    .A3(_04511_),
    .B1(_04512_),
    .C1(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__or2_1 _09730_ (.A(\decoded_imm_j[9] ),
    .B(_04430_),
    .X(_04523_));
 sky130_fd_sc_hd__nand2_1 _09731_ (.A(\decoded_imm_j[9] ),
    .B(_04430_),
    .Y(_04524_));
 sky130_fd_sc_hd__and2_1 _09732_ (.A(_04523_),
    .B(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__nand2_1 _09733_ (.A(_04522_),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__inv_2 _09734_ (.A(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__or2_1 _09735_ (.A(_04522_),
    .B(_04525_),
    .X(_04528_));
 sky130_fd_sc_hd__nand2b_1 _09736_ (.A_N(_04516_),
    .B(_04430_),
    .Y(_04529_));
 sky130_fd_sc_hd__nand2b_1 _09737_ (.A_N(_04430_),
    .B(_04516_),
    .Y(_04530_));
 sky130_fd_sc_hd__a31o_1 _09738_ (.A1(net984),
    .A2(_04529_),
    .A3(_04530_),
    .B1(_02380_),
    .X(_04531_));
 sky130_fd_sc_hd__a31o_1 _09739_ (.A1(net1149),
    .A2(_04526_),
    .A3(_04528_),
    .B1(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__or2_1 _09740_ (.A(net1183),
    .B(_04430_),
    .X(_04533_));
 sky130_fd_sc_hd__a32o_1 _09741_ (.A1(net845),
    .A2(_04532_),
    .A3(_04533_),
    .B1(net875),
    .B2(net2638),
    .X(_00686_));
 sky130_fd_sc_hd__nand2_1 _09742_ (.A(\decoded_imm_j[10] ),
    .B(_04431_),
    .Y(_04534_));
 sky130_fd_sc_hd__or2_1 _09743_ (.A(\decoded_imm_j[10] ),
    .B(_04431_),
    .X(_04535_));
 sky130_fd_sc_hd__nand2_1 _09744_ (.A(_04534_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__nand2_1 _09745_ (.A(_04524_),
    .B(_04526_),
    .Y(_04537_));
 sky130_fd_sc_hd__o21ai_1 _09746_ (.A1(_04536_),
    .A2(_04537_),
    .B1(_02480_),
    .Y(_04538_));
 sky130_fd_sc_hd__a21o_1 _09747_ (.A1(_04536_),
    .A2(_04537_),
    .B1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__and2b_1 _09748_ (.A_N(_04529_),
    .B(_04431_),
    .X(_04540_));
 sky130_fd_sc_hd__xnor2_1 _09749_ (.A(_04431_),
    .B(_04529_),
    .Y(_04541_));
 sky130_fd_sc_hd__o221a_1 _09750_ (.A1(net1183),
    .A2(_04431_),
    .B1(_04541_),
    .B2(_02489_),
    .C1(net846),
    .X(_04542_));
 sky130_fd_sc_hd__a22o_1 _09751_ (.A1(net2689),
    .A2(net875),
    .B1(_04539_),
    .B2(_04542_),
    .X(_00687_));
 sky130_fd_sc_hd__and2_1 _09752_ (.A(\decoded_imm_j[11] ),
    .B(_04432_),
    .X(_04543_));
 sky130_fd_sc_hd__nor2_1 _09753_ (.A(\decoded_imm_j[11] ),
    .B(_04432_),
    .Y(_04544_));
 sky130_fd_sc_hd__nor2_1 _09754_ (.A(_04543_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand2_1 _09755_ (.A(_04524_),
    .B(_04534_),
    .Y(_04546_));
 sky130_fd_sc_hd__nand2_1 _09756_ (.A(_04535_),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__o21ai_1 _09757_ (.A1(_04527_),
    .A2(_04546_),
    .B1(_04535_),
    .Y(_04548_));
 sky130_fd_sc_hd__and2b_1 _09758_ (.A_N(_04548_),
    .B(_04545_),
    .X(_04549_));
 sky130_fd_sc_hd__xnor2_1 _09759_ (.A(_04545_),
    .B(_04548_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand4b_1 _09760_ (.A_N(_04516_),
    .B(_04432_),
    .C(_04431_),
    .D(_04430_),
    .Y(_04551_));
 sky130_fd_sc_hd__or2_1 _09761_ (.A(_04432_),
    .B(_04540_),
    .X(_04552_));
 sky130_fd_sc_hd__a31o_1 _09762_ (.A1(net984),
    .A2(_04551_),
    .A3(_04552_),
    .B1(_02380_),
    .X(_04553_));
 sky130_fd_sc_hd__a21o_1 _09763_ (.A1(net1149),
    .A2(_04550_),
    .B1(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__or2_1 _09764_ (.A(net1183),
    .B(_04432_),
    .X(_04555_));
 sky130_fd_sc_hd__a32o_1 _09765_ (.A1(net845),
    .A2(_04554_),
    .A3(_04555_),
    .B1(net875),
    .B2(net2446),
    .X(_00688_));
 sky130_fd_sc_hd__or2_1 _09766_ (.A(\decoded_imm_j[12] ),
    .B(_04433_),
    .X(_04556_));
 sky130_fd_sc_hd__nand2_1 _09767_ (.A(\decoded_imm_j[12] ),
    .B(_04433_),
    .Y(_04557_));
 sky130_fd_sc_hd__and2_1 _09768_ (.A(_04556_),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__o21ai_1 _09769_ (.A1(_04543_),
    .A2(_04549_),
    .B1(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__o31a_1 _09770_ (.A1(_04543_),
    .A2(_04549_),
    .A3(_04558_),
    .B1(net1149),
    .X(_04560_));
 sky130_fd_sc_hd__nand2b_1 _09771_ (.A_N(_04551_),
    .B(_04433_),
    .Y(_04561_));
 sky130_fd_sc_hd__nand2b_1 _09772_ (.A_N(_04433_),
    .B(_04551_),
    .Y(_04562_));
 sky130_fd_sc_hd__a32o_1 _09773_ (.A1(net984),
    .A2(_04561_),
    .A3(_04562_),
    .B1(_04559_),
    .B2(_04560_),
    .X(_04563_));
 sky130_fd_sc_hd__mux2_1 _09774_ (.A0(_04433_),
    .A1(_04563_),
    .S(net1183),
    .X(_04564_));
 sky130_fd_sc_hd__a22o_1 _09775_ (.A1(net2675),
    .A2(net875),
    .B1(_04564_),
    .B2(net845),
    .X(_00689_));
 sky130_fd_sc_hd__nor2_1 _09776_ (.A(\decoded_imm_j[13] ),
    .B(_04434_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _09777_ (.A(\decoded_imm_j[13] ),
    .B(_04434_),
    .Y(_04566_));
 sky130_fd_sc_hd__and2b_1 _09778_ (.A_N(_04565_),
    .B(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__nand2_1 _09779_ (.A(_04545_),
    .B(_04558_),
    .Y(_04568_));
 sky130_fd_sc_hd__inv_2 _09780_ (.A(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__and3_1 _09781_ (.A(_04525_),
    .B(_04534_),
    .C(_04535_),
    .X(_04570_));
 sky130_fd_sc_hd__or3_1 _09782_ (.A(_04526_),
    .B(_04536_),
    .C(_04568_),
    .X(_04571_));
 sky130_fd_sc_hd__nand2b_1 _09783_ (.A_N(_04543_),
    .B(_04557_),
    .Y(_04572_));
 sky130_fd_sc_hd__o2bb2a_1 _09784_ (.A1_N(_04556_),
    .A2_N(_04572_),
    .B1(_04568_),
    .B2(_04547_),
    .X(_04573_));
 sky130_fd_sc_hd__and2_1 _09785_ (.A(_04571_),
    .B(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__xor2_1 _09786_ (.A(_04567_),
    .B(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__nand2_1 _09787_ (.A(_02480_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__nand2b_1 _09788_ (.A_N(_04561_),
    .B(_04434_),
    .Y(_04577_));
 sky130_fd_sc_hd__xnor2_1 _09789_ (.A(_04434_),
    .B(_04561_),
    .Y(_04578_));
 sky130_fd_sc_hd__o221a_1 _09790_ (.A1(net1183),
    .A2(_04434_),
    .B1(_04578_),
    .B2(_02489_),
    .C1(net846),
    .X(_04579_));
 sky130_fd_sc_hd__a22o_1 _09791_ (.A1(net2741),
    .A2(net875),
    .B1(_04576_),
    .B2(_04579_),
    .X(_00690_));
 sky130_fd_sc_hd__or2_1 _09792_ (.A(\decoded_imm_j[14] ),
    .B(_04435_),
    .X(_04580_));
 sky130_fd_sc_hd__nand2_1 _09793_ (.A(\decoded_imm_j[14] ),
    .B(_04435_),
    .Y(_04581_));
 sky130_fd_sc_hd__and2_1 _09794_ (.A(_04580_),
    .B(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__o21ai_1 _09795_ (.A1(_04565_),
    .A2(_04574_),
    .B1(_04566_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _09796_ (.A(_04582_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__o21a_1 _09797_ (.A1(_04582_),
    .A2(_04583_),
    .B1(net1149),
    .X(_04585_));
 sky130_fd_sc_hd__nand2b_1 _09798_ (.A_N(_04577_),
    .B(_04435_),
    .Y(_04586_));
 sky130_fd_sc_hd__xnor2_1 _09799_ (.A(_04435_),
    .B(_04577_),
    .Y(_04587_));
 sky130_fd_sc_hd__a22o_1 _09800_ (.A1(_04584_),
    .A2(_04585_),
    .B1(_04587_),
    .B2(net984),
    .X(_04588_));
 sky130_fd_sc_hd__mux2_1 _09801_ (.A0(_04435_),
    .A1(_04588_),
    .S(net1183),
    .X(_04589_));
 sky130_fd_sc_hd__a22o_1 _09802_ (.A1(net2642),
    .A2(net875),
    .B1(_04589_),
    .B2(net845),
    .X(_00691_));
 sky130_fd_sc_hd__nand2_1 _09803_ (.A(\decoded_imm_j[15] ),
    .B(_04436_),
    .Y(_04590_));
 sky130_fd_sc_hd__or2_1 _09804_ (.A(\decoded_imm_j[15] ),
    .B(_04436_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_1 _09805_ (.A(_04590_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__inv_2 _09806_ (.A(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__nand2_1 _09807_ (.A(_04566_),
    .B(_04581_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _09808_ (.A(_04567_),
    .B(_04582_),
    .Y(_04595_));
 sky130_fd_sc_hd__a2bb2o_1 _09809_ (.A1_N(_04573_),
    .A2_N(_04595_),
    .B1(_04594_),
    .B2(_04580_),
    .X(_04596_));
 sky130_fd_sc_hd__o21ba_1 _09810_ (.A1(_04571_),
    .A2(_04595_),
    .B1_N(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__xnor2_1 _09811_ (.A(_04592_),
    .B(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_1 _09812_ (.A(_02480_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__and2b_1 _09813_ (.A_N(_04586_),
    .B(_04436_),
    .X(_04600_));
 sky130_fd_sc_hd__and2b_1 _09814_ (.A_N(_04436_),
    .B(_04586_),
    .X(_04601_));
 sky130_fd_sc_hd__nor2_1 _09815_ (.A(_04600_),
    .B(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__o221a_1 _09816_ (.A1(net1183),
    .A2(_04436_),
    .B1(_04602_),
    .B2(_02489_),
    .C1(net846),
    .X(_04603_));
 sky130_fd_sc_hd__a22o_1 _09817_ (.A1(net2617),
    .A2(net876),
    .B1(_04599_),
    .B2(_04603_),
    .X(_00692_));
 sky130_fd_sc_hd__nand2_1 _09818_ (.A(\decoded_imm_j[16] ),
    .B(_04437_),
    .Y(_04604_));
 sky130_fd_sc_hd__or2_1 _09819_ (.A(\decoded_imm_j[16] ),
    .B(_04437_),
    .X(_04605_));
 sky130_fd_sc_hd__and2_1 _09820_ (.A(_04604_),
    .B(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__o21ai_1 _09821_ (.A1(_04592_),
    .A2(_04597_),
    .B1(_04590_),
    .Y(_04607_));
 sky130_fd_sc_hd__o211a_1 _09822_ (.A1(_04592_),
    .A2(_04597_),
    .B1(_04606_),
    .C1(_04590_),
    .X(_04608_));
 sky130_fd_sc_hd__and2b_1 _09823_ (.A_N(_04606_),
    .B(_04607_),
    .X(_04609_));
 sky130_fd_sc_hd__or3_1 _09824_ (.A(_02481_),
    .B(_04608_),
    .C(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__and2_1 _09825_ (.A(_04437_),
    .B(_04600_),
    .X(_04611_));
 sky130_fd_sc_hd__nor2_1 _09826_ (.A(_04437_),
    .B(_04600_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_1 _09827_ (.A(_04611_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__o221a_1 _09828_ (.A1(net1182),
    .A2(_04437_),
    .B1(_04613_),
    .B2(_02489_),
    .C1(net847),
    .X(_04614_));
 sky130_fd_sc_hd__a22o_1 _09829_ (.A1(net2569),
    .A2(net877),
    .B1(_04610_),
    .B2(_04614_),
    .X(_00693_));
 sky130_fd_sc_hd__xnor2_1 _09830_ (.A(\decoded_imm_j[17] ),
    .B(_04438_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand2_1 _09831_ (.A(_04590_),
    .B(_04604_),
    .Y(_04616_));
 sky130_fd_sc_hd__a32o_1 _09832_ (.A1(_04593_),
    .A2(_04596_),
    .A3(_04606_),
    .B1(_04616_),
    .B2(_04605_),
    .X(_04617_));
 sky130_fd_sc_hd__and4_1 _09833_ (.A(_04567_),
    .B(_04582_),
    .C(_04593_),
    .D(_04606_),
    .X(_04618_));
 sky130_fd_sc_hd__and4_1 _09834_ (.A(_04522_),
    .B(_04569_),
    .C(_04570_),
    .D(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__nor2_1 _09835_ (.A(_04617_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _09836_ (.A(_04615_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__a21o_1 _09837_ (.A1(_04615_),
    .A2(_04620_),
    .B1(net984),
    .X(_04622_));
 sky130_fd_sc_hd__nand2_1 _09838_ (.A(_04438_),
    .B(_04611_),
    .Y(_04623_));
 sky130_fd_sc_hd__or2_1 _09839_ (.A(_04438_),
    .B(_04611_),
    .X(_04624_));
 sky130_fd_sc_hd__nand3_1 _09840_ (.A(net984),
    .B(_04623_),
    .C(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__o211a_1 _09841_ (.A1(_04621_),
    .A2(_04622_),
    .B1(_04625_),
    .C1(net1182),
    .X(_04626_));
 sky130_fd_sc_hd__o21ai_1 _09842_ (.A1(net1182),
    .A2(_04438_),
    .B1(net847),
    .Y(_04627_));
 sky130_fd_sc_hd__a2bb2o_1 _09843_ (.A1_N(_04626_),
    .A2_N(_04627_),
    .B1(net2667),
    .B2(net877),
    .X(_00694_));
 sky130_fd_sc_hd__nand2_1 _09844_ (.A(\decoded_imm_j[18] ),
    .B(_04439_),
    .Y(_04628_));
 sky130_fd_sc_hd__or2_1 _09845_ (.A(\decoded_imm_j[18] ),
    .B(_04439_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _09846_ (.A(_04628_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__a21o_1 _09847_ (.A1(\decoded_imm_j[17] ),
    .A2(_04438_),
    .B1(_04621_),
    .X(_04631_));
 sky130_fd_sc_hd__xnor2_1 _09848_ (.A(_04630_),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(net1146),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__and3_1 _09850_ (.A(_04438_),
    .B(_04439_),
    .C(_04611_),
    .X(_04634_));
 sky130_fd_sc_hd__a21oi_1 _09851_ (.A1(_04438_),
    .A2(_04611_),
    .B1(_04439_),
    .Y(_04635_));
 sky130_fd_sc_hd__o311ai_1 _09852_ (.A1(net1146),
    .A2(_04634_),
    .A3(_04635_),
    .B1(_04633_),
    .C1(net1182),
    .Y(_04636_));
 sky130_fd_sc_hd__or2_1 _09853_ (.A(net1182),
    .B(_04439_),
    .X(_04637_));
 sky130_fd_sc_hd__a32o_1 _09854_ (.A1(net847),
    .A2(_04636_),
    .A3(_04637_),
    .B1(net877),
    .B2(net2420),
    .X(_00695_));
 sky130_fd_sc_hd__and2_1 _09855_ (.A(\decoded_imm_j[19] ),
    .B(_04440_),
    .X(_04638_));
 sky130_fd_sc_hd__nor2_1 _09856_ (.A(\decoded_imm_j[19] ),
    .B(_04440_),
    .Y(_04639_));
 sky130_fd_sc_hd__nor2_1 _09857_ (.A(_04638_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__a22o_1 _09858_ (.A1(\decoded_imm_j[17] ),
    .A2(_04438_),
    .B1(_04439_),
    .B2(\decoded_imm_j[18] ),
    .X(_04641_));
 sky130_fd_sc_hd__or2_1 _09859_ (.A(_04621_),
    .B(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__a21oi_1 _09860_ (.A1(_04629_),
    .A2(_04642_),
    .B1(_04640_),
    .Y(_04643_));
 sky130_fd_sc_hd__and3_1 _09861_ (.A(_04629_),
    .B(_04640_),
    .C(_04642_),
    .X(_04644_));
 sky130_fd_sc_hd__nand2_1 _09862_ (.A(_04439_),
    .B(_04440_),
    .Y(_04645_));
 sky130_fd_sc_hd__nor2_1 _09863_ (.A(_04623_),
    .B(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__nor2_1 _09864_ (.A(net1146),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__o21ai_1 _09865_ (.A1(_04440_),
    .A2(_04634_),
    .B1(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__o31ai_1 _09866_ (.A1(net984),
    .A2(_04643_),
    .A3(_04644_),
    .B1(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__mux2_1 _09867_ (.A0(_04440_),
    .A1(_04649_),
    .S(net1187),
    .X(_04650_));
 sky130_fd_sc_hd__a22o_1 _09868_ (.A1(net2578),
    .A2(net877),
    .B1(_04650_),
    .B2(net847),
    .X(_00696_));
 sky130_fd_sc_hd__nand2_1 _09869_ (.A(net1128),
    .B(_04441_),
    .Y(_04651_));
 sky130_fd_sc_hd__inv_2 _09870_ (.A(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__or2_1 _09871_ (.A(net1128),
    .B(_04441_),
    .X(_04653_));
 sky130_fd_sc_hd__and2_1 _09872_ (.A(_04651_),
    .B(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__or3_1 _09873_ (.A(_04638_),
    .B(_04644_),
    .C(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__o21ai_1 _09874_ (.A1(_04638_),
    .A2(_04644_),
    .B1(_04654_),
    .Y(_04656_));
 sky130_fd_sc_hd__nand2b_1 _09875_ (.A_N(_04645_),
    .B(_04441_),
    .Y(_04657_));
 sky130_fd_sc_hd__o22ai_1 _09876_ (.A1(_04441_),
    .A2(_04646_),
    .B1(_04657_),
    .B2(_04623_),
    .Y(_04658_));
 sky130_fd_sc_hd__o21ai_1 _09877_ (.A1(net1146),
    .A2(_04658_),
    .B1(net1182),
    .Y(_04659_));
 sky130_fd_sc_hd__a31o_1 _09878_ (.A1(net1146),
    .A2(_04655_),
    .A3(_04656_),
    .B1(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__or2_1 _09879_ (.A(net1184),
    .B(_04441_),
    .X(_04661_));
 sky130_fd_sc_hd__a32o_1 _09880_ (.A1(net851),
    .A2(_04660_),
    .A3(_04661_),
    .B1(net881),
    .B2(net2296),
    .X(_00697_));
 sky130_fd_sc_hd__and2_1 _09881_ (.A(net1127),
    .B(_04442_),
    .X(_04662_));
 sky130_fd_sc_hd__nor2_1 _09882_ (.A(net1127),
    .B(_04442_),
    .Y(_04663_));
 sky130_fd_sc_hd__nor2_1 _09883_ (.A(_04662_),
    .B(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__and3b_1 _09884_ (.A_N(_04630_),
    .B(_04640_),
    .C(_04654_),
    .X(_04665_));
 sky130_fd_sc_hd__a41o_1 _09885_ (.A1(_04629_),
    .A2(_04640_),
    .A3(_04641_),
    .A4(_04654_),
    .B1(_04652_),
    .X(_04666_));
 sky130_fd_sc_hd__a21o_1 _09886_ (.A1(_04638_),
    .A2(_04653_),
    .B1(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__a21o_1 _09887_ (.A1(_04621_),
    .A2(_04665_),
    .B1(_04667_),
    .X(_04668_));
 sky130_fd_sc_hd__nand2_1 _09888_ (.A(_04664_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__or2_1 _09889_ (.A(_04664_),
    .B(_04668_),
    .X(_04670_));
 sky130_fd_sc_hd__a21oi_1 _09890_ (.A1(_04441_),
    .A2(_04646_),
    .B1(_04442_),
    .Y(_04671_));
 sky130_fd_sc_hd__and4b_1 _09891_ (.A_N(_04657_),
    .B(_04442_),
    .C(_04438_),
    .D(_04611_),
    .X(_04672_));
 sky130_fd_sc_hd__and3_1 _09892_ (.A(_04441_),
    .B(_04442_),
    .C(_04646_),
    .X(_04673_));
 sky130_fd_sc_hd__o31ai_1 _09893_ (.A1(net1147),
    .A2(_04671_),
    .A3(_04673_),
    .B1(net1184),
    .Y(_04674_));
 sky130_fd_sc_hd__a31o_1 _09894_ (.A1(net1147),
    .A2(_04669_),
    .A3(_04670_),
    .B1(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__or2_1 _09895_ (.A(net1184),
    .B(_04442_),
    .X(_04676_));
 sky130_fd_sc_hd__a32o_1 _09896_ (.A1(net851),
    .A2(_04675_),
    .A3(_04676_),
    .B1(net881),
    .B2(net2565),
    .X(_00698_));
 sky130_fd_sc_hd__xor2_1 _09897_ (.A(net1127),
    .B(_04443_),
    .X(_04677_));
 sky130_fd_sc_hd__a21oi_1 _09898_ (.A1(_04664_),
    .A2(_04668_),
    .B1(_04662_),
    .Y(_04678_));
 sky130_fd_sc_hd__xnor2_1 _09899_ (.A(_04677_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__or2_1 _09900_ (.A(_04443_),
    .B(_04672_),
    .X(_04680_));
 sky130_fd_sc_hd__a21oi_1 _09901_ (.A1(_04443_),
    .A2(_04673_),
    .B1(net1150),
    .Y(_04681_));
 sky130_fd_sc_hd__a22o_1 _09902_ (.A1(net1150),
    .A2(_04679_),
    .B1(_04680_),
    .B2(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__mux2_1 _09903_ (.A0(_04443_),
    .A1(_04682_),
    .S(net1184),
    .X(_04683_));
 sky130_fd_sc_hd__a22o_1 _09904_ (.A1(net2564),
    .A2(net881),
    .B1(_04683_),
    .B2(net851),
    .X(_00699_));
 sky130_fd_sc_hd__and2_1 _09905_ (.A(net1128),
    .B(_04444_),
    .X(_04684_));
 sky130_fd_sc_hd__nor2_1 _09906_ (.A(net1127),
    .B(_04444_),
    .Y(_04685_));
 sky130_fd_sc_hd__nor2_1 _09907_ (.A(_04684_),
    .B(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__o21a_1 _09908_ (.A1(_04442_),
    .A2(_04443_),
    .B1(net1127),
    .X(_04687_));
 sky130_fd_sc_hd__a31o_1 _09909_ (.A1(_04664_),
    .A2(_04668_),
    .A3(_04677_),
    .B1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__xnor2_1 _09910_ (.A(_04686_),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__a21oi_1 _09911_ (.A1(_04443_),
    .A2(_04672_),
    .B1(_04444_),
    .Y(_04690_));
 sky130_fd_sc_hd__and3_1 _09912_ (.A(_04443_),
    .B(_04444_),
    .C(_04672_),
    .X(_04691_));
 sky130_fd_sc_hd__o31a_1 _09913_ (.A1(net1150),
    .A2(_04690_),
    .A3(_04691_),
    .B1(net1184),
    .X(_04692_));
 sky130_fd_sc_hd__o21ai_1 _09914_ (.A1(net984),
    .A2(_04689_),
    .B1(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__or2_1 _09915_ (.A(net1184),
    .B(_04444_),
    .X(_04694_));
 sky130_fd_sc_hd__a32o_1 _09916_ (.A1(net851),
    .A2(_04693_),
    .A3(_04694_),
    .B1(net881),
    .B2(net2487),
    .X(_00700_));
 sky130_fd_sc_hd__xor2_1 _09917_ (.A(net1127),
    .B(_04445_),
    .X(_04695_));
 sky130_fd_sc_hd__a21o_1 _09918_ (.A1(_04686_),
    .A2(_04688_),
    .B1(_04684_),
    .X(_04696_));
 sky130_fd_sc_hd__xnor2_1 _09919_ (.A(_04695_),
    .B(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__nor2_1 _09920_ (.A(_04445_),
    .B(_04691_),
    .Y(_04698_));
 sky130_fd_sc_hd__and4_1 _09921_ (.A(_04443_),
    .B(_04444_),
    .C(_04445_),
    .D(_04673_),
    .X(_04699_));
 sky130_fd_sc_hd__o31a_1 _09922_ (.A1(net1150),
    .A2(_04698_),
    .A3(_04699_),
    .B1(net1184),
    .X(_04700_));
 sky130_fd_sc_hd__o21ai_1 _09923_ (.A1(net985),
    .A2(_04697_),
    .B1(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__or2_1 _09924_ (.A(net1184),
    .B(_04445_),
    .X(_04702_));
 sky130_fd_sc_hd__a32o_1 _09925_ (.A1(net851),
    .A2(_04701_),
    .A3(_04702_),
    .B1(net881),
    .B2(net2910),
    .X(_00701_));
 sky130_fd_sc_hd__and4_1 _09926_ (.A(_04664_),
    .B(_04677_),
    .C(_04686_),
    .D(_04695_),
    .X(_04703_));
 sky130_fd_sc_hd__o21a_1 _09927_ (.A1(_04444_),
    .A2(_04445_),
    .B1(net1127),
    .X(_04704_));
 sky130_fd_sc_hd__a211o_1 _09928_ (.A1(_04668_),
    .A2(_04703_),
    .B1(_04704_),
    .C1(_04687_),
    .X(_04705_));
 sky130_fd_sc_hd__and2_1 _09929_ (.A(net1127),
    .B(_04446_),
    .X(_04706_));
 sky130_fd_sc_hd__nor2_1 _09930_ (.A(net1127),
    .B(_04446_),
    .Y(_04707_));
 sky130_fd_sc_hd__nor2_1 _09931_ (.A(_04706_),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__xnor2_1 _09932_ (.A(_04705_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__nand2_1 _09933_ (.A(_02480_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__or2_1 _09934_ (.A(_04446_),
    .B(_04699_),
    .X(_04711_));
 sky130_fd_sc_hd__nand3_1 _09935_ (.A(_04445_),
    .B(_04446_),
    .C(_04691_),
    .Y(_04712_));
 sky130_fd_sc_hd__a21o_1 _09936_ (.A1(_04711_),
    .A2(_04712_),
    .B1(_02489_),
    .X(_04713_));
 sky130_fd_sc_hd__o211a_1 _09937_ (.A1(net1185),
    .A2(_04446_),
    .B1(_04713_),
    .C1(net849),
    .X(_04714_));
 sky130_fd_sc_hd__a22o_1 _09938_ (.A1(net3017),
    .A2(net879),
    .B1(_04710_),
    .B2(_04714_),
    .X(_00702_));
 sky130_fd_sc_hd__xor2_1 _09939_ (.A(net1127),
    .B(_04447_),
    .X(_04715_));
 sky130_fd_sc_hd__a21oi_1 _09940_ (.A1(_04705_),
    .A2(_04708_),
    .B1(_04706_),
    .Y(_04716_));
 sky130_fd_sc_hd__xnor2_1 _09941_ (.A(_04715_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__a31o_1 _09942_ (.A1(_04445_),
    .A2(_04446_),
    .A3(_04691_),
    .B1(_04447_),
    .X(_04718_));
 sky130_fd_sc_hd__and3_1 _09943_ (.A(_04446_),
    .B(_04447_),
    .C(_04699_),
    .X(_04719_));
 sky130_fd_sc_hd__nor2_1 _09944_ (.A(net1150),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__a22o_1 _09945_ (.A1(net1150),
    .A2(_04717_),
    .B1(_04718_),
    .B2(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__mux2_1 _09946_ (.A0(_04447_),
    .A1(_04721_),
    .S(net1185),
    .X(_04722_));
 sky130_fd_sc_hd__a22o_1 _09947_ (.A1(net2644),
    .A2(net879),
    .B1(_04722_),
    .B2(net849),
    .X(_00703_));
 sky130_fd_sc_hd__xor2_1 _09948_ (.A(net1129),
    .B(_04448_),
    .X(_04723_));
 sky130_fd_sc_hd__o21a_1 _09949_ (.A1(_04446_),
    .A2(_04447_),
    .B1(net1129),
    .X(_04724_));
 sky130_fd_sc_hd__and3_1 _09950_ (.A(_04705_),
    .B(_04708_),
    .C(_04715_),
    .X(_04725_));
 sky130_fd_sc_hd__o21a_1 _09951_ (.A1(_04724_),
    .A2(_04725_),
    .B1(_04723_),
    .X(_04726_));
 sky130_fd_sc_hd__o31ai_1 _09952_ (.A1(_04723_),
    .A2(_04724_),
    .A3(_04725_),
    .B1(net1150),
    .Y(_04727_));
 sky130_fd_sc_hd__nand2_1 _09953_ (.A(_04448_),
    .B(_04719_),
    .Y(_04728_));
 sky130_fd_sc_hd__o21a_1 _09954_ (.A1(_04448_),
    .A2(_04719_),
    .B1(net985),
    .X(_04729_));
 sky130_fd_sc_hd__a2bb2o_1 _09955_ (.A1_N(_04726_),
    .A2_N(_04727_),
    .B1(_04728_),
    .B2(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__mux2_1 _09956_ (.A0(_04448_),
    .A1(_04730_),
    .S(net1185),
    .X(_04731_));
 sky130_fd_sc_hd__a22o_1 _09957_ (.A1(net2597),
    .A2(net880),
    .B1(_04731_),
    .B2(net850),
    .X(_00704_));
 sky130_fd_sc_hd__xor2_1 _09958_ (.A(net1129),
    .B(_04449_),
    .X(_04732_));
 sky130_fd_sc_hd__a21o_1 _09959_ (.A1(net1129),
    .A2(_04448_),
    .B1(_04726_),
    .X(_04733_));
 sky130_fd_sc_hd__xnor2_1 _09960_ (.A(_04732_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__a21oi_1 _09961_ (.A1(_04448_),
    .A2(_04719_),
    .B1(_04449_),
    .Y(_04735_));
 sky130_fd_sc_hd__and3_1 _09962_ (.A(_04448_),
    .B(_04449_),
    .C(_04719_),
    .X(_04736_));
 sky130_fd_sc_hd__or3_1 _09963_ (.A(net1150),
    .B(_04735_),
    .C(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__o211a_1 _09964_ (.A1(net985),
    .A2(_04734_),
    .B1(_04737_),
    .C1(net1185),
    .X(_04738_));
 sky130_fd_sc_hd__o21ai_1 _09965_ (.A1(net1185),
    .A2(_04449_),
    .B1(net849),
    .Y(_04739_));
 sky130_fd_sc_hd__a2bb2o_1 _09966_ (.A1_N(_04738_),
    .A2_N(_04739_),
    .B1(net2639),
    .B2(net879),
    .X(_00705_));
 sky130_fd_sc_hd__o21a_1 _09967_ (.A1(_04448_),
    .A2(_04449_),
    .B1(net1129),
    .X(_04740_));
 sky130_fd_sc_hd__a311o_1 _09968_ (.A1(_04723_),
    .A2(_04725_),
    .A3(_04732_),
    .B1(_04740_),
    .C1(_04724_),
    .X(_04741_));
 sky130_fd_sc_hd__and2_1 _09969_ (.A(net1129),
    .B(_04450_),
    .X(_04742_));
 sky130_fd_sc_hd__nor2_1 _09970_ (.A(net1129),
    .B(_04450_),
    .Y(_04743_));
 sky130_fd_sc_hd__nor2_1 _09971_ (.A(_04742_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__o21ai_1 _09972_ (.A1(_04741_),
    .A2(_04744_),
    .B1(net1152),
    .Y(_04745_));
 sky130_fd_sc_hd__a21o_1 _09973_ (.A1(_04741_),
    .A2(_04744_),
    .B1(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__nor2_1 _09974_ (.A(_04450_),
    .B(_04736_),
    .Y(_04747_));
 sky130_fd_sc_hd__and2_1 _09975_ (.A(_04450_),
    .B(_04736_),
    .X(_04748_));
 sky130_fd_sc_hd__o311a_1 _09976_ (.A1(net1152),
    .A2(_04747_),
    .A3(_04748_),
    .B1(_04746_),
    .C1(net1185),
    .X(_04749_));
 sky130_fd_sc_hd__o21ai_1 _09977_ (.A1(net1185),
    .A2(_04450_),
    .B1(net849),
    .Y(_04750_));
 sky130_fd_sc_hd__a2bb2o_1 _09978_ (.A1_N(_04749_),
    .A2_N(_04750_),
    .B1(net2586),
    .B2(net879),
    .X(_00706_));
 sky130_fd_sc_hd__a21o_1 _09979_ (.A1(_04741_),
    .A2(_04744_),
    .B1(_04742_),
    .X(_04751_));
 sky130_fd_sc_hd__nand2_1 _09980_ (.A(net1129),
    .B(_04451_),
    .Y(_04752_));
 sky130_fd_sc_hd__or2_1 _09981_ (.A(net1129),
    .B(_04451_),
    .X(_04753_));
 sky130_fd_sc_hd__nand2_1 _09982_ (.A(_04752_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__xnor2_1 _09983_ (.A(_04751_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _09984_ (.A(net1152),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__nor2_1 _09985_ (.A(_04451_),
    .B(_04748_),
    .Y(_04757_));
 sky130_fd_sc_hd__and3_1 _09986_ (.A(_04450_),
    .B(_04451_),
    .C(_04736_),
    .X(_04758_));
 sky130_fd_sc_hd__o31a_1 _09987_ (.A1(net1152),
    .A2(_04757_),
    .A3(_04758_),
    .B1(net1186),
    .X(_04759_));
 sky130_fd_sc_hd__o2bb2a_1 _09988_ (.A1_N(_04756_),
    .A2_N(_04759_),
    .B1(net1186),
    .B2(_04451_),
    .X(_04760_));
 sky130_fd_sc_hd__a22o_1 _09989_ (.A1(net2607),
    .A2(net879),
    .B1(_04760_),
    .B2(net849),
    .X(_00707_));
 sky130_fd_sc_hd__a21bo_1 _09990_ (.A1(_04751_),
    .A2(_04753_),
    .B1_N(_04752_),
    .X(_04761_));
 sky130_fd_sc_hd__xnor2_1 _09991_ (.A(net1129),
    .B(_04452_),
    .Y(_04762_));
 sky130_fd_sc_hd__xnor2_1 _09992_ (.A(_04452_),
    .B(_04758_),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2_1 _09993_ (.A(net1152),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__xnor2_1 _09994_ (.A(_04761_),
    .B(_04762_),
    .Y(_04765_));
 sky130_fd_sc_hd__a211o_1 _09995_ (.A1(net1152),
    .A2(_04765_),
    .B1(_04764_),
    .C1(_02380_),
    .X(_04766_));
 sky130_fd_sc_hd__or2_1 _09996_ (.A(net1185),
    .B(_04452_),
    .X(_04767_));
 sky130_fd_sc_hd__a32o_1 _09997_ (.A1(net849),
    .A2(_04766_),
    .A3(_04767_),
    .B1(net879),
    .B2(net2512),
    .X(_00708_));
 sky130_fd_sc_hd__nor2_1 _09998_ (.A(net1206),
    .B(net2605),
    .Y(_00709_));
 sky130_fd_sc_hd__o21ai_1 _09999_ (.A1(\count_cycle[0] ),
    .A2(\count_cycle[1] ),
    .B1(net1231),
    .Y(_04768_));
 sky130_fd_sc_hd__a21oi_1 _10000_ (.A1(net2605),
    .A2(net2906),
    .B1(_04768_),
    .Y(_00710_));
 sky130_fd_sc_hd__a21o_1 _10001_ (.A1(\count_cycle[0] ),
    .A2(\count_cycle[1] ),
    .B1(\count_cycle[2] ),
    .X(_04769_));
 sky130_fd_sc_hd__and3_1 _10002_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .X(_04770_));
 sky130_fd_sc_hd__and3b_1 _10003_ (.A_N(_04770_),
    .B(net1231),
    .C(_04769_),
    .X(_00711_));
 sky130_fd_sc_hd__and4_1 _10004_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .C(\count_cycle[2] ),
    .D(\count_cycle[3] ),
    .X(_04771_));
 sky130_fd_sc_hd__o21ai_1 _10005_ (.A1(net2857),
    .A2(_04770_),
    .B1(net1231),
    .Y(_04772_));
 sky130_fd_sc_hd__nor2_1 _10006_ (.A(_04771_),
    .B(_04772_),
    .Y(_00712_));
 sky130_fd_sc_hd__a21oi_1 _10007_ (.A1(\count_cycle[4] ),
    .A2(_04771_),
    .B1(net1205),
    .Y(_04773_));
 sky130_fd_sc_hd__o21a_1 _10008_ (.A1(net3039),
    .A2(_04771_),
    .B1(_04773_),
    .X(_00713_));
 sky130_fd_sc_hd__a21o_1 _10009_ (.A1(\count_cycle[4] ),
    .A2(_04771_),
    .B1(\count_cycle[5] ),
    .X(_04774_));
 sky130_fd_sc_hd__and3_1 _10010_ (.A(\count_cycle[4] ),
    .B(\count_cycle[5] ),
    .C(_04771_),
    .X(_04775_));
 sky130_fd_sc_hd__and3b_1 _10011_ (.A_N(_04775_),
    .B(net1223),
    .C(_04774_),
    .X(_00714_));
 sky130_fd_sc_hd__and4_1 _10012_ (.A(\count_cycle[4] ),
    .B(\count_cycle[5] ),
    .C(\count_cycle[6] ),
    .D(_04771_),
    .X(_04776_));
 sky130_fd_sc_hd__o21ai_1 _10013_ (.A1(net2848),
    .A2(_04775_),
    .B1(net1223),
    .Y(_04777_));
 sky130_fd_sc_hd__nor2_1 _10014_ (.A(_04776_),
    .B(_04777_),
    .Y(_00715_));
 sky130_fd_sc_hd__a21oi_1 _10015_ (.A1(\count_cycle[7] ),
    .A2(_04776_),
    .B1(net1204),
    .Y(_04778_));
 sky130_fd_sc_hd__o21a_1 _10016_ (.A1(\count_cycle[7] ),
    .A2(_04776_),
    .B1(_04778_),
    .X(_00716_));
 sky130_fd_sc_hd__a21o_1 _10017_ (.A1(\count_cycle[7] ),
    .A2(_04776_),
    .B1(\count_cycle[8] ),
    .X(_04779_));
 sky130_fd_sc_hd__and3_1 _10018_ (.A(\count_cycle[7] ),
    .B(\count_cycle[8] ),
    .C(_04776_),
    .X(_04780_));
 sky130_fd_sc_hd__and3b_1 _10019_ (.A_N(_04780_),
    .B(net1223),
    .C(_04779_),
    .X(_00717_));
 sky130_fd_sc_hd__and4_1 _10020_ (.A(\count_cycle[7] ),
    .B(\count_cycle[8] ),
    .C(\count_cycle[9] ),
    .D(_04776_),
    .X(_04781_));
 sky130_fd_sc_hd__o21ai_1 _10021_ (.A1(net2790),
    .A2(_04780_),
    .B1(net1223),
    .Y(_04782_));
 sky130_fd_sc_hd__nor2_1 _10022_ (.A(_04781_),
    .B(_04782_),
    .Y(_00718_));
 sky130_fd_sc_hd__a21oi_1 _10023_ (.A1(\count_cycle[10] ),
    .A2(_04781_),
    .B1(net1205),
    .Y(_04783_));
 sky130_fd_sc_hd__o21a_1 _10024_ (.A1(net3054),
    .A2(_04781_),
    .B1(_04783_),
    .X(_00719_));
 sky130_fd_sc_hd__a21o_1 _10025_ (.A1(\count_cycle[10] ),
    .A2(_04781_),
    .B1(\count_cycle[11] ),
    .X(_04784_));
 sky130_fd_sc_hd__and3_1 _10026_ (.A(\count_cycle[10] ),
    .B(\count_cycle[11] ),
    .C(_04781_),
    .X(_04785_));
 sky130_fd_sc_hd__and3b_1 _10027_ (.A_N(_04785_),
    .B(net1224),
    .C(_04784_),
    .X(_00720_));
 sky130_fd_sc_hd__and4_1 _10028_ (.A(\count_cycle[10] ),
    .B(\count_cycle[11] ),
    .C(\count_cycle[12] ),
    .D(_04781_),
    .X(_04786_));
 sky130_fd_sc_hd__o21ai_1 _10029_ (.A1(net2784),
    .A2(_04785_),
    .B1(net1224),
    .Y(_04787_));
 sky130_fd_sc_hd__nor2_1 _10030_ (.A(_04786_),
    .B(_04787_),
    .Y(_00721_));
 sky130_fd_sc_hd__a21oi_1 _10031_ (.A1(\count_cycle[13] ),
    .A2(_04786_),
    .B1(net1191),
    .Y(_04788_));
 sky130_fd_sc_hd__o21a_1 _10032_ (.A1(net3041),
    .A2(_04786_),
    .B1(_04788_),
    .X(_00722_));
 sky130_fd_sc_hd__a21o_1 _10033_ (.A1(\count_cycle[13] ),
    .A2(_04786_),
    .B1(\count_cycle[14] ),
    .X(_04789_));
 sky130_fd_sc_hd__and3_1 _10034_ (.A(\count_cycle[13] ),
    .B(\count_cycle[14] ),
    .C(_04786_),
    .X(_04790_));
 sky130_fd_sc_hd__and3b_1 _10035_ (.A_N(_04790_),
    .B(net1224),
    .C(_04789_),
    .X(_00723_));
 sky130_fd_sc_hd__and4_2 _10036_ (.A(\count_cycle[13] ),
    .B(\count_cycle[14] ),
    .C(\count_cycle[15] ),
    .D(_04786_),
    .X(_04791_));
 sky130_fd_sc_hd__o21ai_1 _10037_ (.A1(net2720),
    .A2(_04790_),
    .B1(net1224),
    .Y(_04792_));
 sky130_fd_sc_hd__nor2_1 _10038_ (.A(_04791_),
    .B(_04792_),
    .Y(_00724_));
 sky130_fd_sc_hd__a21oi_1 _10039_ (.A1(\count_cycle[16] ),
    .A2(_04791_),
    .B1(net1206),
    .Y(_04793_));
 sky130_fd_sc_hd__o21a_1 _10040_ (.A1(net2988),
    .A2(_04791_),
    .B1(_04793_),
    .X(_00725_));
 sky130_fd_sc_hd__a21oi_1 _10041_ (.A1(\count_cycle[16] ),
    .A2(_04791_),
    .B1(net2787),
    .Y(_04794_));
 sky130_fd_sc_hd__and2_1 _10042_ (.A(\count_cycle[16] ),
    .B(\count_cycle[17] ),
    .X(_04795_));
 sky130_fd_sc_hd__a211oi_1 _10043_ (.A1(_04791_),
    .A2(_04795_),
    .B1(_04794_),
    .C1(net1206),
    .Y(_00726_));
 sky130_fd_sc_hd__a21o_1 _10044_ (.A1(_04791_),
    .A2(_04795_),
    .B1(\count_cycle[18] ),
    .X(_04796_));
 sky130_fd_sc_hd__and3_1 _10045_ (.A(\count_cycle[18] ),
    .B(_04791_),
    .C(_04795_),
    .X(_04797_));
 sky130_fd_sc_hd__and3b_1 _10046_ (.A_N(_04797_),
    .B(net1229),
    .C(_04796_),
    .X(_00727_));
 sky130_fd_sc_hd__and4_1 _10047_ (.A(\count_cycle[18] ),
    .B(\count_cycle[19] ),
    .C(_04791_),
    .D(_04795_),
    .X(_04798_));
 sky130_fd_sc_hd__o21ai_1 _10048_ (.A1(net2885),
    .A2(_04797_),
    .B1(net1229),
    .Y(_04799_));
 sky130_fd_sc_hd__nor2_1 _10049_ (.A(_04798_),
    .B(_04799_),
    .Y(_00728_));
 sky130_fd_sc_hd__and2_1 _10050_ (.A(\count_cycle[20] ),
    .B(_04798_),
    .X(_04800_));
 sky130_fd_sc_hd__o21ai_1 _10051_ (.A1(\count_cycle[20] ),
    .A2(_04798_),
    .B1(net1235),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _10052_ (.A(_04800_),
    .B(_04801_),
    .Y(_00729_));
 sky130_fd_sc_hd__and3_1 _10053_ (.A(\count_cycle[20] ),
    .B(\count_cycle[21] ),
    .C(_04798_),
    .X(_04802_));
 sky130_fd_sc_hd__o21ai_1 _10054_ (.A1(net2972),
    .A2(_04800_),
    .B1(net1235),
    .Y(_04803_));
 sky130_fd_sc_hd__nor2_1 _10055_ (.A(_04802_),
    .B(_04803_),
    .Y(_00730_));
 sky130_fd_sc_hd__and4_1 _10056_ (.A(\count_cycle[20] ),
    .B(\count_cycle[21] ),
    .C(\count_cycle[22] ),
    .D(_04798_),
    .X(_04804_));
 sky130_fd_sc_hd__o21ai_1 _10057_ (.A1(net2851),
    .A2(_04802_),
    .B1(net1235),
    .Y(_04805_));
 sky130_fd_sc_hd__nor2_1 _10058_ (.A(_04804_),
    .B(_04805_),
    .Y(_00731_));
 sky130_fd_sc_hd__and2_1 _10059_ (.A(\count_cycle[23] ),
    .B(_04804_),
    .X(_04806_));
 sky130_fd_sc_hd__o21ai_1 _10060_ (.A1(net3038),
    .A2(_04804_),
    .B1(net1236),
    .Y(_04807_));
 sky130_fd_sc_hd__nor2_1 _10061_ (.A(_04806_),
    .B(_04807_),
    .Y(_00732_));
 sky130_fd_sc_hd__and3_1 _10062_ (.A(\count_cycle[23] ),
    .B(\count_cycle[24] ),
    .C(_04804_),
    .X(_04808_));
 sky130_fd_sc_hd__o21ai_1 _10063_ (.A1(net2996),
    .A2(_04806_),
    .B1(net1236),
    .Y(_04809_));
 sky130_fd_sc_hd__nor2_1 _10064_ (.A(_04808_),
    .B(_04809_),
    .Y(_00733_));
 sky130_fd_sc_hd__or2_1 _10065_ (.A(\count_cycle[25] ),
    .B(_04808_),
    .X(_04810_));
 sky130_fd_sc_hd__and4_1 _10066_ (.A(\count_cycle[23] ),
    .B(\count_cycle[24] ),
    .C(\count_cycle[25] ),
    .D(_04804_),
    .X(_04811_));
 sky130_fd_sc_hd__and3b_1 _10067_ (.A_N(_04811_),
    .B(net1236),
    .C(_04810_),
    .X(_00734_));
 sky130_fd_sc_hd__or2_1 _10068_ (.A(\count_cycle[26] ),
    .B(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__and2_1 _10069_ (.A(\count_cycle[26] ),
    .B(_04811_),
    .X(_04813_));
 sky130_fd_sc_hd__and3b_1 _10070_ (.A_N(_04813_),
    .B(net1236),
    .C(_04812_),
    .X(_00735_));
 sky130_fd_sc_hd__and3_1 _10071_ (.A(\count_cycle[26] ),
    .B(\count_cycle[27] ),
    .C(_04811_),
    .X(_04814_));
 sky130_fd_sc_hd__o21ai_1 _10072_ (.A1(net2987),
    .A2(_04813_),
    .B1(net1236),
    .Y(_04815_));
 sky130_fd_sc_hd__nor2_1 _10073_ (.A(_04814_),
    .B(_04815_),
    .Y(_00736_));
 sky130_fd_sc_hd__and4_1 _10074_ (.A(\count_cycle[26] ),
    .B(\count_cycle[27] ),
    .C(\count_cycle[28] ),
    .D(_04811_),
    .X(_04816_));
 sky130_fd_sc_hd__o21ai_1 _10075_ (.A1(net2747),
    .A2(_04814_),
    .B1(net1236),
    .Y(_04817_));
 sky130_fd_sc_hd__nor2_1 _10076_ (.A(_04816_),
    .B(_04817_),
    .Y(_00737_));
 sky130_fd_sc_hd__a21oi_1 _10077_ (.A1(\count_cycle[29] ),
    .A2(_04816_),
    .B1(net1209),
    .Y(_04818_));
 sky130_fd_sc_hd__o21a_1 _10078_ (.A1(\count_cycle[29] ),
    .A2(_04816_),
    .B1(_04818_),
    .X(_00738_));
 sky130_fd_sc_hd__a21o_1 _10079_ (.A1(\count_cycle[29] ),
    .A2(_04816_),
    .B1(\count_cycle[30] ),
    .X(_04819_));
 sky130_fd_sc_hd__and3_1 _10080_ (.A(\count_cycle[29] ),
    .B(\count_cycle[30] ),
    .C(_04816_),
    .X(_04820_));
 sky130_fd_sc_hd__and3b_1 _10081_ (.A_N(_04820_),
    .B(net1235),
    .C(_04819_),
    .X(_00739_));
 sky130_fd_sc_hd__and4_2 _10082_ (.A(\count_cycle[29] ),
    .B(\count_cycle[30] ),
    .C(\count_cycle[31] ),
    .D(_04816_),
    .X(_04821_));
 sky130_fd_sc_hd__o21ai_1 _10083_ (.A1(net2788),
    .A2(_04820_),
    .B1(net1235),
    .Y(_04822_));
 sky130_fd_sc_hd__nor2_1 _10084_ (.A(_04821_),
    .B(_04822_),
    .Y(_00740_));
 sky130_fd_sc_hd__a21oi_1 _10085_ (.A1(\count_cycle[32] ),
    .A2(_04821_),
    .B1(net1207),
    .Y(_04823_));
 sky130_fd_sc_hd__o21a_1 _10086_ (.A1(net3062),
    .A2(_04821_),
    .B1(_04823_),
    .X(_00741_));
 sky130_fd_sc_hd__a21o_1 _10087_ (.A1(\count_cycle[32] ),
    .A2(_04821_),
    .B1(\count_cycle[33] ),
    .X(_04824_));
 sky130_fd_sc_hd__and3_1 _10088_ (.A(\count_cycle[32] ),
    .B(\count_cycle[33] ),
    .C(_04821_),
    .X(_04825_));
 sky130_fd_sc_hd__and3b_1 _10089_ (.A_N(_04825_),
    .B(net1228),
    .C(_04824_),
    .X(_00742_));
 sky130_fd_sc_hd__and4_2 _10090_ (.A(\count_cycle[32] ),
    .B(\count_cycle[33] ),
    .C(\count_cycle[34] ),
    .D(_04821_),
    .X(_04826_));
 sky130_fd_sc_hd__o21ai_1 _10091_ (.A1(net2940),
    .A2(_04825_),
    .B1(net1228),
    .Y(_04827_));
 sky130_fd_sc_hd__nor2_1 _10092_ (.A(_04826_),
    .B(_04827_),
    .Y(_00743_));
 sky130_fd_sc_hd__a21oi_1 _10093_ (.A1(\count_cycle[35] ),
    .A2(_04826_),
    .B1(net1206),
    .Y(_04828_));
 sky130_fd_sc_hd__o21a_1 _10094_ (.A1(net3030),
    .A2(_04826_),
    .B1(_04828_),
    .X(_00744_));
 sky130_fd_sc_hd__a21o_1 _10095_ (.A1(\count_cycle[35] ),
    .A2(_04826_),
    .B1(\count_cycle[36] ),
    .X(_04829_));
 sky130_fd_sc_hd__and3_1 _10096_ (.A(\count_cycle[35] ),
    .B(\count_cycle[36] ),
    .C(_04826_),
    .X(_04830_));
 sky130_fd_sc_hd__and3b_1 _10097_ (.A_N(_04830_),
    .B(net1225),
    .C(_04829_),
    .X(_00745_));
 sky130_fd_sc_hd__and4_1 _10098_ (.A(\count_cycle[35] ),
    .B(\count_cycle[36] ),
    .C(\count_cycle[37] ),
    .D(_04826_),
    .X(_04831_));
 sky130_fd_sc_hd__o21ai_1 _10099_ (.A1(net2745),
    .A2(_04830_),
    .B1(net1225),
    .Y(_04832_));
 sky130_fd_sc_hd__nor2_1 _10100_ (.A(_04831_),
    .B(_04832_),
    .Y(_00746_));
 sky130_fd_sc_hd__a21oi_1 _10101_ (.A1(\count_cycle[38] ),
    .A2(_04831_),
    .B1(net1206),
    .Y(_04833_));
 sky130_fd_sc_hd__o21a_1 _10102_ (.A1(\count_cycle[38] ),
    .A2(_04831_),
    .B1(_04833_),
    .X(_00747_));
 sky130_fd_sc_hd__a21o_1 _10103_ (.A1(\count_cycle[38] ),
    .A2(_04831_),
    .B1(\count_cycle[39] ),
    .X(_04834_));
 sky130_fd_sc_hd__and3_1 _10104_ (.A(\count_cycle[38] ),
    .B(\count_cycle[39] ),
    .C(_04831_),
    .X(_04835_));
 sky130_fd_sc_hd__and3b_1 _10105_ (.A_N(_04835_),
    .B(net1225),
    .C(_04834_),
    .X(_00748_));
 sky130_fd_sc_hd__and4_1 _10106_ (.A(\count_cycle[38] ),
    .B(\count_cycle[39] ),
    .C(\count_cycle[40] ),
    .D(_04831_),
    .X(_04836_));
 sky130_fd_sc_hd__o21ai_1 _10107_ (.A1(net2841),
    .A2(_04835_),
    .B1(net1225),
    .Y(_04837_));
 sky130_fd_sc_hd__nor2_1 _10108_ (.A(_04836_),
    .B(_04837_),
    .Y(_00749_));
 sky130_fd_sc_hd__a21oi_1 _10109_ (.A1(\count_cycle[41] ),
    .A2(_04836_),
    .B1(net1204),
    .Y(_04838_));
 sky130_fd_sc_hd__o21a_1 _10110_ (.A1(net3067),
    .A2(_04836_),
    .B1(_04838_),
    .X(_00750_));
 sky130_fd_sc_hd__a21o_1 _10111_ (.A1(\count_cycle[41] ),
    .A2(_04836_),
    .B1(\count_cycle[42] ),
    .X(_04839_));
 sky130_fd_sc_hd__and3_1 _10112_ (.A(\count_cycle[41] ),
    .B(\count_cycle[42] ),
    .C(_04836_),
    .X(_04840_));
 sky130_fd_sc_hd__and3b_1 _10113_ (.A_N(_04840_),
    .B(net1225),
    .C(_04839_),
    .X(_00751_));
 sky130_fd_sc_hd__and4_2 _10114_ (.A(\count_cycle[41] ),
    .B(\count_cycle[42] ),
    .C(\count_cycle[43] ),
    .D(_04836_),
    .X(_04841_));
 sky130_fd_sc_hd__o21ai_1 _10115_ (.A1(net2860),
    .A2(_04840_),
    .B1(net1225),
    .Y(_04842_));
 sky130_fd_sc_hd__nor2_1 _10116_ (.A(_04841_),
    .B(_04842_),
    .Y(_00752_));
 sky130_fd_sc_hd__a21oi_1 _10117_ (.A1(\count_cycle[44] ),
    .A2(_04841_),
    .B1(net1206),
    .Y(_04843_));
 sky130_fd_sc_hd__o21a_1 _10118_ (.A1(\count_cycle[44] ),
    .A2(_04841_),
    .B1(_04843_),
    .X(_00753_));
 sky130_fd_sc_hd__a21o_1 _10119_ (.A1(\count_cycle[44] ),
    .A2(_04841_),
    .B1(\count_cycle[45] ),
    .X(_04844_));
 sky130_fd_sc_hd__and3_1 _10120_ (.A(\count_cycle[44] ),
    .B(\count_cycle[45] ),
    .C(_04841_),
    .X(_04845_));
 sky130_fd_sc_hd__and3b_1 _10121_ (.A_N(_04845_),
    .B(net1228),
    .C(_04844_),
    .X(_00754_));
 sky130_fd_sc_hd__and4_1 _10122_ (.A(\count_cycle[44] ),
    .B(\count_cycle[45] ),
    .C(\count_cycle[46] ),
    .D(_04841_),
    .X(_04846_));
 sky130_fd_sc_hd__o21ai_1 _10123_ (.A1(net2824),
    .A2(_04845_),
    .B1(net1228),
    .Y(_04847_));
 sky130_fd_sc_hd__nor2_1 _10124_ (.A(_04846_),
    .B(_04847_),
    .Y(_00755_));
 sky130_fd_sc_hd__and2_1 _10125_ (.A(\count_cycle[47] ),
    .B(_04846_),
    .X(_04848_));
 sky130_fd_sc_hd__o21ai_1 _10126_ (.A1(\count_cycle[47] ),
    .A2(_04846_),
    .B1(net1228),
    .Y(_04849_));
 sky130_fd_sc_hd__nor2_1 _10127_ (.A(_04848_),
    .B(_04849_),
    .Y(_00756_));
 sky130_fd_sc_hd__o21ai_1 _10128_ (.A1(net2701),
    .A2(_04848_),
    .B1(net1228),
    .Y(_04850_));
 sky130_fd_sc_hd__a21oi_1 _10129_ (.A1(net2701),
    .A2(_04848_),
    .B1(_04850_),
    .Y(_00757_));
 sky130_fd_sc_hd__a31o_1 _10130_ (.A1(\count_cycle[47] ),
    .A2(\count_cycle[48] ),
    .A3(_04846_),
    .B1(\count_cycle[49] ),
    .X(_04851_));
 sky130_fd_sc_hd__and2_1 _10131_ (.A(\count_cycle[48] ),
    .B(\count_cycle[49] ),
    .X(_04852_));
 sky130_fd_sc_hd__and3_1 _10132_ (.A(\count_cycle[47] ),
    .B(_04846_),
    .C(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__and3b_1 _10133_ (.A_N(_04853_),
    .B(net1229),
    .C(_04851_),
    .X(_00758_));
 sky130_fd_sc_hd__and4_1 _10134_ (.A(\count_cycle[47] ),
    .B(\count_cycle[50] ),
    .C(_04846_),
    .D(_04852_),
    .X(_04854_));
 sky130_fd_sc_hd__o21ai_1 _10135_ (.A1(net2783),
    .A2(_04853_),
    .B1(net1229),
    .Y(_04855_));
 sky130_fd_sc_hd__nor2_1 _10136_ (.A(_04854_),
    .B(_04855_),
    .Y(_00759_));
 sky130_fd_sc_hd__and2_1 _10137_ (.A(\count_cycle[51] ),
    .B(_04854_),
    .X(_04856_));
 sky130_fd_sc_hd__o21ai_1 _10138_ (.A1(\count_cycle[51] ),
    .A2(_04854_),
    .B1(net1235),
    .Y(_04857_));
 sky130_fd_sc_hd__nor2_1 _10139_ (.A(_04856_),
    .B(_04857_),
    .Y(_00760_));
 sky130_fd_sc_hd__and3_1 _10140_ (.A(\count_cycle[51] ),
    .B(\count_cycle[52] ),
    .C(_04854_),
    .X(_04858_));
 sky130_fd_sc_hd__o21ai_1 _10141_ (.A1(net3001),
    .A2(_04856_),
    .B1(net1235),
    .Y(_04859_));
 sky130_fd_sc_hd__nor2_1 _10142_ (.A(_04858_),
    .B(_04859_),
    .Y(_00761_));
 sky130_fd_sc_hd__and4_2 _10143_ (.A(\count_cycle[51] ),
    .B(\count_cycle[52] ),
    .C(\count_cycle[53] ),
    .D(_04854_),
    .X(_04860_));
 sky130_fd_sc_hd__o21ai_1 _10144_ (.A1(net2862),
    .A2(_04858_),
    .B1(net1235),
    .Y(_04861_));
 sky130_fd_sc_hd__nor2_1 _10145_ (.A(_04860_),
    .B(_04861_),
    .Y(_00762_));
 sky130_fd_sc_hd__a21oi_1 _10146_ (.A1(\count_cycle[54] ),
    .A2(_04860_),
    .B1(net1215),
    .Y(_04862_));
 sky130_fd_sc_hd__o21a_1 _10147_ (.A1(net3045),
    .A2(_04860_),
    .B1(_04862_),
    .X(_00763_));
 sky130_fd_sc_hd__a21o_1 _10148_ (.A1(\count_cycle[54] ),
    .A2(_04860_),
    .B1(\count_cycle[55] ),
    .X(_04863_));
 sky130_fd_sc_hd__and3_1 _10149_ (.A(\count_cycle[54] ),
    .B(\count_cycle[55] ),
    .C(_04860_),
    .X(_04864_));
 sky130_fd_sc_hd__and3b_1 _10150_ (.A_N(_04864_),
    .B(net1238),
    .C(_04863_),
    .X(_00764_));
 sky130_fd_sc_hd__o21ai_1 _10151_ (.A1(\count_cycle[56] ),
    .A2(_04864_),
    .B1(net1238),
    .Y(_04865_));
 sky130_fd_sc_hd__a21oi_1 _10152_ (.A1(net2758),
    .A2(_04864_),
    .B1(_04865_),
    .Y(_00765_));
 sky130_fd_sc_hd__a21o_1 _10153_ (.A1(\count_cycle[56] ),
    .A2(_04864_),
    .B1(\count_cycle[57] ),
    .X(_04866_));
 sky130_fd_sc_hd__and2_1 _10154_ (.A(\count_cycle[56] ),
    .B(\count_cycle[57] ),
    .X(_04867_));
 sky130_fd_sc_hd__and4_1 _10155_ (.A(\count_cycle[54] ),
    .B(\count_cycle[55] ),
    .C(_04860_),
    .D(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__and3b_1 _10156_ (.A_N(_04868_),
    .B(net1238),
    .C(_04866_),
    .X(_00766_));
 sky130_fd_sc_hd__and2_1 _10157_ (.A(\count_cycle[58] ),
    .B(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__o21ai_1 _10158_ (.A1(\count_cycle[58] ),
    .A2(_04868_),
    .B1(net1239),
    .Y(_04870_));
 sky130_fd_sc_hd__nor2_1 _10159_ (.A(_04869_),
    .B(_04870_),
    .Y(_00767_));
 sky130_fd_sc_hd__and3_1 _10160_ (.A(\count_cycle[58] ),
    .B(\count_cycle[59] ),
    .C(_04868_),
    .X(_04871_));
 sky130_fd_sc_hd__o21ai_1 _10161_ (.A1(net2968),
    .A2(_04869_),
    .B1(net1238),
    .Y(_04872_));
 sky130_fd_sc_hd__nor2_1 _10162_ (.A(_04871_),
    .B(_04872_),
    .Y(_00768_));
 sky130_fd_sc_hd__and4_2 _10163_ (.A(\count_cycle[58] ),
    .B(\count_cycle[59] ),
    .C(\count_cycle[60] ),
    .D(_04868_),
    .X(_04873_));
 sky130_fd_sc_hd__o21ai_1 _10164_ (.A1(net2797),
    .A2(_04871_),
    .B1(net1238),
    .Y(_04874_));
 sky130_fd_sc_hd__nor2_1 _10165_ (.A(_04873_),
    .B(_04874_),
    .Y(_00769_));
 sky130_fd_sc_hd__a21oi_1 _10166_ (.A1(\count_cycle[61] ),
    .A2(_04873_),
    .B1(net1209),
    .Y(_04875_));
 sky130_fd_sc_hd__o21a_1 _10167_ (.A1(\count_cycle[61] ),
    .A2(_04873_),
    .B1(_04875_),
    .X(_00770_));
 sky130_fd_sc_hd__a21oi_1 _10168_ (.A1(\count_cycle[61] ),
    .A2(_04873_),
    .B1(net2991),
    .Y(_04876_));
 sky130_fd_sc_hd__a311oi_1 _10169_ (.A1(\count_cycle[61] ),
    .A2(net2991),
    .A3(_04873_),
    .B1(_04876_),
    .C1(net1209),
    .Y(_00771_));
 sky130_fd_sc_hd__a31o_1 _10170_ (.A1(\count_cycle[61] ),
    .A2(\count_cycle[62] ),
    .A3(_04873_),
    .B1(\count_cycle[63] ),
    .X(_04877_));
 sky130_fd_sc_hd__a41o_1 _10171_ (.A1(\count_cycle[61] ),
    .A2(\count_cycle[62] ),
    .A3(\count_cycle[63] ),
    .A4(_04873_),
    .B1(net1209),
    .X(_04878_));
 sky130_fd_sc_hd__and2b_1 _10172_ (.A_N(_04878_),
    .B(_04877_),
    .X(_00772_));
 sky130_fd_sc_hd__nor2_2 _10173_ (.A(net1068),
    .B(net958),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_1 _10174_ (.A(net1068),
    .B(net958),
    .X(_04880_));
 sky130_fd_sc_hd__nor2_1 _10175_ (.A(net1088),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__or3_1 _10176_ (.A(net1207),
    .B(_02478_),
    .C(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__or2_2 _10177_ (.A(instr_sra),
    .B(instr_srai),
    .X(_04883_));
 sky130_fd_sc_hd__nor3_4 _10178_ (.A(instr_srl),
    .B(instr_srli),
    .C(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__or3_1 _10179_ (.A(instr_srl),
    .B(instr_srli),
    .C(_04883_),
    .X(_04885_));
 sky130_fd_sc_hd__or4b_1 _10180_ (.A(instr_sll),
    .B(net756),
    .C(instr_slli),
    .D_N(net1068),
    .X(_04886_));
 sky130_fd_sc_hd__and4bb_1 _10181_ (.A_N(_02464_),
    .B_N(_04882_),
    .C(_04886_),
    .D(_02459_),
    .X(_04887_));
 sky130_fd_sc_hd__or4bb_2 _10182_ (.A(_02464_),
    .B(_04882_),
    .C_N(_04886_),
    .D_N(_02459_),
    .X(_04888_));
 sky130_fd_sc_hd__a31o_1 _10183_ (.A1(net1068),
    .A2(_02477_),
    .A3(_04883_),
    .B1(net393),
    .X(_04889_));
 sky130_fd_sc_hd__nand2b_1 _10184_ (.A_N(net1188),
    .B(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__and2_1 _10185_ (.A(\decoded_imm[30] ),
    .B(net992),
    .X(_04891_));
 sky130_fd_sc_hd__nor2_1 _10186_ (.A(\decoded_imm[30] ),
    .B(net992),
    .Y(_04892_));
 sky130_fd_sc_hd__or2_1 _10187_ (.A(_04891_),
    .B(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__nor2_1 _10188_ (.A(\decoded_imm[29] ),
    .B(net994),
    .Y(_04894_));
 sky130_fd_sc_hd__and2_1 _10189_ (.A(\decoded_imm[29] ),
    .B(net994),
    .X(_04895_));
 sky130_fd_sc_hd__xor2_1 _10190_ (.A(\decoded_imm[28] ),
    .B(net996),
    .X(_04896_));
 sky130_fd_sc_hd__or2_1 _10191_ (.A(\decoded_imm[27] ),
    .B(net998),
    .X(_04897_));
 sky130_fd_sc_hd__and2_1 _10192_ (.A(\decoded_imm[26] ),
    .B(net1000),
    .X(_04898_));
 sky130_fd_sc_hd__nor2_1 _10193_ (.A(\decoded_imm[26] ),
    .B(net1000),
    .Y(_04899_));
 sky130_fd_sc_hd__or2_1 _10194_ (.A(_04898_),
    .B(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__inv_2 _10195_ (.A(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__nor2_1 _10196_ (.A(\decoded_imm[25] ),
    .B(net1002),
    .Y(_04902_));
 sky130_fd_sc_hd__inv_2 _10197_ (.A(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__and2_1 _10198_ (.A(\decoded_imm[25] ),
    .B(net1002),
    .X(_04904_));
 sky130_fd_sc_hd__nand2_1 _10199_ (.A(\decoded_imm[24] ),
    .B(net1004),
    .Y(_04905_));
 sky130_fd_sc_hd__and2_1 _10200_ (.A(\decoded_imm[23] ),
    .B(net1006),
    .X(_04906_));
 sky130_fd_sc_hd__nor2_1 _10201_ (.A(\decoded_imm[23] ),
    .B(net218),
    .Y(_04907_));
 sky130_fd_sc_hd__nand2_1 _10202_ (.A(\decoded_imm[22] ),
    .B(net1007),
    .Y(_04908_));
 sky130_fd_sc_hd__or2_1 _10203_ (.A(\decoded_imm[22] ),
    .B(net1007),
    .X(_04909_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(_04908_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(\decoded_imm[21] ),
    .B(net1009),
    .Y(_04911_));
 sky130_fd_sc_hd__and2_1 _10206_ (.A(\decoded_imm[21] ),
    .B(net216),
    .X(_04912_));
 sky130_fd_sc_hd__nand2_1 _10207_ (.A(\decoded_imm[20] ),
    .B(net1010),
    .Y(_04913_));
 sky130_fd_sc_hd__nor2_1 _10208_ (.A(\decoded_imm[17] ),
    .B(net1017),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_1 _10209_ (.A(\decoded_imm[17] ),
    .B(net1017),
    .Y(_04915_));
 sky130_fd_sc_hd__nor2_1 _10210_ (.A(\decoded_imm[15] ),
    .B(net1020),
    .Y(_04916_));
 sky130_fd_sc_hd__nand2_1 _10211_ (.A(\decoded_imm[14] ),
    .B(net1022),
    .Y(_04917_));
 sky130_fd_sc_hd__nor2_1 _10212_ (.A(_04916_),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__and2_1 _10213_ (.A(\decoded_imm[15] ),
    .B(net1020),
    .X(_04919_));
 sky130_fd_sc_hd__nor2_1 _10214_ (.A(_04916_),
    .B(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__or2_1 _10215_ (.A(\decoded_imm[14] ),
    .B(net1022),
    .X(_04921_));
 sky130_fd_sc_hd__nand2_1 _10216_ (.A(_04917_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__and3_1 _10217_ (.A(_04917_),
    .B(_04920_),
    .C(_04921_),
    .X(_04923_));
 sky130_fd_sc_hd__nand2_1 _10218_ (.A(\decoded_imm[13] ),
    .B(net1024),
    .Y(_04924_));
 sky130_fd_sc_hd__a22o_1 _10219_ (.A1(\decoded_imm[12] ),
    .A2(net1026),
    .B1(net1024),
    .B2(\decoded_imm[13] ),
    .X(_04925_));
 sky130_fd_sc_hd__or2_1 _10220_ (.A(\decoded_imm[13] ),
    .B(net1024),
    .X(_04926_));
 sky130_fd_sc_hd__nand2_1 _10221_ (.A(_04924_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__xnor2_1 _10222_ (.A(\decoded_imm[12] ),
    .B(net1026),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _10223_ (.A(\decoded_imm[11] ),
    .B(net1028),
    .Y(_04929_));
 sky130_fd_sc_hd__or2_1 _10224_ (.A(\decoded_imm[11] ),
    .B(net1028),
    .X(_04930_));
 sky130_fd_sc_hd__nand2_1 _10225_ (.A(\decoded_imm[10] ),
    .B(net1029),
    .Y(_04931_));
 sky130_fd_sc_hd__or2_1 _10226_ (.A(\decoded_imm[10] ),
    .B(net1029),
    .X(_04932_));
 sky130_fd_sc_hd__nand2_1 _10227_ (.A(_04931_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nor2_1 _10228_ (.A(\decoded_imm[9] ),
    .B(net1031),
    .Y(_04934_));
 sky130_fd_sc_hd__nand2_1 _10229_ (.A(\decoded_imm[9] ),
    .B(net1031),
    .Y(_04935_));
 sky130_fd_sc_hd__nand2_2 _10230_ (.A(\decoded_imm[8] ),
    .B(net1033),
    .Y(_04936_));
 sky130_fd_sc_hd__and2_1 _10231_ (.A(\decoded_imm[7] ),
    .B(net1035),
    .X(_04937_));
 sky130_fd_sc_hd__nand2_1 _10232_ (.A(\decoded_imm[7] ),
    .B(net1035),
    .Y(_04938_));
 sky130_fd_sc_hd__nor2_1 _10233_ (.A(\decoded_imm[7] ),
    .B(net1035),
    .Y(_04939_));
 sky130_fd_sc_hd__or2_1 _10234_ (.A(\decoded_imm[7] ),
    .B(net1035),
    .X(_04940_));
 sky130_fd_sc_hd__nand2_1 _10235_ (.A(\decoded_imm[6] ),
    .B(net1038),
    .Y(_04941_));
 sky130_fd_sc_hd__or2_1 _10236_ (.A(\decoded_imm[6] ),
    .B(net1038),
    .X(_04942_));
 sky130_fd_sc_hd__nand2_1 _10237_ (.A(_04941_),
    .B(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__and2_1 _10238_ (.A(\decoded_imm[5] ),
    .B(net1040),
    .X(_04944_));
 sky130_fd_sc_hd__nand2_1 _10239_ (.A(\decoded_imm[5] ),
    .B(net1040),
    .Y(_04945_));
 sky130_fd_sc_hd__nor2_1 _10240_ (.A(\decoded_imm[5] ),
    .B(net1040),
    .Y(_04946_));
 sky130_fd_sc_hd__nand2_2 _10241_ (.A(\decoded_imm[4] ),
    .B(net1042),
    .Y(_04947_));
 sky130_fd_sc_hd__and2_2 _10242_ (.A(\decoded_imm[3] ),
    .B(net1044),
    .X(_04948_));
 sky130_fd_sc_hd__nand2_1 _10243_ (.A(\decoded_imm[2] ),
    .B(net1045),
    .Y(_04949_));
 sky130_fd_sc_hd__and2_1 _10244_ (.A(net1047),
    .B(\decoded_imm[1] ),
    .X(_04950_));
 sky130_fd_sc_hd__nand2_1 _10245_ (.A(net1047),
    .B(\decoded_imm[1] ),
    .Y(_04951_));
 sky130_fd_sc_hd__or2_1 _10246_ (.A(net1047),
    .B(\decoded_imm[1] ),
    .X(_04952_));
 sky130_fd_sc_hd__nand4_1 _10247_ (.A(net1051),
    .B(\decoded_imm[0] ),
    .C(_04951_),
    .D(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__a31o_1 _10248_ (.A1(net1051),
    .A2(\decoded_imm[0] ),
    .A3(_04952_),
    .B1(_04950_),
    .X(_04954_));
 sky130_fd_sc_hd__or2_1 _10249_ (.A(\decoded_imm[2] ),
    .B(net1045),
    .X(_04955_));
 sky130_fd_sc_hd__nand3_1 _10250_ (.A(_04949_),
    .B(_04954_),
    .C(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__nor2_1 _10251_ (.A(\decoded_imm[3] ),
    .B(net1044),
    .Y(_04957_));
 sky130_fd_sc_hd__a211oi_2 _10252_ (.A1(_04949_),
    .A2(_04956_),
    .B1(_04957_),
    .C1(_04948_),
    .Y(_04958_));
 sky130_fd_sc_hd__or2_1 _10253_ (.A(\decoded_imm[4] ),
    .B(net1042),
    .X(_04959_));
 sky130_fd_sc_hd__o211ai_2 _10254_ (.A1(_04948_),
    .A2(_04958_),
    .B1(_04959_),
    .C1(_04947_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_1 _10255_ (.A(_04947_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__a31o_1 _10256_ (.A1(_04945_),
    .A2(_04947_),
    .A3(_04960_),
    .B1(_04946_),
    .X(_04962_));
 sky130_fd_sc_hd__o21ai_1 _10257_ (.A1(_04943_),
    .A2(_04962_),
    .B1(_04941_),
    .Y(_04963_));
 sky130_fd_sc_hd__nand3_1 _10258_ (.A(\decoded_imm[6] ),
    .B(net1038),
    .C(_04940_),
    .Y(_04964_));
 sky130_fd_sc_hd__nor2_1 _10259_ (.A(_04937_),
    .B(_04939_),
    .Y(_04965_));
 sky130_fd_sc_hd__or3_1 _10260_ (.A(_04937_),
    .B(_04939_),
    .C(_04943_),
    .X(_04966_));
 sky130_fd_sc_hd__a211o_1 _10261_ (.A1(_04945_),
    .A2(_04947_),
    .B1(_04966_),
    .C1(_04946_),
    .X(_04967_));
 sky130_fd_sc_hd__nor2_1 _10262_ (.A(_04944_),
    .B(_04946_),
    .Y(_04968_));
 sky130_fd_sc_hd__and2b_1 _10263_ (.A_N(_04966_),
    .B(_04968_),
    .X(_04969_));
 sky130_fd_sc_hd__o2111ai_1 _10264_ (.A1(_04948_),
    .A2(_04958_),
    .B1(_04959_),
    .C1(_04969_),
    .D1(_04947_),
    .Y(_04970_));
 sky130_fd_sc_hd__or2_1 _10265_ (.A(\decoded_imm[8] ),
    .B(net1033),
    .X(_04971_));
 sky130_fd_sc_hd__nand2_1 _10266_ (.A(_04936_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__a41o_1 _10267_ (.A1(_04938_),
    .A2(_04964_),
    .A3(_04967_),
    .A4(_04970_),
    .B1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__nand2_1 _10268_ (.A(_04936_),
    .B(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__a31o_1 _10269_ (.A1(_04935_),
    .A2(_04936_),
    .A3(_04973_),
    .B1(_04934_),
    .X(_04975_));
 sky130_fd_sc_hd__or2_1 _10270_ (.A(_04933_),
    .B(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__nand2_1 _10271_ (.A(_04931_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__a21bo_1 _10272_ (.A1(_04929_),
    .A2(_04931_),
    .B1_N(_04930_),
    .X(_04978_));
 sky130_fd_sc_hd__nand2_1 _10273_ (.A(_04929_),
    .B(_04930_),
    .Y(_04979_));
 sky130_fd_sc_hd__or2_1 _10274_ (.A(_04933_),
    .B(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__and2b_1 _10275_ (.A_N(_04934_),
    .B(_04935_),
    .X(_04981_));
 sky130_fd_sc_hd__a311o_1 _10276_ (.A1(_04935_),
    .A2(_04936_),
    .A3(_04973_),
    .B1(_04980_),
    .C1(_04934_),
    .X(_04982_));
 sky130_fd_sc_hd__a21oi_1 _10277_ (.A1(_04978_),
    .A2(_04982_),
    .B1(_04928_),
    .Y(_04983_));
 sky130_fd_sc_hd__o21ai_1 _10278_ (.A1(_04925_),
    .A2(_04983_),
    .B1(_04926_),
    .Y(_04984_));
 sky130_fd_sc_hd__and3_1 _10279_ (.A(_04923_),
    .B(_04924_),
    .C(_04926_),
    .X(_04985_));
 sky130_fd_sc_hd__inv_2 _10280_ (.A(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__a211o_1 _10281_ (.A1(_04978_),
    .A2(_04982_),
    .B1(_04986_),
    .C1(_04928_),
    .X(_04987_));
 sky130_fd_sc_hd__a311o_1 _10282_ (.A1(_04923_),
    .A2(_04925_),
    .A3(_04926_),
    .B1(_04919_),
    .C1(_04918_),
    .X(_04988_));
 sky130_fd_sc_hd__inv_2 _10283_ (.A(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__xnor2_1 _10284_ (.A(\decoded_imm[16] ),
    .B(net1018),
    .Y(_04990_));
 sky130_fd_sc_hd__a21oi_1 _10285_ (.A1(_04987_),
    .A2(_04989_),
    .B1(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__a21oi_1 _10286_ (.A1(\decoded_imm[16] ),
    .A2(net1018),
    .B1(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__o211a_1 _10287_ (.A1(\decoded_imm[17] ),
    .A2(net1017),
    .B1(net1018),
    .C1(\decoded_imm[16] ),
    .X(_04993_));
 sky130_fd_sc_hd__nand2b_1 _10288_ (.A_N(_04914_),
    .B(_04915_),
    .Y(_04994_));
 sky130_fd_sc_hd__a211o_1 _10289_ (.A1(_04987_),
    .A2(_04989_),
    .B1(_04990_),
    .C1(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__a21o_1 _10290_ (.A1(_04915_),
    .A2(_04992_),
    .B1(_04914_),
    .X(_04996_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(\decoded_imm[19] ),
    .B(net1012),
    .Y(_04997_));
 sky130_fd_sc_hd__inv_2 _10292_ (.A(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__nor2_1 _10293_ (.A(\decoded_imm[19] ),
    .B(net1012),
    .Y(_04999_));
 sky130_fd_sc_hd__and2_1 _10294_ (.A(\decoded_imm[18] ),
    .B(net1014),
    .X(_05000_));
 sky130_fd_sc_hd__nand2_1 _10295_ (.A(\decoded_imm[18] ),
    .B(net1014),
    .Y(_05001_));
 sky130_fd_sc_hd__o21a_1 _10296_ (.A1(_04999_),
    .A2(_05001_),
    .B1(_04997_),
    .X(_05002_));
 sky130_fd_sc_hd__and4b_1 _10297_ (.A_N(_04993_),
    .B(_05002_),
    .C(_04995_),
    .D(_04915_),
    .X(_05003_));
 sky130_fd_sc_hd__nor2_1 _10298_ (.A(\decoded_imm[18] ),
    .B(net1014),
    .Y(_05004_));
 sky130_fd_sc_hd__a21o_1 _10299_ (.A1(_04997_),
    .A2(_05004_),
    .B1(_04999_),
    .X(_05005_));
 sky130_fd_sc_hd__or2_1 _10300_ (.A(\decoded_imm[20] ),
    .B(net1010),
    .X(_05006_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(_04913_),
    .B(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__or3_1 _10302_ (.A(_05003_),
    .B(_05005_),
    .C(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__nand2_1 _10303_ (.A(_04913_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__and2b_1 _10304_ (.A_N(_04912_),
    .B(_04913_),
    .X(_05010_));
 sky130_fd_sc_hd__a21o_1 _10305_ (.A1(_05008_),
    .A2(_05010_),
    .B1(_04911_),
    .X(_05011_));
 sky130_fd_sc_hd__or2_1 _10306_ (.A(_04910_),
    .B(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__nand2_1 _10307_ (.A(_04908_),
    .B(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__and2b_1 _10308_ (.A_N(_04906_),
    .B(_04908_),
    .X(_05014_));
 sky130_fd_sc_hd__or2_1 _10309_ (.A(_04906_),
    .B(_04907_),
    .X(_05015_));
 sky130_fd_sc_hd__or2_1 _10310_ (.A(_04910_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__or3_1 _10311_ (.A(_04911_),
    .B(_05010_),
    .C(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__nor2_1 _10312_ (.A(_04911_),
    .B(_04912_),
    .Y(_05018_));
 sky130_fd_sc_hd__or3b_1 _10313_ (.A(_05007_),
    .B(_05016_),
    .C_N(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__or3_1 _10314_ (.A(_05003_),
    .B(_05005_),
    .C(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__o211a_1 _10315_ (.A1(_04907_),
    .A2(_05014_),
    .B1(_05017_),
    .C1(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__or2_1 _10316_ (.A(\decoded_imm[24] ),
    .B(net1004),
    .X(_05022_));
 sky130_fd_sc_hd__nand2_1 _10317_ (.A(_04905_),
    .B(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__o21ai_2 _10318_ (.A1(_05021_),
    .A2(_05023_),
    .B1(_04905_),
    .Y(_05024_));
 sky130_fd_sc_hd__nor2_1 _10319_ (.A(_04904_),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__o211a_1 _10320_ (.A1(_04904_),
    .A2(_05024_),
    .B1(_04901_),
    .C1(_04903_),
    .X(_05026_));
 sky130_fd_sc_hd__and2_1 _10321_ (.A(\decoded_imm[27] ),
    .B(net998),
    .X(_05027_));
 sky130_fd_sc_hd__nand2_1 _10322_ (.A(\decoded_imm[27] ),
    .B(net998),
    .Y(_05028_));
 sky130_fd_sc_hd__nor2_1 _10323_ (.A(_04902_),
    .B(_04904_),
    .Y(_05029_));
 sky130_fd_sc_hd__o31a_1 _10324_ (.A1(_04898_),
    .A2(_05026_),
    .A3(_05027_),
    .B1(_04897_),
    .X(_05030_));
 sky130_fd_sc_hd__a22o_1 _10325_ (.A1(\decoded_imm[28] ),
    .A2(net996),
    .B1(_04896_),
    .B2(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__nor2_1 _10326_ (.A(_04895_),
    .B(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__nor2_1 _10327_ (.A(_04894_),
    .B(_04895_),
    .Y(_05033_));
 sky130_fd_sc_hd__nor3_1 _10328_ (.A(_04893_),
    .B(_04894_),
    .C(_05032_),
    .Y(_05034_));
 sky130_fd_sc_hd__or2_1 _10329_ (.A(net1188),
    .B(\decoded_imm[31] ),
    .X(_05035_));
 sky130_fd_sc_hd__nand2_1 _10330_ (.A(net1188),
    .B(\decoded_imm[31] ),
    .Y(_05036_));
 sky130_fd_sc_hd__a211o_1 _10331_ (.A1(_05035_),
    .A2(_05036_),
    .B1(_04891_),
    .C1(_05034_),
    .X(_05037_));
 sky130_fd_sc_hd__o211ai_1 _10332_ (.A1(_04891_),
    .A2(_05034_),
    .B1(_05035_),
    .C1(_05036_),
    .Y(_05038_));
 sky130_fd_sc_hd__and3_1 _10333_ (.A(net958),
    .B(_05037_),
    .C(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__or2_1 _10334_ (.A(is_lui_auipc_jal),
    .B(_04880_),
    .X(_05040_));
 sky130_fd_sc_hd__mux2_1 _10335_ (.A0(\cpuregs[6][31] ),
    .A1(\cpuregs[7][31] ),
    .S(net692),
    .X(_05041_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(\cpuregs[4][31] ),
    .A1(\cpuregs[5][31] ),
    .S(net695),
    .X(_05042_));
 sky130_fd_sc_hd__mux2_1 _10337_ (.A0(_05041_),
    .A1(_05042_),
    .S(net818),
    .X(_05043_));
 sky130_fd_sc_hd__or2_1 _10338_ (.A(\cpuregs[0][31] ),
    .B(net694),
    .X(_05044_));
 sky130_fd_sc_hd__o211a_1 _10339_ (.A1(\cpuregs[1][31] ),
    .A2(net639),
    .B1(net613),
    .C1(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__or2_1 _10340_ (.A(\cpuregs[2][31] ),
    .B(net695),
    .X(_05046_));
 sky130_fd_sc_hd__o211a_1 _10341_ (.A1(\cpuregs[3][31] ),
    .A2(net638),
    .B1(net599),
    .C1(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__a211o_1 _10342_ (.A1(net833),
    .A2(_05043_),
    .B1(_05047_),
    .C1(net784),
    .X(_05048_));
 sky130_fd_sc_hd__mux2_1 _10343_ (.A0(\cpuregs[14][31] ),
    .A1(\cpuregs[15][31] ),
    .S(net695),
    .X(_05049_));
 sky130_fd_sc_hd__mux2_1 _10344_ (.A0(\cpuregs[12][31] ),
    .A1(\cpuregs[13][31] ),
    .S(net694),
    .X(_05050_));
 sky130_fd_sc_hd__or2_1 _10345_ (.A(net806),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__o211a_1 _10346_ (.A1(net817),
    .A2(_05049_),
    .B1(_05051_),
    .C1(net833),
    .X(_05052_));
 sky130_fd_sc_hd__or2_1 _10347_ (.A(\cpuregs[8][31] ),
    .B(net694),
    .X(_05053_));
 sky130_fd_sc_hd__o211a_1 _10348_ (.A1(\cpuregs[9][31] ),
    .A2(net638),
    .B1(net612),
    .C1(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__or2_1 _10349_ (.A(\cpuregs[10][31] ),
    .B(net694),
    .X(_05055_));
 sky130_fd_sc_hd__o211a_1 _10350_ (.A1(\cpuregs[11][31] ),
    .A2(net638),
    .B1(net599),
    .C1(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__or4_1 _10351_ (.A(net792),
    .B(_05052_),
    .C(_05054_),
    .D(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__o21a_1 _10352_ (.A1(_05045_),
    .A2(_05048_),
    .B1(_03171_),
    .X(_05058_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(\cpuregs[20][31] ),
    .A1(\cpuregs[21][31] ),
    .S(net693),
    .X(_05059_));
 sky130_fd_sc_hd__mux2_1 _10354_ (.A0(\cpuregs[22][31] ),
    .A1(\cpuregs[23][31] ),
    .S(net693),
    .X(_05060_));
 sky130_fd_sc_hd__mux2_1 _10355_ (.A0(_05059_),
    .A1(_05060_),
    .S(net806),
    .X(_05061_));
 sky130_fd_sc_hd__or2_1 _10356_ (.A(\cpuregs[16][31] ),
    .B(net692),
    .X(_05062_));
 sky130_fd_sc_hd__o211a_1 _10357_ (.A1(\cpuregs[17][31] ),
    .A2(net638),
    .B1(net613),
    .C1(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__o21a_1 _10358_ (.A1(\cpuregs[19][31] ),
    .A2(net638),
    .B1(net599),
    .X(_05064_));
 sky130_fd_sc_hd__o22a_1 _10359_ (.A1(\cpuregs[18][31] ),
    .A2(net554),
    .B1(_05064_),
    .B2(net783),
    .X(_05065_));
 sky130_fd_sc_hd__a211o_1 _10360_ (.A1(net833),
    .A2(_05061_),
    .B1(_05063_),
    .C1(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__mux2_1 _10361_ (.A0(\cpuregs[30][31] ),
    .A1(\cpuregs[31][31] ),
    .S(net694),
    .X(_05067_));
 sky130_fd_sc_hd__mux2_1 _10362_ (.A0(\cpuregs[28][31] ),
    .A1(\cpuregs[29][31] ),
    .S(net694),
    .X(_05068_));
 sky130_fd_sc_hd__mux2_1 _10363_ (.A0(_05067_),
    .A1(_05068_),
    .S(net817),
    .X(_05069_));
 sky130_fd_sc_hd__or2_1 _10364_ (.A(\cpuregs[24][31] ),
    .B(net693),
    .X(_05070_));
 sky130_fd_sc_hd__o211a_1 _10365_ (.A1(\cpuregs[25][31] ),
    .A2(net638),
    .B1(net613),
    .C1(_05070_),
    .X(_05071_));
 sky130_fd_sc_hd__or2_1 _10366_ (.A(\cpuregs[26][31] ),
    .B(net693),
    .X(_05072_));
 sky130_fd_sc_hd__o211a_1 _10367_ (.A1(\cpuregs[27][31] ),
    .A2(net638),
    .B1(net599),
    .C1(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__a2111o_1 _10368_ (.A1(net833),
    .A2(_05069_),
    .B1(_05071_),
    .C1(_05073_),
    .D1(net793),
    .X(_05074_));
 sky130_fd_sc_hd__and3_1 _10369_ (.A(net774),
    .B(_05066_),
    .C(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a21oi_4 _10370_ (.A1(_05057_),
    .A2(_05058_),
    .B1(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__nor2_1 _10371_ (.A(net569),
    .B(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__mux2_1 _10372_ (.A0(net999),
    .A1(net992),
    .S(_02474_),
    .X(_05078_));
 sky130_fd_sc_hd__and2b_1 _10373_ (.A_N(instr_lui),
    .B(is_lui_auipc_jal),
    .X(_05079_));
 sky130_fd_sc_hd__and2_1 _10374_ (.A(_04879_),
    .B(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__a32o_1 _10375_ (.A1(net1068),
    .A2(net760),
    .A3(_05078_),
    .B1(net566),
    .B2(\reg_pc[31] ),
    .X(_05081_));
 sky130_fd_sc_hd__o41a_1 _10376_ (.A1(_04889_),
    .A2(_05039_),
    .A3(_05077_),
    .A4(_05081_),
    .B1(_04890_),
    .X(_00773_));
 sky130_fd_sc_hd__and2b_2 _10377_ (.A_N(\genblk2.pcpi_div.pcpi_wait_q ),
    .B(\genblk2.pcpi_div.pcpi_wait ),
    .X(_05082_));
 sky130_fd_sc_hd__nand2b_1 _10378_ (.A_N(\genblk2.pcpi_div.pcpi_wait_q ),
    .B(\genblk2.pcpi_div.pcpi_wait ),
    .Y(_05083_));
 sky130_fd_sc_hd__or4_1 _10379_ (.A(\genblk2.pcpi_div.quotient_msk[11] ),
    .B(\genblk2.pcpi_div.quotient_msk[10] ),
    .C(\genblk2.pcpi_div.quotient_msk[9] ),
    .D(\genblk2.pcpi_div.quotient_msk[8] ),
    .X(_05084_));
 sky130_fd_sc_hd__or4_1 _10380_ (.A(\genblk2.pcpi_div.quotient_msk[15] ),
    .B(\genblk2.pcpi_div.quotient_msk[14] ),
    .C(\genblk2.pcpi_div.quotient_msk[13] ),
    .D(\genblk2.pcpi_div.quotient_msk[12] ),
    .X(_05085_));
 sky130_fd_sc_hd__or4_1 _10381_ (.A(\genblk2.pcpi_div.quotient_msk[7] ),
    .B(\genblk2.pcpi_div.quotient_msk[6] ),
    .C(\genblk2.pcpi_div.quotient_msk[5] ),
    .D(\genblk2.pcpi_div.quotient_msk[4] ),
    .X(_05086_));
 sky130_fd_sc_hd__or4_1 _10382_ (.A(\genblk2.pcpi_div.quotient_msk[3] ),
    .B(\genblk2.pcpi_div.quotient_msk[2] ),
    .C(\genblk2.pcpi_div.quotient_msk[1] ),
    .D(\genblk2.pcpi_div.quotient_msk[0] ),
    .X(_05087_));
 sky130_fd_sc_hd__or3_1 _10383_ (.A(_05084_),
    .B(_05085_),
    .C(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__or4_1 _10384_ (.A(\genblk2.pcpi_div.quotient_msk[27] ),
    .B(\genblk2.pcpi_div.quotient_msk[26] ),
    .C(\genblk2.pcpi_div.quotient_msk[25] ),
    .D(\genblk2.pcpi_div.quotient_msk[24] ),
    .X(_05089_));
 sky130_fd_sc_hd__or4_1 _10385_ (.A(\genblk2.pcpi_div.quotient_msk[31] ),
    .B(\genblk2.pcpi_div.quotient_msk[30] ),
    .C(\genblk2.pcpi_div.quotient_msk[29] ),
    .D(\genblk2.pcpi_div.quotient_msk[28] ),
    .X(_05090_));
 sky130_fd_sc_hd__or4_1 _10386_ (.A(\genblk2.pcpi_div.quotient_msk[23] ),
    .B(\genblk2.pcpi_div.quotient_msk[22] ),
    .C(\genblk2.pcpi_div.quotient_msk[21] ),
    .D(\genblk2.pcpi_div.quotient_msk[20] ),
    .X(_05091_));
 sky130_fd_sc_hd__or4_1 _10387_ (.A(\genblk2.pcpi_div.quotient_msk[19] ),
    .B(\genblk2.pcpi_div.quotient_msk[18] ),
    .C(\genblk2.pcpi_div.quotient_msk[17] ),
    .D(\genblk2.pcpi_div.quotient_msk[16] ),
    .X(_05092_));
 sky130_fd_sc_hd__or3_1 _10388_ (.A(_05089_),
    .B(_05090_),
    .C(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__or4_1 _10389_ (.A(_05086_),
    .B(_05088_),
    .C(_05091_),
    .D(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_1 _10390_ (.A(_02362_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _10391_ (.A(net864),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__nand2_1 _10392_ (.A(net1223),
    .B(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__or4_2 _10393_ (.A(net1180),
    .B(net1178),
    .C(net1176),
    .D(net1177),
    .X(_05098_));
 sky130_fd_sc_hd__or2_1 _10394_ (.A(net1174),
    .B(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__or4_1 _10395_ (.A(net1172),
    .B(net1174),
    .C(net1171),
    .D(_05098_),
    .X(_05100_));
 sky130_fd_sc_hd__or3_1 _10396_ (.A(net1169),
    .B(net1168),
    .C(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__or2_1 _10397_ (.A(net1167),
    .B(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__nor2_1 _10398_ (.A(net1166),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__or3_1 _10399_ (.A(net1165),
    .B(net1166),
    .C(_05102_),
    .X(_05104_));
 sky130_fd_sc_hd__or2_1 _10400_ (.A(net1164),
    .B(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__nor2_1 _10401_ (.A(net1163),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__or3_1 _10402_ (.A(net1163),
    .B(net240),
    .C(_05105_),
    .X(_05107_));
 sky130_fd_sc_hd__or2_1 _10403_ (.A(net1162),
    .B(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__nor2_1 _10404_ (.A(net1161),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__or3_1 _10405_ (.A(net1160),
    .B(net1161),
    .C(_05108_),
    .X(_05110_));
 sky130_fd_sc_hd__or2_1 _10406_ (.A(net244),
    .B(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__or3_1 _10407_ (.A(net1159),
    .B(net247),
    .C(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__or2_1 _10408_ (.A(net248),
    .B(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__or3_2 _10409_ (.A(net250),
    .B(net1158),
    .C(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__or3_1 _10410_ (.A(net252),
    .B(net251),
    .C(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__or2_1 _10411_ (.A(net253),
    .B(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__or2_1 _10412_ (.A(net254),
    .B(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__or3_1 _10413_ (.A(net256),
    .B(net255),
    .C(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__o21ai_1 _10414_ (.A1(net258),
    .A2(_05118_),
    .B1(_02507_),
    .Y(_05119_));
 sky130_fd_sc_hd__nor2_2 _10415_ (.A(net1214),
    .B(_05083_),
    .Y(_05120_));
 sky130_fd_sc_hd__a32o_1 _10416_ (.A1(net1157),
    .A2(_05119_),
    .A3(_05120_),
    .B1(net389),
    .B2(net2455),
    .X(_00774_));
 sky130_fd_sc_hd__nor2_1 _10417_ (.A(net1208),
    .B(_02451_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand2_1 _10418_ (.A(net2852),
    .B(_02490_),
    .Y(_05122_));
 sky130_fd_sc_hd__o211a_1 _10419_ (.A1(mem_do_prefetch),
    .A2(_02490_),
    .B1(_05121_),
    .C1(_05122_),
    .X(_00775_));
 sky130_fd_sc_hd__nor2_1 _10420_ (.A(net1088),
    .B(\cpu_state[0] ),
    .Y(_05123_));
 sky130_fd_sc_hd__and3_1 _10421_ (.A(_02379_),
    .B(net880),
    .C(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__or3_2 _10422_ (.A(net1081),
    .B(net1088),
    .C(net1068),
    .X(_05125_));
 sky130_fd_sc_hd__o21ai_1 _10423_ (.A1(net1089),
    .A2(_05125_),
    .B1(_02503_),
    .Y(_05126_));
 sky130_fd_sc_hd__o31a_1 _10424_ (.A1(_02439_),
    .A2(_02493_),
    .A3(_05126_),
    .B1(_05121_),
    .X(_05127_));
 sky130_fd_sc_hd__a21oi_1 _10425_ (.A1(net1087),
    .A2(is_sb_sh_sw),
    .B1(mem_do_prefetch),
    .Y(_05128_));
 sky130_fd_sc_hd__nand4_1 _10426_ (.A(_02437_),
    .B(_02491_),
    .C(_05125_),
    .D(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__o211a_1 _10427_ (.A1(_02489_),
    .A2(_05125_),
    .B1(_05129_),
    .C1(_05121_),
    .X(_05130_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(_05130_),
    .A1(mem_do_rinst),
    .S(_05127_),
    .X(_05131_));
 sky130_fd_sc_hd__a41o_1 _10429_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(_03457_),
    .A3(_04881_),
    .A4(_05124_),
    .B1(_05131_),
    .X(_00776_));
 sky130_fd_sc_hd__a21o_1 _10430_ (.A1(net3008),
    .A2(_05121_),
    .B1(net410),
    .X(_00777_));
 sky130_fd_sc_hd__and3b_1 _10431_ (.A_N(mem_do_wdata),
    .B(_02702_),
    .C(_05124_),
    .X(_05132_));
 sky130_fd_sc_hd__a22o_1 _10432_ (.A1(mem_do_wdata),
    .A2(_05121_),
    .B1(_05132_),
    .B2(_02453_),
    .X(_00778_));
 sky130_fd_sc_hd__o21a_1 _10433_ (.A1(net1083),
    .A2(net1088),
    .B1(net1231),
    .X(_05133_));
 sky130_fd_sc_hd__o21ai_2 _10434_ (.A1(net1083),
    .A2(net1088),
    .B1(net1231),
    .Y(_05134_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(\cpuregs[6][0] ),
    .A1(\cpuregs[7][0] ),
    .S(net684),
    .X(_05135_));
 sky130_fd_sc_hd__mux2_1 _10436_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .S(net697),
    .X(_05136_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(_05135_),
    .A1(_05136_),
    .S(net818),
    .X(_05137_));
 sky130_fd_sc_hd__or2_1 _10438_ (.A(\cpuregs[2][0] ),
    .B(net685),
    .X(_05138_));
 sky130_fd_sc_hd__o211a_1 _10439_ (.A1(\cpuregs[3][0] ),
    .A2(net634),
    .B1(net597),
    .C1(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__o21a_1 _10440_ (.A1(\cpuregs[1][0] ),
    .A2(net635),
    .B1(net611),
    .X(_05140_));
 sky130_fd_sc_hd__o22a_1 _10441_ (.A1(\cpuregs[0][0] ),
    .A2(net555),
    .B1(_05140_),
    .B2(net785),
    .X(_05141_));
 sky130_fd_sc_hd__a211o_1 _10442_ (.A1(net831),
    .A2(_05137_),
    .B1(_05139_),
    .C1(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .S(net685),
    .X(_05143_));
 sky130_fd_sc_hd__mux2_1 _10444_ (.A0(\cpuregs[14][0] ),
    .A1(\cpuregs[15][0] ),
    .S(net685),
    .X(_05144_));
 sky130_fd_sc_hd__mux2_1 _10445_ (.A0(_05143_),
    .A1(_05144_),
    .S(net804),
    .X(_05145_));
 sky130_fd_sc_hd__or2_1 _10446_ (.A(\cpuregs[10][0] ),
    .B(net684),
    .X(_05146_));
 sky130_fd_sc_hd__o211a_1 _10447_ (.A1(\cpuregs[11][0] ),
    .A2(net634),
    .B1(net600),
    .C1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__mux2_1 _10448_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .S(net686),
    .X(_05148_));
 sky130_fd_sc_hd__a31o_1 _10449_ (.A1(net839),
    .A2(net816),
    .A3(_05148_),
    .B1(net792),
    .X(_05149_));
 sky130_fd_sc_hd__a211o_1 _10450_ (.A1(net834),
    .A2(_05145_),
    .B1(_05147_),
    .C1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__mux2_1 _10451_ (.A0(\cpuregs[22][0] ),
    .A1(\cpuregs[23][0] ),
    .S(net687),
    .X(_05151_));
 sky130_fd_sc_hd__mux2_1 _10452_ (.A0(\cpuregs[20][0] ),
    .A1(\cpuregs[21][0] ),
    .S(net687),
    .X(_05152_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(_05151_),
    .A1(_05152_),
    .S(net816),
    .X(_05153_));
 sky130_fd_sc_hd__or2_1 _10454_ (.A(\cpuregs[18][0] ),
    .B(net686),
    .X(_05154_));
 sky130_fd_sc_hd__o211a_1 _10455_ (.A1(\cpuregs[19][0] ),
    .A2(net635),
    .B1(net600),
    .C1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__o21a_1 _10456_ (.A1(\cpuregs[17][0] ),
    .A2(net635),
    .B1(net611),
    .X(_05156_));
 sky130_fd_sc_hd__o22a_1 _10457_ (.A1(\cpuregs[16][0] ),
    .A2(net554),
    .B1(_05156_),
    .B2(net784),
    .X(_05157_));
 sky130_fd_sc_hd__a211o_1 _10458_ (.A1(net834),
    .A2(_05153_),
    .B1(_05155_),
    .C1(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(\cpuregs[28][0] ),
    .A1(\cpuregs[29][0] ),
    .S(net684),
    .X(_05159_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(\cpuregs[30][0] ),
    .A1(\cpuregs[31][0] ),
    .S(net684),
    .X(_05160_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(_05159_),
    .A1(_05160_),
    .S(net804),
    .X(_05161_));
 sky130_fd_sc_hd__or2_1 _10462_ (.A(\cpuregs[24][0] ),
    .B(net684),
    .X(_05162_));
 sky130_fd_sc_hd__o211a_1 _10463_ (.A1(\cpuregs[25][0] ),
    .A2(net634),
    .B1(net611),
    .C1(_05162_),
    .X(_05163_));
 sky130_fd_sc_hd__or2_1 _10464_ (.A(\cpuregs[26][0] ),
    .B(net684),
    .X(_05164_));
 sky130_fd_sc_hd__o211a_1 _10465_ (.A1(\cpuregs[27][0] ),
    .A2(net634),
    .B1(net600),
    .C1(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__a211o_1 _10466_ (.A1(net834),
    .A2(_05161_),
    .B1(_05163_),
    .C1(net792),
    .X(_05166_));
 sky130_fd_sc_hd__o211a_1 _10467_ (.A1(_05165_),
    .A2(_05166_),
    .B1(net774),
    .C1(_05158_),
    .X(_05167_));
 sky130_fd_sc_hd__a31oi_4 _10468_ (.A1(_03171_),
    .A2(_05142_),
    .A3(_05150_),
    .B1(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__nor2_1 _10469_ (.A(net987),
    .B(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__a21o_1 _10470_ (.A1(net987),
    .A2(\decoded_imm[0] ),
    .B1(net856),
    .X(_05170_));
 sky130_fd_sc_hd__o22a_1 _10471_ (.A1(net1181),
    .A2(net860),
    .B1(_05169_),
    .B2(_05170_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(\cpuregs[6][1] ),
    .A1(\cpuregs[7][1] ),
    .S(net686),
    .X(_05171_));
 sky130_fd_sc_hd__or2_1 _10473_ (.A(\cpuregs[4][1] ),
    .B(net692),
    .X(_05172_));
 sky130_fd_sc_hd__o211a_1 _10474_ (.A1(\cpuregs[5][1] ),
    .A2(net636),
    .B1(net817),
    .C1(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__a211o_1 _10475_ (.A1(net806),
    .A2(_05171_),
    .B1(_05173_),
    .C1(net839),
    .X(_05174_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(\cpuregs[2][1] ),
    .A1(\cpuregs[3][1] ),
    .S(net688),
    .X(_05175_));
 sky130_fd_sc_hd__a221o_1 _10477_ (.A1(\cpuregs[1][1] ),
    .A2(net551),
    .B1(_05175_),
    .B2(net805),
    .C1(net832),
    .X(_05176_));
 sky130_fd_sc_hd__a21o_1 _10478_ (.A1(_05174_),
    .A2(_05176_),
    .B1(net783),
    .X(_05177_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\cpuregs[12][1] ),
    .A1(\cpuregs[13][1] ),
    .S(net682),
    .X(_05178_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(\cpuregs[14][1] ),
    .A1(\cpuregs[15][1] ),
    .S(net683),
    .X(_05179_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(_05178_),
    .A1(_05179_),
    .S(net804),
    .X(_05180_));
 sky130_fd_sc_hd__or2_1 _10482_ (.A(\cpuregs[8][1] ),
    .B(net682),
    .X(_05181_));
 sky130_fd_sc_hd__o211a_1 _10483_ (.A1(\cpuregs[9][1] ),
    .A2(net632),
    .B1(net610),
    .C1(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__or2_1 _10484_ (.A(\cpuregs[10][1] ),
    .B(net682),
    .X(_05183_));
 sky130_fd_sc_hd__o211a_1 _10485_ (.A1(\cpuregs[11][1] ),
    .A2(net633),
    .B1(net597),
    .C1(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__a211o_1 _10486_ (.A1(net831),
    .A2(_05180_),
    .B1(_05182_),
    .C1(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__o211a_1 _10487_ (.A1(net792),
    .A2(_05185_),
    .B1(_05177_),
    .C1(net778),
    .X(_05186_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(\cpuregs[30][1] ),
    .A1(\cpuregs[31][1] ),
    .S(net686),
    .X(_05187_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(\cpuregs[28][1] ),
    .A1(\cpuregs[29][1] ),
    .S(net683),
    .X(_05188_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(_05187_),
    .A1(_05188_),
    .S(net816),
    .X(_05189_));
 sky130_fd_sc_hd__or2_1 _10491_ (.A(\cpuregs[24][1] ),
    .B(net683),
    .X(_05190_));
 sky130_fd_sc_hd__o211a_1 _10492_ (.A1(\cpuregs[25][1] ),
    .A2(net636),
    .B1(net612),
    .C1(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__or2_1 _10493_ (.A(\cpuregs[26][1] ),
    .B(net691),
    .X(_05192_));
 sky130_fd_sc_hd__o211a_1 _10494_ (.A1(\cpuregs[27][1] ),
    .A2(net636),
    .B1(net598),
    .C1(_05192_),
    .X(_05193_));
 sky130_fd_sc_hd__a2111o_1 _10495_ (.A1(net832),
    .A2(_05189_),
    .B1(_05191_),
    .C1(_05193_),
    .D1(net793),
    .X(_05194_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(\cpuregs[20][1] ),
    .A1(\cpuregs[21][1] ),
    .S(net688),
    .X(_05195_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(\cpuregs[22][1] ),
    .A1(\cpuregs[23][1] ),
    .S(net688),
    .X(_05196_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(_05195_),
    .A1(_05196_),
    .S(net805),
    .X(_05197_));
 sky130_fd_sc_hd__or2_1 _10499_ (.A(\cpuregs[16][1] ),
    .B(net688),
    .X(_05198_));
 sky130_fd_sc_hd__o211a_1 _10500_ (.A1(\cpuregs[17][1] ),
    .A2(net636),
    .B1(net612),
    .C1(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__o21a_1 _10501_ (.A1(\cpuregs[19][1] ),
    .A2(net636),
    .B1(net598),
    .X(_05200_));
 sky130_fd_sc_hd__o22a_1 _10502_ (.A1(\cpuregs[18][1] ),
    .A2(net554),
    .B1(_05200_),
    .B2(net783),
    .X(_05201_));
 sky130_fd_sc_hd__a211o_1 _10503_ (.A1(net832),
    .A2(_05197_),
    .B1(_05199_),
    .C1(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__a31oi_4 _10504_ (.A1(net774),
    .A2(_05194_),
    .A3(_05202_),
    .B1(_05186_),
    .Y(_05203_));
 sky130_fd_sc_hd__nor2_1 _10505_ (.A(net987),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__a21o_1 _10506_ (.A1(net986),
    .A2(\decoded_imm[1] ),
    .B1(net856),
    .X(_05205_));
 sky130_fd_sc_hd__o22a_1 _10507_ (.A1(net1179),
    .A2(net860),
    .B1(_05204_),
    .B2(_05205_),
    .X(_00780_));
 sky130_fd_sc_hd__a21o_1 _10508_ (.A1(net987),
    .A2(\decoded_imm[2] ),
    .B1(net856),
    .X(_05206_));
 sky130_fd_sc_hd__o22a_1 _10509_ (.A1(net119),
    .A2(net860),
    .B1(_05206_),
    .B2(_03190_),
    .X(_00781_));
 sky130_fd_sc_hd__a21o_1 _10510_ (.A1(net987),
    .A2(\decoded_imm[3] ),
    .B1(net856),
    .X(_05207_));
 sky130_fd_sc_hd__o22a_1 _10511_ (.A1(net1176),
    .A2(net860),
    .B1(_05207_),
    .B2(_03228_),
    .X(_00782_));
 sky130_fd_sc_hd__a21o_1 _10512_ (.A1(net987),
    .A2(\decoded_imm[4] ),
    .B1(net858),
    .X(_05208_));
 sky130_fd_sc_hd__o22a_1 _10513_ (.A1(net1175),
    .A2(net860),
    .B1(_05208_),
    .B2(_03264_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(\cpuregs[6][5] ),
    .A1(\cpuregs[7][5] ),
    .S(net676),
    .X(_05209_));
 sky130_fd_sc_hd__or2_1 _10515_ (.A(\cpuregs[4][5] ),
    .B(net676),
    .X(_05210_));
 sky130_fd_sc_hd__o211a_1 _10516_ (.A1(\cpuregs[5][5] ),
    .A2(net630),
    .B1(net815),
    .C1(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__a211o_1 _10517_ (.A1(net801),
    .A2(_05209_),
    .B1(_05211_),
    .C1(net838),
    .X(_05212_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(\cpuregs[2][5] ),
    .A1(\cpuregs[3][5] ),
    .S(net675),
    .X(_05213_));
 sky130_fd_sc_hd__a221o_1 _10519_ (.A1(\cpuregs[1][5] ),
    .A2(net550),
    .B1(_05213_),
    .B2(net801),
    .C1(net829),
    .X(_05214_));
 sky130_fd_sc_hd__a21o_1 _10520_ (.A1(_05212_),
    .A2(_05214_),
    .B1(net785),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(\cpuregs[14][5] ),
    .A1(\cpuregs[15][5] ),
    .S(net675),
    .X(_05216_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(\cpuregs[12][5] ),
    .A1(\cpuregs[13][5] ),
    .S(net675),
    .X(_05217_));
 sky130_fd_sc_hd__or2_1 _10523_ (.A(net801),
    .B(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__o211a_1 _10524_ (.A1(net815),
    .A2(_05216_),
    .B1(_05218_),
    .C1(net829),
    .X(_05219_));
 sky130_fd_sc_hd__or2_1 _10525_ (.A(\cpuregs[8][5] ),
    .B(net675),
    .X(_05220_));
 sky130_fd_sc_hd__o211a_1 _10526_ (.A1(\cpuregs[9][5] ),
    .A2(net630),
    .B1(net609),
    .C1(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__or2_1 _10527_ (.A(\cpuregs[10][5] ),
    .B(net675),
    .X(_05222_));
 sky130_fd_sc_hd__o211a_1 _10528_ (.A1(\cpuregs[11][5] ),
    .A2(net630),
    .B1(net595),
    .C1(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__o41a_1 _10529_ (.A1(net790),
    .A2(_05219_),
    .A3(_05221_),
    .A4(_05223_),
    .B1(net776),
    .X(_05224_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(\cpuregs[28][5] ),
    .A1(\cpuregs[29][5] ),
    .S(net678),
    .X(_05225_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(\cpuregs[30][5] ),
    .A1(\cpuregs[31][5] ),
    .S(net678),
    .X(_05226_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(_05225_),
    .A1(_05226_),
    .S(net802),
    .X(_05227_));
 sky130_fd_sc_hd__or2_1 _10533_ (.A(\cpuregs[24][5] ),
    .B(net678),
    .X(_05228_));
 sky130_fd_sc_hd__o211a_1 _10534_ (.A1(\cpuregs[25][5] ),
    .A2(net629),
    .B1(net609),
    .C1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__or2_1 _10535_ (.A(\cpuregs[26][5] ),
    .B(net678),
    .X(_05230_));
 sky130_fd_sc_hd__o211a_1 _10536_ (.A1(\cpuregs[27][5] ),
    .A2(net629),
    .B1(net595),
    .C1(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__a2111o_1 _10537_ (.A1(net830),
    .A2(_05227_),
    .B1(_05229_),
    .C1(_05231_),
    .D1(net790),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(\cpuregs[20][5] ),
    .A1(\cpuregs[21][5] ),
    .S(net678),
    .X(_05233_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(\cpuregs[22][5] ),
    .A1(\cpuregs[23][5] ),
    .S(net678),
    .X(_05234_));
 sky130_fd_sc_hd__mux2_1 _10540_ (.A0(_05233_),
    .A1(_05234_),
    .S(net802),
    .X(_05235_));
 sky130_fd_sc_hd__or2_1 _10541_ (.A(\cpuregs[16][5] ),
    .B(net676),
    .X(_05236_));
 sky130_fd_sc_hd__o211a_1 _10542_ (.A1(\cpuregs[17][5] ),
    .A2(net629),
    .B1(net609),
    .C1(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__o21a_1 _10543_ (.A1(\cpuregs[19][5] ),
    .A2(net631),
    .B1(net595),
    .X(_05238_));
 sky130_fd_sc_hd__o22a_1 _10544_ (.A1(\cpuregs[18][5] ),
    .A2(net552),
    .B1(_05238_),
    .B2(net781),
    .X(_05239_));
 sky130_fd_sc_hd__a211o_1 _10545_ (.A1(net829),
    .A2(_05235_),
    .B1(_05237_),
    .C1(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__and3_1 _10546_ (.A(net772),
    .B(_05232_),
    .C(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__a21oi_2 _10547_ (.A1(_05215_),
    .A2(_05224_),
    .B1(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__or2_1 _10548_ (.A(net1078),
    .B(\decoded_imm[5] ),
    .X(_05243_));
 sky130_fd_sc_hd__a21oi_1 _10549_ (.A1(net1078),
    .A2(_05242_),
    .B1(net855),
    .Y(_05244_));
 sky130_fd_sc_hd__a22o_1 _10550_ (.A1(net1172),
    .A2(net855),
    .B1(_05243_),
    .B2(_05244_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(\cpuregs[6][6] ),
    .A1(\cpuregs[7][6] ),
    .S(net677),
    .X(_05245_));
 sky130_fd_sc_hd__or2_1 _10552_ (.A(\cpuregs[4][6] ),
    .B(net677),
    .X(_05246_));
 sky130_fd_sc_hd__o211a_1 _10553_ (.A1(\cpuregs[5][6] ),
    .A2(net629),
    .B1(net815),
    .C1(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__a211o_1 _10554_ (.A1(net801),
    .A2(_05245_),
    .B1(_05247_),
    .C1(net839),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(\cpuregs[2][6] ),
    .A1(\cpuregs[3][6] ),
    .S(net674),
    .X(_05249_));
 sky130_fd_sc_hd__a221o_1 _10556_ (.A1(\cpuregs[1][6] ),
    .A2(net549),
    .B1(_05249_),
    .B2(net802),
    .C1(net830),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_1 _10557_ (.A1(_05248_),
    .A2(_05250_),
    .B1(net781),
    .X(_05251_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(\cpuregs[14][6] ),
    .A1(\cpuregs[15][6] ),
    .S(net673),
    .X(_05252_));
 sky130_fd_sc_hd__mux2_1 _10559_ (.A0(\cpuregs[12][6] ),
    .A1(\cpuregs[13][6] ),
    .S(net673),
    .X(_05253_));
 sky130_fd_sc_hd__or2_1 _10560_ (.A(net801),
    .B(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__o211a_1 _10561_ (.A1(net815),
    .A2(_05252_),
    .B1(_05254_),
    .C1(net829),
    .X(_05255_));
 sky130_fd_sc_hd__or2_1 _10562_ (.A(\cpuregs[8][6] ),
    .B(net674),
    .X(_05256_));
 sky130_fd_sc_hd__o211a_1 _10563_ (.A1(\cpuregs[9][6] ),
    .A2(net629),
    .B1(net609),
    .C1(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__or2_1 _10564_ (.A(\cpuregs[10][6] ),
    .B(net674),
    .X(_05258_));
 sky130_fd_sc_hd__o211a_1 _10565_ (.A1(\cpuregs[11][6] ),
    .A2(net629),
    .B1(net596),
    .C1(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__o41a_1 _10566_ (.A1(net789),
    .A2(_05255_),
    .A3(_05257_),
    .A4(_05259_),
    .B1(net777),
    .X(_05260_));
 sky130_fd_sc_hd__mux2_1 _10567_ (.A0(\cpuregs[28][6] ),
    .A1(\cpuregs[29][6] ),
    .S(net670),
    .X(_05261_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(\cpuregs[30][6] ),
    .A1(\cpuregs[31][6] ),
    .S(net670),
    .X(_05262_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(_05261_),
    .A1(_05262_),
    .S(net800),
    .X(_05263_));
 sky130_fd_sc_hd__or2_1 _10570_ (.A(\cpuregs[24][6] ),
    .B(net677),
    .X(_05264_));
 sky130_fd_sc_hd__o211a_1 _10571_ (.A1(\cpuregs[25][6] ),
    .A2(net629),
    .B1(net609),
    .C1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__or2_1 _10572_ (.A(\cpuregs[26][6] ),
    .B(net677),
    .X(_05266_));
 sky130_fd_sc_hd__o211a_1 _10573_ (.A1(\cpuregs[27][6] ),
    .A2(net629),
    .B1(net595),
    .C1(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__a2111o_1 _10574_ (.A1(net830),
    .A2(_05263_),
    .B1(_05265_),
    .C1(_05267_),
    .D1(net790),
    .X(_05268_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(\cpuregs[22][6] ),
    .A1(\cpuregs[23][6] ),
    .S(net671),
    .X(_05269_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(\cpuregs[20][6] ),
    .A1(\cpuregs[21][6] ),
    .S(net670),
    .X(_05270_));
 sky130_fd_sc_hd__mux2_1 _10577_ (.A0(_05269_),
    .A1(_05270_),
    .S(net814),
    .X(_05271_));
 sky130_fd_sc_hd__or2_1 _10578_ (.A(\cpuregs[16][6] ),
    .B(net671),
    .X(_05272_));
 sky130_fd_sc_hd__o211a_1 _10579_ (.A1(\cpuregs[17][6] ),
    .A2(net627),
    .B1(net608),
    .C1(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__o21a_1 _10580_ (.A1(\cpuregs[19][6] ),
    .A2(net627),
    .B1(net594),
    .X(_05274_));
 sky130_fd_sc_hd__o22a_1 _10581_ (.A1(\cpuregs[18][6] ),
    .A2(net553),
    .B1(_05274_),
    .B2(net780),
    .X(_05275_));
 sky130_fd_sc_hd__a211o_1 _10582_ (.A1(net827),
    .A2(_05271_),
    .B1(_05273_),
    .C1(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__and3_1 _10583_ (.A(net773),
    .B(_05268_),
    .C(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__a21oi_2 _10584_ (.A1(_05251_),
    .A2(_05260_),
    .B1(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__nand2_1 _10585_ (.A(net1077),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__o21a_1 _10586_ (.A1(net1077),
    .A2(\decoded_imm[6] ),
    .B1(net860),
    .X(_05280_));
 sky130_fd_sc_hd__a22o_1 _10587_ (.A1(net1171),
    .A2(net855),
    .B1(_05279_),
    .B2(_05280_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\cpuregs[6][7] ),
    .A1(\cpuregs[7][7] ),
    .S(net673),
    .X(_05281_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(\cpuregs[4][7] ),
    .A1(\cpuregs[5][7] ),
    .S(net659),
    .X(_05282_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(_05281_),
    .A1(_05282_),
    .S(net815),
    .X(_05283_));
 sky130_fd_sc_hd__or2_1 _10591_ (.A(\cpuregs[0][7] ),
    .B(net673),
    .X(_05284_));
 sky130_fd_sc_hd__o211a_1 _10592_ (.A1(\cpuregs[1][7] ),
    .A2(net630),
    .B1(net609),
    .C1(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__or2_1 _10593_ (.A(\cpuregs[2][7] ),
    .B(net673),
    .X(_05286_));
 sky130_fd_sc_hd__o211a_1 _10594_ (.A1(\cpuregs[3][7] ),
    .A2(net630),
    .B1(net595),
    .C1(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__a211o_1 _10595_ (.A1(net829),
    .A2(_05283_),
    .B1(_05287_),
    .C1(net781),
    .X(_05288_));
 sky130_fd_sc_hd__mux2_1 _10596_ (.A0(\cpuregs[12][7] ),
    .A1(\cpuregs[13][7] ),
    .S(net673),
    .X(_05289_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(\cpuregs[14][7] ),
    .A1(\cpuregs[15][7] ),
    .S(net673),
    .X(_05290_));
 sky130_fd_sc_hd__or2_1 _10598_ (.A(net815),
    .B(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__o211a_1 _10599_ (.A1(net801),
    .A2(_05289_),
    .B1(_05291_),
    .C1(net829),
    .X(_05292_));
 sky130_fd_sc_hd__or2_1 _10600_ (.A(\cpuregs[8][7] ),
    .B(net673),
    .X(_05293_));
 sky130_fd_sc_hd__o211a_1 _10601_ (.A1(\cpuregs[9][7] ),
    .A2(net630),
    .B1(net609),
    .C1(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__or2_1 _10602_ (.A(\cpuregs[10][7] ),
    .B(net673),
    .X(_05295_));
 sky130_fd_sc_hd__o211a_1 _10603_ (.A1(\cpuregs[11][7] ),
    .A2(net630),
    .B1(net595),
    .C1(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__or4_1 _10604_ (.A(net790),
    .B(_05292_),
    .C(_05294_),
    .D(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__o21a_1 _10605_ (.A1(_05285_),
    .A2(_05288_),
    .B1(_03171_),
    .X(_05298_));
 sky130_fd_sc_hd__mux2_1 _10606_ (.A0(\cpuregs[22][7] ),
    .A1(\cpuregs[23][7] ),
    .S(net668),
    .X(_05299_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(\cpuregs[20][7] ),
    .A1(\cpuregs[21][7] ),
    .S(net668),
    .X(_05300_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(_05299_),
    .A1(_05300_),
    .S(net814),
    .X(_05301_));
 sky130_fd_sc_hd__or2_1 _10609_ (.A(\cpuregs[16][7] ),
    .B(net665),
    .X(_05302_));
 sky130_fd_sc_hd__o211a_1 _10610_ (.A1(\cpuregs[17][7] ),
    .A2(net626),
    .B1(net608),
    .C1(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__o21a_1 _10611_ (.A1(\cpuregs[19][7] ),
    .A2(net626),
    .B1(net593),
    .X(_05304_));
 sky130_fd_sc_hd__o22a_1 _10612_ (.A1(\cpuregs[18][7] ),
    .A2(net553),
    .B1(_05304_),
    .B2(net780),
    .X(_05305_));
 sky130_fd_sc_hd__a211o_1 _10613_ (.A1(net827),
    .A2(_05301_),
    .B1(_05303_),
    .C1(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__mux2_1 _10614_ (.A0(\cpuregs[30][7] ),
    .A1(\cpuregs[31][7] ),
    .S(net669),
    .X(_05307_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\cpuregs[28][7] ),
    .A1(\cpuregs[29][7] ),
    .S(net669),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(_05307_),
    .A1(_05308_),
    .S(net814),
    .X(_05309_));
 sky130_fd_sc_hd__or2_1 _10617_ (.A(\cpuregs[24][7] ),
    .B(net669),
    .X(_05310_));
 sky130_fd_sc_hd__o211a_1 _10618_ (.A1(\cpuregs[25][7] ),
    .A2(net626),
    .B1(net608),
    .C1(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__or2_1 _10619_ (.A(\cpuregs[26][7] ),
    .B(net668),
    .X(_05312_));
 sky130_fd_sc_hd__o211a_1 _10620_ (.A1(\cpuregs[27][7] ),
    .A2(net626),
    .B1(net594),
    .C1(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__a2111o_1 _10621_ (.A1(net827),
    .A2(_05309_),
    .B1(_05311_),
    .C1(_05313_),
    .D1(net789),
    .X(_05314_));
 sky130_fd_sc_hd__and3_1 _10622_ (.A(net773),
    .B(_05306_),
    .C(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__a21oi_2 _10623_ (.A1(_05297_),
    .A2(_05298_),
    .B1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_1 _10624_ (.A(net1077),
    .B(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__o21a_1 _10625_ (.A1(net1077),
    .A2(\decoded_imm[7] ),
    .B1(net860),
    .X(_05318_));
 sky130_fd_sc_hd__a22o_1 _10626_ (.A1(net1169),
    .A2(net854),
    .B1(_05317_),
    .B2(_05318_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(\cpuregs[6][8] ),
    .A1(\cpuregs[7][8] ),
    .S(net677),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\cpuregs[4][8] ),
    .A1(\cpuregs[5][8] ),
    .S(net677),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _10629_ (.A0(_05319_),
    .A1(_05320_),
    .S(net815),
    .X(_05321_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\cpuregs[2][8] ),
    .A1(\cpuregs[3][8] ),
    .S(net674),
    .X(_05322_));
 sky130_fd_sc_hd__a221o_1 _10631_ (.A1(\cpuregs[1][8] ),
    .A2(net550),
    .B1(_05322_),
    .B2(net800),
    .C1(net827),
    .X(_05323_));
 sky130_fd_sc_hd__o21a_1 _10632_ (.A1(net838),
    .A2(_05321_),
    .B1(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__mux2_1 _10633_ (.A0(\cpuregs[12][8] ),
    .A1(\cpuregs[13][8] ),
    .S(net665),
    .X(_05325_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(\cpuregs[14][8] ),
    .A1(\cpuregs[15][8] ),
    .S(net664),
    .X(_05326_));
 sky130_fd_sc_hd__or2_1 _10635_ (.A(net813),
    .B(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__o211a_1 _10636_ (.A1(net800),
    .A2(_05325_),
    .B1(_05327_),
    .C1(net827),
    .X(_05328_));
 sky130_fd_sc_hd__or2_1 _10637_ (.A(\cpuregs[8][8] ),
    .B(net667),
    .X(_05329_));
 sky130_fd_sc_hd__o211a_1 _10638_ (.A1(\cpuregs[9][8] ),
    .A2(net628),
    .B1(net608),
    .C1(_05329_),
    .X(_05330_));
 sky130_fd_sc_hd__or2_1 _10639_ (.A(\cpuregs[10][8] ),
    .B(net666),
    .X(_05331_));
 sky130_fd_sc_hd__o211a_1 _10640_ (.A1(\cpuregs[11][8] ),
    .A2(net626),
    .B1(net593),
    .C1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__or4_1 _10641_ (.A(net789),
    .B(_05328_),
    .C(_05330_),
    .D(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__o211a_1 _10642_ (.A1(net781),
    .A2(_05324_),
    .B1(_05333_),
    .C1(net777),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\cpuregs[30][8] ),
    .A1(\cpuregs[31][8] ),
    .S(net670),
    .X(_05335_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(\cpuregs[28][8] ),
    .A1(\cpuregs[29][8] ),
    .S(net670),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(_05335_),
    .A1(_05336_),
    .S(net814),
    .X(_05337_));
 sky130_fd_sc_hd__or2_1 _10646_ (.A(\cpuregs[24][8] ),
    .B(net670),
    .X(_05338_));
 sky130_fd_sc_hd__o211a_1 _10647_ (.A1(\cpuregs[25][8] ),
    .A2(net627),
    .B1(net608),
    .C1(_05338_),
    .X(_05339_));
 sky130_fd_sc_hd__or2_1 _10648_ (.A(\cpuregs[26][8] ),
    .B(net670),
    .X(_05340_));
 sky130_fd_sc_hd__o211a_1 _10649_ (.A1(\cpuregs[27][8] ),
    .A2(net626),
    .B1(net594),
    .C1(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__a2111o_1 _10650_ (.A1(net827),
    .A2(_05337_),
    .B1(_05339_),
    .C1(_05341_),
    .D1(net789),
    .X(_05342_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\cpuregs[22][8] ),
    .A1(\cpuregs[23][8] ),
    .S(net668),
    .X(_05343_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(\cpuregs[20][8] ),
    .A1(\cpuregs[21][8] ),
    .S(net669),
    .X(_05344_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(_05343_),
    .A1(_05344_),
    .S(net814),
    .X(_05345_));
 sky130_fd_sc_hd__or2_1 _10654_ (.A(\cpuregs[16][8] ),
    .B(net668),
    .X(_05346_));
 sky130_fd_sc_hd__o211a_1 _10655_ (.A1(\cpuregs[17][8] ),
    .A2(net626),
    .B1(net607),
    .C1(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__o21a_1 _10656_ (.A1(\cpuregs[19][8] ),
    .A2(net626),
    .B1(net594),
    .X(_05348_));
 sky130_fd_sc_hd__o22a_1 _10657_ (.A1(\cpuregs[18][8] ),
    .A2(net553),
    .B1(_05348_),
    .B2(net780),
    .X(_05349_));
 sky130_fd_sc_hd__a211o_1 _10658_ (.A1(net827),
    .A2(_05345_),
    .B1(_05347_),
    .C1(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__a31oi_4 _10659_ (.A1(net773),
    .A2(_05342_),
    .A3(_05350_),
    .B1(_05334_),
    .Y(_05351_));
 sky130_fd_sc_hd__or2_1 _10660_ (.A(net1076),
    .B(\decoded_imm[8] ),
    .X(_05352_));
 sky130_fd_sc_hd__a21oi_1 _10661_ (.A1(net1076),
    .A2(_05351_),
    .B1(net853),
    .Y(_05353_));
 sky130_fd_sc_hd__a22o_1 _10662_ (.A1(net1168),
    .A2(net853),
    .B1(_05352_),
    .B2(_05353_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _10663_ (.A0(\cpuregs[6][9] ),
    .A1(\cpuregs[7][9] ),
    .S(net671),
    .X(_05354_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\cpuregs[4][9] ),
    .A1(\cpuregs[5][9] ),
    .S(net666),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _10665_ (.A0(_05354_),
    .A1(_05355_),
    .S(net813),
    .X(_05356_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\cpuregs[2][9] ),
    .A1(\cpuregs[3][9] ),
    .S(net667),
    .X(_05357_));
 sky130_fd_sc_hd__a221o_1 _10667_ (.A1(\cpuregs[1][9] ),
    .A2(net550),
    .B1(_05357_),
    .B2(net800),
    .C1(net828),
    .X(_05358_));
 sky130_fd_sc_hd__o21a_1 _10668_ (.A1(net839),
    .A2(_05356_),
    .B1(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__mux2_1 _10669_ (.A0(\cpuregs[14][9] ),
    .A1(\cpuregs[15][9] ),
    .S(net667),
    .X(_05360_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\cpuregs[12][9] ),
    .A1(\cpuregs[13][9] ),
    .S(net667),
    .X(_05361_));
 sky130_fd_sc_hd__or2_1 _10671_ (.A(net800),
    .B(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__o211a_1 _10672_ (.A1(net813),
    .A2(_05360_),
    .B1(_05362_),
    .C1(net828),
    .X(_05363_));
 sky130_fd_sc_hd__or2_1 _10673_ (.A(\cpuregs[8][9] ),
    .B(net667),
    .X(_05364_));
 sky130_fd_sc_hd__o211a_1 _10674_ (.A1(\cpuregs[9][9] ),
    .A2(net628),
    .B1(net607),
    .C1(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__or2_1 _10675_ (.A(\cpuregs[10][9] ),
    .B(net667),
    .X(_05366_));
 sky130_fd_sc_hd__o211a_1 _10676_ (.A1(\cpuregs[11][9] ),
    .A2(net628),
    .B1(net593),
    .C1(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__or4_1 _10677_ (.A(net789),
    .B(_05363_),
    .C(_05365_),
    .D(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__o211a_1 _10678_ (.A1(net780),
    .A2(_05359_),
    .B1(_05368_),
    .C1(net777),
    .X(_05369_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(\cpuregs[30][9] ),
    .A1(\cpuregs[31][9] ),
    .S(net670),
    .X(_05370_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\cpuregs[28][9] ),
    .A1(\cpuregs[29][9] ),
    .S(net670),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(_05370_),
    .A1(_05371_),
    .S(net814),
    .X(_05372_));
 sky130_fd_sc_hd__or2_1 _10682_ (.A(\cpuregs[24][9] ),
    .B(net671),
    .X(_05373_));
 sky130_fd_sc_hd__o211a_1 _10683_ (.A1(\cpuregs[25][9] ),
    .A2(net627),
    .B1(net608),
    .C1(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__or2_1 _10684_ (.A(\cpuregs[26][9] ),
    .B(net670),
    .X(_05375_));
 sky130_fd_sc_hd__o211a_1 _10685_ (.A1(\cpuregs[27][9] ),
    .A2(net627),
    .B1(net594),
    .C1(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__a2111o_1 _10686_ (.A1(net830),
    .A2(_05372_),
    .B1(_05374_),
    .C1(_05376_),
    .D1(net789),
    .X(_05377_));
 sky130_fd_sc_hd__mux2_1 _10687_ (.A0(\cpuregs[20][9] ),
    .A1(\cpuregs[21][9] ),
    .S(net671),
    .X(_05378_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(\cpuregs[22][9] ),
    .A1(\cpuregs[23][9] ),
    .S(net671),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(_05378_),
    .A1(_05379_),
    .S(net800),
    .X(_05380_));
 sky130_fd_sc_hd__or2_1 _10690_ (.A(\cpuregs[16][9] ),
    .B(net671),
    .X(_05381_));
 sky130_fd_sc_hd__o211a_1 _10691_ (.A1(\cpuregs[17][9] ),
    .A2(net627),
    .B1(net607),
    .C1(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__o21a_1 _10692_ (.A1(\cpuregs[19][9] ),
    .A2(net627),
    .B1(net594),
    .X(_05383_));
 sky130_fd_sc_hd__o22a_1 _10693_ (.A1(\cpuregs[18][9] ),
    .A2(net553),
    .B1(_05383_),
    .B2(net780),
    .X(_05384_));
 sky130_fd_sc_hd__a211o_1 _10694_ (.A1(net827),
    .A2(_05380_),
    .B1(_05382_),
    .C1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__a31oi_4 _10695_ (.A1(net773),
    .A2(_05377_),
    .A3(_05385_),
    .B1(_05369_),
    .Y(_05386_));
 sky130_fd_sc_hd__or2_1 _10696_ (.A(net1076),
    .B(\decoded_imm[9] ),
    .X(_05387_));
 sky130_fd_sc_hd__a21oi_1 _10697_ (.A1(net1076),
    .A2(_05386_),
    .B1(net853),
    .Y(_05388_));
 sky130_fd_sc_hd__a22o_1 _10698_ (.A1(net1167),
    .A2(net853),
    .B1(_05387_),
    .B2(_05388_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(\cpuregs[6][10] ),
    .A1(\cpuregs[7][10] ),
    .S(net666),
    .X(_05389_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(\cpuregs[4][10] ),
    .A1(\cpuregs[5][10] ),
    .S(net666),
    .X(_05390_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(_05389_),
    .A1(_05390_),
    .S(net813),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(\cpuregs[2][10] ),
    .A1(\cpuregs[3][10] ),
    .S(net673),
    .X(_05392_));
 sky130_fd_sc_hd__a221o_1 _10703_ (.A1(\cpuregs[1][10] ),
    .A2(net550),
    .B1(_05392_),
    .B2(net800),
    .C1(net828),
    .X(_05393_));
 sky130_fd_sc_hd__o21a_1 _10704_ (.A1(net839),
    .A2(_05391_),
    .B1(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__mux2_1 _10705_ (.A0(\cpuregs[14][10] ),
    .A1(\cpuregs[15][10] ),
    .S(net664),
    .X(_05395_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(\cpuregs[12][10] ),
    .A1(\cpuregs[13][10] ),
    .S(net664),
    .X(_05396_));
 sky130_fd_sc_hd__or2_1 _10707_ (.A(net800),
    .B(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__o211a_1 _10708_ (.A1(net813),
    .A2(_05395_),
    .B1(_05397_),
    .C1(net828),
    .X(_05398_));
 sky130_fd_sc_hd__or2_1 _10709_ (.A(\cpuregs[8][10] ),
    .B(net666),
    .X(_05399_));
 sky130_fd_sc_hd__o211a_1 _10710_ (.A1(\cpuregs[9][10] ),
    .A2(net628),
    .B1(net607),
    .C1(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__or2_1 _10711_ (.A(\cpuregs[10][10] ),
    .B(net666),
    .X(_05401_));
 sky130_fd_sc_hd__o211a_1 _10712_ (.A1(\cpuregs[11][10] ),
    .A2(net625),
    .B1(net593),
    .C1(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__or4_1 _10713_ (.A(net789),
    .B(_05398_),
    .C(_05400_),
    .D(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__o211a_1 _10714_ (.A1(net780),
    .A2(_05394_),
    .B1(_05403_),
    .C1(net777),
    .X(_05404_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(\cpuregs[28][10] ),
    .A1(\cpuregs[29][10] ),
    .S(net669),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\cpuregs[30][10] ),
    .A1(\cpuregs[31][10] ),
    .S(net669),
    .X(_05406_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(_05405_),
    .A1(_05406_),
    .S(net802),
    .X(_05407_));
 sky130_fd_sc_hd__or2_1 _10718_ (.A(\cpuregs[24][10] ),
    .B(net668),
    .X(_05408_));
 sky130_fd_sc_hd__o211a_1 _10719_ (.A1(\cpuregs[25][10] ),
    .A2(net627),
    .B1(net608),
    .C1(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__or2_1 _10720_ (.A(\cpuregs[26][10] ),
    .B(net668),
    .X(_05410_));
 sky130_fd_sc_hd__o211a_1 _10721_ (.A1(\cpuregs[27][10] ),
    .A2(net627),
    .B1(net594),
    .C1(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__a2111o_1 _10722_ (.A1(net827),
    .A2(_05407_),
    .B1(_05409_),
    .C1(_05411_),
    .D1(net789),
    .X(_05412_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(\cpuregs[22][10] ),
    .A1(\cpuregs[23][10] ),
    .S(net668),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(\cpuregs[20][10] ),
    .A1(\cpuregs[21][10] ),
    .S(net668),
    .X(_05414_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(_05413_),
    .A1(_05414_),
    .S(net814),
    .X(_05415_));
 sky130_fd_sc_hd__or2_1 _10726_ (.A(\cpuregs[16][10] ),
    .B(net668),
    .X(_05416_));
 sky130_fd_sc_hd__o211a_1 _10727_ (.A1(\cpuregs[17][10] ),
    .A2(net626),
    .B1(net607),
    .C1(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__o21a_1 _10728_ (.A1(\cpuregs[19][10] ),
    .A2(net626),
    .B1(net593),
    .X(_05418_));
 sky130_fd_sc_hd__o22a_1 _10729_ (.A1(\cpuregs[18][10] ),
    .A2(net553),
    .B1(_05418_),
    .B2(net780),
    .X(_05419_));
 sky130_fd_sc_hd__a211o_1 _10730_ (.A1(net827),
    .A2(_05415_),
    .B1(_05417_),
    .C1(_05419_),
    .X(_05420_));
 sky130_fd_sc_hd__a31oi_4 _10731_ (.A1(net773),
    .A2(_05412_),
    .A3(_05420_),
    .B1(_05404_),
    .Y(_05421_));
 sky130_fd_sc_hd__or2_1 _10732_ (.A(net1076),
    .B(\decoded_imm[10] ),
    .X(_05422_));
 sky130_fd_sc_hd__a21oi_1 _10733_ (.A1(net1076),
    .A2(_05421_),
    .B1(net853),
    .Y(_05423_));
 sky130_fd_sc_hd__a22o_1 _10734_ (.A1(net1166),
    .A2(net853),
    .B1(_05422_),
    .B2(_05423_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _10735_ (.A0(\cpuregs[28][11] ),
    .A1(\cpuregs[29][11] ),
    .S(net665),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\cpuregs[30][11] ),
    .A1(\cpuregs[31][11] ),
    .S(net665),
    .X(_05425_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(_05424_),
    .A1(_05425_),
    .S(net800),
    .X(_05426_));
 sky130_fd_sc_hd__or2_1 _10738_ (.A(\cpuregs[24][11] ),
    .B(net664),
    .X(_05427_));
 sky130_fd_sc_hd__o211a_1 _10739_ (.A1(\cpuregs[25][11] ),
    .A2(net625),
    .B1(net607),
    .C1(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__or2_1 _10740_ (.A(\cpuregs[26][11] ),
    .B(net665),
    .X(_05429_));
 sky130_fd_sc_hd__o211a_1 _10741_ (.A1(\cpuregs[27][11] ),
    .A2(net625),
    .B1(net593),
    .C1(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__a2111o_1 _10742_ (.A1(net828),
    .A2(_05426_),
    .B1(_05428_),
    .C1(_05430_),
    .D1(net789),
    .X(_05431_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\cpuregs[22][11] ),
    .A1(\cpuregs[23][11] ),
    .S(net664),
    .X(_05432_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(\cpuregs[20][11] ),
    .A1(\cpuregs[21][11] ),
    .S(net665),
    .X(_05433_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(_05432_),
    .A1(_05433_),
    .S(net813),
    .X(_05434_));
 sky130_fd_sc_hd__or2_1 _10746_ (.A(\cpuregs[16][11] ),
    .B(net665),
    .X(_05435_));
 sky130_fd_sc_hd__o211a_1 _10747_ (.A1(\cpuregs[17][11] ),
    .A2(net625),
    .B1(net607),
    .C1(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__o21a_1 _10748_ (.A1(\cpuregs[19][11] ),
    .A2(net625),
    .B1(net593),
    .X(_05437_));
 sky130_fd_sc_hd__o22a_1 _10749_ (.A1(\cpuregs[18][11] ),
    .A2(net553),
    .B1(_05437_),
    .B2(net780),
    .X(_05438_));
 sky130_fd_sc_hd__a211o_1 _10750_ (.A1(net828),
    .A2(_05434_),
    .B1(_05436_),
    .C1(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(\cpuregs[6][11] ),
    .A1(\cpuregs[7][11] ),
    .S(net666),
    .X(_05440_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\cpuregs[4][11] ),
    .A1(\cpuregs[5][11] ),
    .S(net666),
    .X(_05441_));
 sky130_fd_sc_hd__mux2_1 _10753_ (.A0(_05440_),
    .A1(_05441_),
    .S(net813),
    .X(_05442_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\cpuregs[2][11] ),
    .A1(\cpuregs[3][11] ),
    .S(net653),
    .X(_05443_));
 sky130_fd_sc_hd__a221o_1 _10755_ (.A1(\cpuregs[1][11] ),
    .A2(net549),
    .B1(_05443_),
    .B2(net796),
    .C1(net823),
    .X(_05444_));
 sky130_fd_sc_hd__o21a_1 _10756_ (.A1(net839),
    .A2(_05442_),
    .B1(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__mux2_1 _10757_ (.A0(\cpuregs[14][11] ),
    .A1(\cpuregs[15][11] ),
    .S(net666),
    .X(_05446_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\cpuregs[12][11] ),
    .A1(\cpuregs[13][11] ),
    .S(net651),
    .X(_05447_));
 sky130_fd_sc_hd__or2_1 _10759_ (.A(net800),
    .B(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__o211a_1 _10760_ (.A1(net813),
    .A2(_05446_),
    .B1(_05448_),
    .C1(net828),
    .X(_05449_));
 sky130_fd_sc_hd__or2_1 _10761_ (.A(\cpuregs[8][11] ),
    .B(net666),
    .X(_05450_));
 sky130_fd_sc_hd__o211a_1 _10762_ (.A1(\cpuregs[9][11] ),
    .A2(net628),
    .B1(net607),
    .C1(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__or2_1 _10763_ (.A(\cpuregs[10][11] ),
    .B(net653),
    .X(_05452_));
 sky130_fd_sc_hd__o211a_1 _10764_ (.A1(\cpuregs[11][11] ),
    .A2(net625),
    .B1(net593),
    .C1(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__or4_1 _10765_ (.A(net789),
    .B(_05449_),
    .C(_05451_),
    .D(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__o211a_1 _10766_ (.A1(net780),
    .A2(_05445_),
    .B1(_05454_),
    .C1(net777),
    .X(_05455_));
 sky130_fd_sc_hd__a31oi_4 _10767_ (.A1(net773),
    .A2(_05431_),
    .A3(_05439_),
    .B1(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__nand2_1 _10768_ (.A(net1076),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__o21a_1 _10769_ (.A1(net1076),
    .A2(\decoded_imm[11] ),
    .B1(net860),
    .X(_05458_));
 sky130_fd_sc_hd__a22o_1 _10770_ (.A1(net1165),
    .A2(net853),
    .B1(_05457_),
    .B2(_05458_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(\cpuregs[28][12] ),
    .A1(\cpuregs[29][12] ),
    .S(net650),
    .X(_05459_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(\cpuregs[30][12] ),
    .A1(\cpuregs[31][12] ),
    .S(net650),
    .X(_05460_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(_05459_),
    .A1(_05460_),
    .S(net797),
    .X(_05461_));
 sky130_fd_sc_hd__or2_1 _10774_ (.A(\cpuregs[24][12] ),
    .B(net650),
    .X(_05462_));
 sky130_fd_sc_hd__o211a_1 _10775_ (.A1(\cpuregs[25][12] ),
    .A2(net619),
    .B1(net604),
    .C1(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__or2_1 _10776_ (.A(\cpuregs[26][12] ),
    .B(net650),
    .X(_05464_));
 sky130_fd_sc_hd__o211a_1 _10777_ (.A1(\cpuregs[27][12] ),
    .A2(net619),
    .B1(net590),
    .C1(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__a2111o_1 _10778_ (.A1(net826),
    .A2(_05461_),
    .B1(_05463_),
    .C1(_05465_),
    .D1(net787),
    .X(_05466_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\cpuregs[22][12] ),
    .A1(\cpuregs[23][12] ),
    .S(net650),
    .X(_05467_));
 sky130_fd_sc_hd__mux2_1 _10780_ (.A0(\cpuregs[20][12] ),
    .A1(\cpuregs[21][12] ),
    .S(net646),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(_05467_),
    .A1(_05468_),
    .S(net809),
    .X(_05469_));
 sky130_fd_sc_hd__or2_1 _10782_ (.A(\cpuregs[16][12] ),
    .B(net646),
    .X(_05470_));
 sky130_fd_sc_hd__o211a_1 _10783_ (.A1(\cpuregs[17][12] ),
    .A2(net617),
    .B1(net603),
    .C1(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__o21a_1 _10784_ (.A1(\cpuregs[19][12] ),
    .A2(net617),
    .B1(net589),
    .X(_05472_));
 sky130_fd_sc_hd__o22a_1 _10785_ (.A1(\cpuregs[18][12] ),
    .A2(net552),
    .B1(_05472_),
    .B2(net779),
    .X(_05473_));
 sky130_fd_sc_hd__a211o_1 _10786_ (.A1(net822),
    .A2(_05469_),
    .B1(_05471_),
    .C1(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\cpuregs[6][12] ),
    .A1(\cpuregs[7][12] ),
    .S(net652),
    .X(_05475_));
 sky130_fd_sc_hd__mux2_1 _10788_ (.A0(\cpuregs[4][12] ),
    .A1(\cpuregs[5][12] ),
    .S(net652),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(_05475_),
    .A1(_05476_),
    .S(net809),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(\cpuregs[2][12] ),
    .A1(\cpuregs[3][12] ),
    .S(net659),
    .X(_05478_));
 sky130_fd_sc_hd__a221o_1 _10791_ (.A1(\cpuregs[1][12] ),
    .A2(net549),
    .B1(_05478_),
    .B2(net797),
    .C1(net823),
    .X(_05479_));
 sky130_fd_sc_hd__o21a_1 _10792_ (.A1(net838),
    .A2(_05477_),
    .B1(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\cpuregs[14][12] ),
    .A1(\cpuregs[15][12] ),
    .S(net652),
    .X(_05481_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(\cpuregs[12][12] ),
    .A1(\cpuregs[13][12] ),
    .S(net650),
    .X(_05482_));
 sky130_fd_sc_hd__or2_1 _10795_ (.A(net797),
    .B(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__o211a_1 _10796_ (.A1(net812),
    .A2(_05481_),
    .B1(_05483_),
    .C1(net826),
    .X(_05484_));
 sky130_fd_sc_hd__or2_1 _10797_ (.A(\cpuregs[8][12] ),
    .B(net652),
    .X(_05485_));
 sky130_fd_sc_hd__o211a_1 _10798_ (.A1(\cpuregs[9][12] ),
    .A2(net620),
    .B1(net604),
    .C1(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__or2_1 _10799_ (.A(\cpuregs[10][12] ),
    .B(net652),
    .X(_05487_));
 sky130_fd_sc_hd__o211a_1 _10800_ (.A1(\cpuregs[11][12] ),
    .A2(net619),
    .B1(net589),
    .C1(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__or4_1 _10801_ (.A(net787),
    .B(_05484_),
    .C(_05486_),
    .D(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__o211a_1 _10802_ (.A1(net779),
    .A2(_05480_),
    .B1(_05489_),
    .C1(net776),
    .X(_05490_));
 sky130_fd_sc_hd__a31oi_4 _10803_ (.A1(net772),
    .A2(_05466_),
    .A3(_05474_),
    .B1(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__or2_1 _10804_ (.A(net1075),
    .B(\decoded_imm[12] ),
    .X(_05492_));
 sky130_fd_sc_hd__a21oi_1 _10805_ (.A1(net1075),
    .A2(_05491_),
    .B1(net854),
    .Y(_05493_));
 sky130_fd_sc_hd__a22o_1 _10806_ (.A1(net1164),
    .A2(net854),
    .B1(_05492_),
    .B2(_05493_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\cpuregs[6][13] ),
    .A1(\cpuregs[7][13] ),
    .S(net653),
    .X(_05494_));
 sky130_fd_sc_hd__or2_1 _10808_ (.A(\cpuregs[4][13] ),
    .B(net653),
    .X(_05495_));
 sky130_fd_sc_hd__o211a_1 _10809_ (.A1(\cpuregs[5][13] ),
    .A2(net620),
    .B1(net812),
    .C1(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__a211o_1 _10810_ (.A1(net797),
    .A2(_05494_),
    .B1(_05496_),
    .C1(net838),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(\cpuregs[2][13] ),
    .A1(\cpuregs[3][13] ),
    .S(net660),
    .X(_05498_));
 sky130_fd_sc_hd__a221o_1 _10812_ (.A1(\cpuregs[1][13] ),
    .A2(net549),
    .B1(_05498_),
    .B2(net799),
    .C1(net823),
    .X(_05499_));
 sky130_fd_sc_hd__a21o_1 _10813_ (.A1(_05497_),
    .A2(_05499_),
    .B1(net779),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\cpuregs[12][13] ),
    .A1(\cpuregs[13][13] ),
    .S(net651),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\cpuregs[14][13] ),
    .A1(\cpuregs[15][13] ),
    .S(net652),
    .X(_05502_));
 sky130_fd_sc_hd__or2_1 _10816_ (.A(net809),
    .B(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__o211a_1 _10817_ (.A1(net796),
    .A2(_05501_),
    .B1(_05503_),
    .C1(net823),
    .X(_05504_));
 sky130_fd_sc_hd__or2_1 _10818_ (.A(\cpuregs[8][13] ),
    .B(net652),
    .X(_05505_));
 sky130_fd_sc_hd__o211a_1 _10819_ (.A1(\cpuregs[9][13] ),
    .A2(net619),
    .B1(net603),
    .C1(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__or2_1 _10820_ (.A(\cpuregs[10][13] ),
    .B(net652),
    .X(_05507_));
 sky130_fd_sc_hd__o211a_1 _10821_ (.A1(\cpuregs[11][13] ),
    .A2(net619),
    .B1(net590),
    .C1(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__o41a_1 _10822_ (.A1(net788),
    .A2(_05504_),
    .A3(_05506_),
    .A4(_05508_),
    .B1(net776),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\cpuregs[28][13] ),
    .A1(\cpuregs[29][13] ),
    .S(net651),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(\cpuregs[30][13] ),
    .A1(\cpuregs[31][13] ),
    .S(net651),
    .X(_05511_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(_05510_),
    .A1(_05511_),
    .S(net796),
    .X(_05512_));
 sky130_fd_sc_hd__or2_1 _10826_ (.A(\cpuregs[24][13] ),
    .B(net650),
    .X(_05513_));
 sky130_fd_sc_hd__o211a_1 _10827_ (.A1(\cpuregs[25][13] ),
    .A2(net619),
    .B1(net604),
    .C1(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__or2_1 _10828_ (.A(\cpuregs[26][13] ),
    .B(net650),
    .X(_05515_));
 sky130_fd_sc_hd__o211a_1 _10829_ (.A1(\cpuregs[27][13] ),
    .A2(net619),
    .B1(net590),
    .C1(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__a2111o_1 _10830_ (.A1(net823),
    .A2(_05512_),
    .B1(_05514_),
    .C1(_05516_),
    .D1(net787),
    .X(_05517_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\cpuregs[20][13] ),
    .A1(\cpuregs[21][13] ),
    .S(net651),
    .X(_05518_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(\cpuregs[22][13] ),
    .A1(\cpuregs[23][13] ),
    .S(net651),
    .X(_05519_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(_05518_),
    .A1(_05519_),
    .S(net797),
    .X(_05520_));
 sky130_fd_sc_hd__or2_1 _10834_ (.A(\cpuregs[16][13] ),
    .B(net650),
    .X(_05521_));
 sky130_fd_sc_hd__o211a_1 _10835_ (.A1(\cpuregs[17][13] ),
    .A2(net619),
    .B1(net604),
    .C1(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__o21a_1 _10836_ (.A1(\cpuregs[19][13] ),
    .A2(net619),
    .B1(net590),
    .X(_05523_));
 sky130_fd_sc_hd__o22a_1 _10837_ (.A1(\cpuregs[18][13] ),
    .A2(net552),
    .B1(_05523_),
    .B2(net779),
    .X(_05524_));
 sky130_fd_sc_hd__a211o_1 _10838_ (.A1(net823),
    .A2(_05520_),
    .B1(_05522_),
    .C1(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__and3_1 _10839_ (.A(net772),
    .B(_05517_),
    .C(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__a21oi_2 _10840_ (.A1(_05500_),
    .A2(_05509_),
    .B1(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__or2_1 _10841_ (.A(net1075),
    .B(\decoded_imm[13] ),
    .X(_05528_));
 sky130_fd_sc_hd__a21oi_1 _10842_ (.A1(net1075),
    .A2(_05527_),
    .B1(net854),
    .Y(_05529_));
 sky130_fd_sc_hd__a22o_1 _10843_ (.A1(net1163),
    .A2(net854),
    .B1(_05528_),
    .B2(_05529_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(\cpuregs[6][14] ),
    .A1(\cpuregs[7][14] ),
    .S(net660),
    .X(_05530_));
 sky130_fd_sc_hd__or2_1 _10845_ (.A(\cpuregs[4][14] ),
    .B(net660),
    .X(_05531_));
 sky130_fd_sc_hd__o211a_1 _10846_ (.A1(\cpuregs[5][14] ),
    .A2(net623),
    .B1(net811),
    .C1(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__a211o_1 _10847_ (.A1(net799),
    .A2(_05530_),
    .B1(_05532_),
    .C1(net838),
    .X(_05533_));
 sky130_fd_sc_hd__mux2_1 _10848_ (.A0(\cpuregs[2][14] ),
    .A1(\cpuregs[3][14] ),
    .S(net660),
    .X(_05534_));
 sky130_fd_sc_hd__a221o_1 _10849_ (.A1(\cpuregs[1][14] ),
    .A2(net549),
    .B1(_05534_),
    .B2(net799),
    .C1(net826),
    .X(_05535_));
 sky130_fd_sc_hd__a21o_1 _10850_ (.A1(_05533_),
    .A2(_05535_),
    .B1(net781),
    .X(_05536_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\cpuregs[14][14] ),
    .A1(\cpuregs[15][14] ),
    .S(net653),
    .X(_05537_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(\cpuregs[12][14] ),
    .A1(\cpuregs[13][14] ),
    .S(net651),
    .X(_05538_));
 sky130_fd_sc_hd__or2_1 _10853_ (.A(net797),
    .B(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__o211a_1 _10854_ (.A1(net812),
    .A2(_05537_),
    .B1(_05539_),
    .C1(net823),
    .X(_05540_));
 sky130_fd_sc_hd__or2_1 _10855_ (.A(\cpuregs[8][14] ),
    .B(net653),
    .X(_05541_));
 sky130_fd_sc_hd__o211a_1 _10856_ (.A1(\cpuregs[9][14] ),
    .A2(net619),
    .B1(net604),
    .C1(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__or2_1 _10857_ (.A(\cpuregs[10][14] ),
    .B(net653),
    .X(_05543_));
 sky130_fd_sc_hd__o211a_1 _10858_ (.A1(\cpuregs[11][14] ),
    .A2(net620),
    .B1(net590),
    .C1(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__o41a_1 _10859_ (.A1(net787),
    .A2(_05540_),
    .A3(_05542_),
    .A4(_05544_),
    .B1(net777),
    .X(_05545_));
 sky130_fd_sc_hd__mux2_1 _10860_ (.A0(\cpuregs[30][14] ),
    .A1(\cpuregs[31][14] ),
    .S(net664),
    .X(_05546_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(\cpuregs[28][14] ),
    .A1(\cpuregs[29][14] ),
    .S(net664),
    .X(_05547_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(_05546_),
    .A1(_05547_),
    .S(net813),
    .X(_05548_));
 sky130_fd_sc_hd__or2_1 _10863_ (.A(\cpuregs[24][14] ),
    .B(net651),
    .X(_05549_));
 sky130_fd_sc_hd__o211a_1 _10864_ (.A1(\cpuregs[25][14] ),
    .A2(net625),
    .B1(net607),
    .C1(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__or2_1 _10865_ (.A(\cpuregs[26][14] ),
    .B(net664),
    .X(_05551_));
 sky130_fd_sc_hd__o211a_1 _10866_ (.A1(\cpuregs[27][14] ),
    .A2(net625),
    .B1(net593),
    .C1(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__a2111o_1 _10867_ (.A1(net828),
    .A2(_05548_),
    .B1(_05550_),
    .C1(_05552_),
    .D1(net787),
    .X(_05553_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(\cpuregs[22][14] ),
    .A1(\cpuregs[23][14] ),
    .S(net664),
    .X(_05554_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(\cpuregs[20][14] ),
    .A1(\cpuregs[21][14] ),
    .S(net664),
    .X(_05555_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(_05554_),
    .A1(_05555_),
    .S(net813),
    .X(_05556_));
 sky130_fd_sc_hd__or2_1 _10871_ (.A(\cpuregs[16][14] ),
    .B(net650),
    .X(_05557_));
 sky130_fd_sc_hd__o211a_1 _10872_ (.A1(\cpuregs[17][14] ),
    .A2(net625),
    .B1(net607),
    .C1(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__o21a_1 _10873_ (.A1(\cpuregs[19][14] ),
    .A2(net625),
    .B1(net593),
    .X(_05559_));
 sky130_fd_sc_hd__o22a_1 _10874_ (.A1(\cpuregs[18][14] ),
    .A2(net553),
    .B1(_05559_),
    .B2(net780),
    .X(_05560_));
 sky130_fd_sc_hd__a211o_1 _10875_ (.A1(net828),
    .A2(_05556_),
    .B1(_05558_),
    .C1(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__and3_1 _10876_ (.A(net772),
    .B(_05553_),
    .C(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__a21oi_2 _10877_ (.A1(_05536_),
    .A2(_05545_),
    .B1(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__or2_1 _10878_ (.A(net1075),
    .B(\decoded_imm[14] ),
    .X(_05564_));
 sky130_fd_sc_hd__a21oi_1 _10879_ (.A1(net1076),
    .A2(_05563_),
    .B1(net853),
    .Y(_05565_));
 sky130_fd_sc_hd__a22o_1 _10880_ (.A1(net240),
    .A2(net855),
    .B1(_05564_),
    .B2(_05565_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(\cpuregs[6][15] ),
    .A1(\cpuregs[7][15] ),
    .S(net659),
    .X(_05566_));
 sky130_fd_sc_hd__or2_1 _10882_ (.A(\cpuregs[4][15] ),
    .B(net659),
    .X(_05567_));
 sky130_fd_sc_hd__o211a_1 _10883_ (.A1(\cpuregs[5][15] ),
    .A2(net621),
    .B1(net811),
    .C1(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__a211o_1 _10884_ (.A1(net799),
    .A2(_05566_),
    .B1(_05568_),
    .C1(net838),
    .X(_05569_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(\cpuregs[2][15] ),
    .A1(\cpuregs[3][15] ),
    .S(net656),
    .X(_05570_));
 sky130_fd_sc_hd__a221o_1 _10886_ (.A1(\cpuregs[1][15] ),
    .A2(net549),
    .B1(_05570_),
    .B2(net798),
    .C1(net822),
    .X(_05571_));
 sky130_fd_sc_hd__a21o_1 _10887_ (.A1(_05569_),
    .A2(_05571_),
    .B1(net782),
    .X(_05572_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(\cpuregs[12][15] ),
    .A1(\cpuregs[13][15] ),
    .S(net647),
    .X(_05573_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\cpuregs[14][15] ),
    .A1(\cpuregs[15][15] ),
    .S(net647),
    .X(_05574_));
 sky130_fd_sc_hd__or2_1 _10890_ (.A(net809),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__o211a_1 _10891_ (.A1(net796),
    .A2(_05573_),
    .B1(_05575_),
    .C1(net822),
    .X(_05576_));
 sky130_fd_sc_hd__or2_1 _10892_ (.A(\cpuregs[8][15] ),
    .B(net648),
    .X(_05577_));
 sky130_fd_sc_hd__o211a_1 _10893_ (.A1(\cpuregs[9][15] ),
    .A2(net618),
    .B1(net603),
    .C1(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__or2_1 _10894_ (.A(\cpuregs[10][15] ),
    .B(net647),
    .X(_05579_));
 sky130_fd_sc_hd__o211a_1 _10895_ (.A1(\cpuregs[11][15] ),
    .A2(net618),
    .B1(net589),
    .C1(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__o41a_1 _10896_ (.A1(net787),
    .A2(_05576_),
    .A3(_05578_),
    .A4(_05580_),
    .B1(net776),
    .X(_05581_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\cpuregs[28][15] ),
    .A1(\cpuregs[29][15] ),
    .S(net646),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_1 _10898_ (.A0(\cpuregs[30][15] ),
    .A1(\cpuregs[31][15] ),
    .S(net649),
    .X(_05583_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(_05582_),
    .A1(_05583_),
    .S(net796),
    .X(_05584_));
 sky130_fd_sc_hd__or2_1 _10900_ (.A(\cpuregs[24][15] ),
    .B(net649),
    .X(_05585_));
 sky130_fd_sc_hd__o211a_1 _10901_ (.A1(\cpuregs[25][15] ),
    .A2(net617),
    .B1(net603),
    .C1(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__or2_1 _10902_ (.A(\cpuregs[26][15] ),
    .B(net646),
    .X(_05587_));
 sky130_fd_sc_hd__o211a_1 _10903_ (.A1(\cpuregs[27][15] ),
    .A2(net617),
    .B1(net589),
    .C1(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a2111o_1 _10904_ (.A1(net822),
    .A2(_05584_),
    .B1(_05586_),
    .C1(_05588_),
    .D1(net787),
    .X(_05589_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\cpuregs[22][15] ),
    .A1(\cpuregs[23][15] ),
    .S(net646),
    .X(_05590_));
 sky130_fd_sc_hd__mux2_1 _10906_ (.A0(\cpuregs[20][15] ),
    .A1(\cpuregs[21][15] ),
    .S(net646),
    .X(_05591_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(_05590_),
    .A1(_05591_),
    .S(net809),
    .X(_05592_));
 sky130_fd_sc_hd__or2_1 _10908_ (.A(\cpuregs[16][15] ),
    .B(net646),
    .X(_05593_));
 sky130_fd_sc_hd__o211a_1 _10909_ (.A1(\cpuregs[17][15] ),
    .A2(net617),
    .B1(net603),
    .C1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__o21a_1 _10910_ (.A1(\cpuregs[19][15] ),
    .A2(net617),
    .B1(net589),
    .X(_05595_));
 sky130_fd_sc_hd__o22a_1 _10911_ (.A1(\cpuregs[18][15] ),
    .A2(net552),
    .B1(_05595_),
    .B2(net779),
    .X(_05596_));
 sky130_fd_sc_hd__a211o_1 _10912_ (.A1(net822),
    .A2(_05592_),
    .B1(_05594_),
    .C1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__and3_1 _10913_ (.A(net772),
    .B(_05589_),
    .C(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__a21oi_4 _10914_ (.A1(_05572_),
    .A2(_05581_),
    .B1(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__or2_1 _10915_ (.A(net1075),
    .B(\decoded_imm[15] ),
    .X(_05600_));
 sky130_fd_sc_hd__a21oi_1 _10916_ (.A1(net1076),
    .A2(_05599_),
    .B1(net853),
    .Y(_05601_));
 sky130_fd_sc_hd__a22o_1 _10917_ (.A1(net1162),
    .A2(net853),
    .B1(_05600_),
    .B2(_05601_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(\cpuregs[6][16] ),
    .A1(\cpuregs[7][16] ),
    .S(net659),
    .X(_05602_));
 sky130_fd_sc_hd__mux2_1 _10919_ (.A0(\cpuregs[4][16] ),
    .A1(\cpuregs[5][16] ),
    .S(net659),
    .X(_05603_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(_05602_),
    .A1(_05603_),
    .S(net811),
    .X(_05604_));
 sky130_fd_sc_hd__or2_1 _10921_ (.A(\cpuregs[0][16] ),
    .B(net658),
    .X(_05605_));
 sky130_fd_sc_hd__o211a_1 _10922_ (.A1(\cpuregs[1][16] ),
    .A2(net622),
    .B1(net605),
    .C1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__or2_1 _10923_ (.A(\cpuregs[2][16] ),
    .B(net659),
    .X(_05607_));
 sky130_fd_sc_hd__o211a_1 _10924_ (.A1(\cpuregs[3][16] ),
    .A2(net623),
    .B1(net591),
    .C1(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__a211o_1 _10925_ (.A1(net825),
    .A2(_05604_),
    .B1(_05608_),
    .C1(net782),
    .X(_05609_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\cpuregs[14][16] ),
    .A1(\cpuregs[15][16] ),
    .S(net657),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(\cpuregs[12][16] ),
    .A1(\cpuregs[13][16] ),
    .S(net655),
    .X(_05611_));
 sky130_fd_sc_hd__or2_1 _10928_ (.A(net798),
    .B(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__o211a_1 _10929_ (.A1(net810),
    .A2(_05610_),
    .B1(_05612_),
    .C1(net824),
    .X(_05613_));
 sky130_fd_sc_hd__or2_1 _10930_ (.A(\cpuregs[8][16] ),
    .B(net657),
    .X(_05614_));
 sky130_fd_sc_hd__o211a_1 _10931_ (.A1(\cpuregs[9][16] ),
    .A2(net621),
    .B1(net605),
    .C1(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__or2_1 _10932_ (.A(\cpuregs[10][16] ),
    .B(net655),
    .X(_05616_));
 sky130_fd_sc_hd__o211a_1 _10933_ (.A1(\cpuregs[11][16] ),
    .A2(net621),
    .B1(net591),
    .C1(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__or4_1 _10934_ (.A(net788),
    .B(_05613_),
    .C(_05615_),
    .D(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__o21a_1 _10935_ (.A1(_05606_),
    .A2(_05609_),
    .B1(_03171_),
    .X(_05619_));
 sky130_fd_sc_hd__mux2_1 _10936_ (.A0(\cpuregs[20][16] ),
    .A1(\cpuregs[21][16] ),
    .S(net655),
    .X(_05620_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(\cpuregs[22][16] ),
    .A1(\cpuregs[23][16] ),
    .S(net655),
    .X(_05621_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(_05620_),
    .A1(_05621_),
    .S(net798),
    .X(_05622_));
 sky130_fd_sc_hd__or2_1 _10939_ (.A(\cpuregs[16][16] ),
    .B(net655),
    .X(_05623_));
 sky130_fd_sc_hd__o211a_1 _10940_ (.A1(\cpuregs[17][16] ),
    .A2(net621),
    .B1(net605),
    .C1(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__o21a_1 _10941_ (.A1(\cpuregs[19][16] ),
    .A2(net621),
    .B1(net591),
    .X(_05625_));
 sky130_fd_sc_hd__o22a_1 _10942_ (.A1(\cpuregs[18][16] ),
    .A2(net552),
    .B1(_05625_),
    .B2(net779),
    .X(_05626_));
 sky130_fd_sc_hd__a211o_1 _10943_ (.A1(net824),
    .A2(_05622_),
    .B1(_05624_),
    .C1(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__mux2_1 _10944_ (.A0(\cpuregs[30][16] ),
    .A1(\cpuregs[31][16] ),
    .S(net656),
    .X(_05628_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(\cpuregs[28][16] ),
    .A1(\cpuregs[29][16] ),
    .S(net656),
    .X(_05629_));
 sky130_fd_sc_hd__mux2_1 _10946_ (.A0(_05628_),
    .A1(_05629_),
    .S(net810),
    .X(_05630_));
 sky130_fd_sc_hd__or2_1 _10947_ (.A(\cpuregs[24][16] ),
    .B(net656),
    .X(_05631_));
 sky130_fd_sc_hd__o211a_1 _10948_ (.A1(\cpuregs[25][16] ),
    .A2(net621),
    .B1(net605),
    .C1(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__or2_1 _10949_ (.A(\cpuregs[26][16] ),
    .B(net656),
    .X(_05633_));
 sky130_fd_sc_hd__o211a_1 _10950_ (.A1(\cpuregs[27][16] ),
    .A2(net621),
    .B1(net591),
    .C1(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__a2111o_1 _10951_ (.A1(net824),
    .A2(_05630_),
    .B1(_05632_),
    .C1(_05634_),
    .D1(net788),
    .X(_05635_));
 sky130_fd_sc_hd__and3_1 _10952_ (.A(net772),
    .B(_05627_),
    .C(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__a21oi_4 _10953_ (.A1(_05618_),
    .A2(_05619_),
    .B1(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__or2_1 _10954_ (.A(net1075),
    .B(\decoded_imm[16] ),
    .X(_05638_));
 sky130_fd_sc_hd__a21oi_1 _10955_ (.A1(net1078),
    .A2(_05637_),
    .B1(net855),
    .Y(_05639_));
 sky130_fd_sc_hd__a22o_1 _10956_ (.A1(net1161),
    .A2(net855),
    .B1(_05638_),
    .B2(_05639_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(\cpuregs[6][17] ),
    .A1(\cpuregs[7][17] ),
    .S(net659),
    .X(_05640_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(\cpuregs[4][17] ),
    .A1(\cpuregs[5][17] ),
    .S(net659),
    .X(_05641_));
 sky130_fd_sc_hd__mux2_1 _10959_ (.A0(_05640_),
    .A1(_05641_),
    .S(net811),
    .X(_05642_));
 sky130_fd_sc_hd__or2_1 _10960_ (.A(\cpuregs[0][17] ),
    .B(net656),
    .X(_05643_));
 sky130_fd_sc_hd__o211a_1 _10961_ (.A1(\cpuregs[1][17] ),
    .A2(net621),
    .B1(net605),
    .C1(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__or2_1 _10962_ (.A(\cpuregs[2][17] ),
    .B(net659),
    .X(_05645_));
 sky130_fd_sc_hd__o211a_1 _10963_ (.A1(\cpuregs[3][17] ),
    .A2(net623),
    .B1(net592),
    .C1(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__a211o_1 _10964_ (.A1(net825),
    .A2(_05642_),
    .B1(_05646_),
    .C1(net779),
    .X(_05647_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(\cpuregs[12][17] ),
    .A1(\cpuregs[13][17] ),
    .S(net655),
    .X(_05648_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(\cpuregs[14][17] ),
    .A1(\cpuregs[15][17] ),
    .S(net655),
    .X(_05649_));
 sky130_fd_sc_hd__or2_1 _10967_ (.A(net810),
    .B(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__o211a_1 _10968_ (.A1(net798),
    .A2(_05648_),
    .B1(_05650_),
    .C1(net824),
    .X(_05651_));
 sky130_fd_sc_hd__or2_1 _10969_ (.A(\cpuregs[8][17] ),
    .B(net655),
    .X(_05652_));
 sky130_fd_sc_hd__o211a_1 _10970_ (.A1(\cpuregs[9][17] ),
    .A2(net621),
    .B1(net605),
    .C1(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__or2_1 _10971_ (.A(\cpuregs[10][17] ),
    .B(net655),
    .X(_05654_));
 sky130_fd_sc_hd__o211a_1 _10972_ (.A1(\cpuregs[11][17] ),
    .A2(net621),
    .B1(net590),
    .C1(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__or4_1 _10973_ (.A(net791),
    .B(_05651_),
    .C(_05653_),
    .D(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__o21a_1 _10974_ (.A1(_05644_),
    .A2(_05647_),
    .B1(_03171_),
    .X(_05657_));
 sky130_fd_sc_hd__mux2_1 _10975_ (.A0(\cpuregs[22][17] ),
    .A1(\cpuregs[23][17] ),
    .S(net646),
    .X(_05658_));
 sky130_fd_sc_hd__mux2_1 _10976_ (.A0(\cpuregs[20][17] ),
    .A1(\cpuregs[21][17] ),
    .S(net646),
    .X(_05659_));
 sky130_fd_sc_hd__mux2_1 _10977_ (.A0(_05658_),
    .A1(_05659_),
    .S(net809),
    .X(_05660_));
 sky130_fd_sc_hd__or2_1 _10978_ (.A(\cpuregs[16][17] ),
    .B(net647),
    .X(_05661_));
 sky130_fd_sc_hd__o211a_1 _10979_ (.A1(\cpuregs[17][17] ),
    .A2(net617),
    .B1(net603),
    .C1(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__o21a_1 _10980_ (.A1(\cpuregs[19][17] ),
    .A2(net617),
    .B1(net589),
    .X(_05663_));
 sky130_fd_sc_hd__o22a_1 _10981_ (.A1(\cpuregs[18][17] ),
    .A2(net552),
    .B1(_05663_),
    .B2(net779),
    .X(_05664_));
 sky130_fd_sc_hd__a211o_1 _10982_ (.A1(net822),
    .A2(_05660_),
    .B1(_05662_),
    .C1(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__mux2_1 _10983_ (.A0(\cpuregs[28][17] ),
    .A1(\cpuregs[29][17] ),
    .S(net646),
    .X(_05666_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\cpuregs[30][17] ),
    .A1(\cpuregs[31][17] ),
    .S(net647),
    .X(_05667_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(_05666_),
    .A1(_05667_),
    .S(net796),
    .X(_05668_));
 sky130_fd_sc_hd__or2_1 _10986_ (.A(\cpuregs[24][17] ),
    .B(net648),
    .X(_05669_));
 sky130_fd_sc_hd__o211a_1 _10987_ (.A1(\cpuregs[25][17] ),
    .A2(net617),
    .B1(net603),
    .C1(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__or2_1 _10988_ (.A(\cpuregs[26][17] ),
    .B(net649),
    .X(_05671_));
 sky130_fd_sc_hd__o211a_1 _10989_ (.A1(\cpuregs[27][17] ),
    .A2(net617),
    .B1(net589),
    .C1(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__a2111o_1 _10990_ (.A1(net822),
    .A2(_05668_),
    .B1(_05670_),
    .C1(_05672_),
    .D1(net787),
    .X(_05673_));
 sky130_fd_sc_hd__and3_1 _10991_ (.A(net772),
    .B(_05665_),
    .C(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__a21oi_4 _10992_ (.A1(_05656_),
    .A2(_05657_),
    .B1(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(net1078),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__o21a_1 _10994_ (.A1(net1078),
    .A2(\decoded_imm[17] ),
    .B1(net860),
    .X(_05677_));
 sky130_fd_sc_hd__a22o_1 _10995_ (.A1(net1160),
    .A2(net855),
    .B1(_05676_),
    .B2(_05677_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(\cpuregs[6][18] ),
    .A1(\cpuregs[7][18] ),
    .S(net652),
    .X(_05678_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(\cpuregs[4][18] ),
    .A1(\cpuregs[5][18] ),
    .S(net652),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(_05678_),
    .A1(_05679_),
    .S(net809),
    .X(_05680_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(\cpuregs[2][18] ),
    .A1(\cpuregs[3][18] ),
    .S(net648),
    .X(_05681_));
 sky130_fd_sc_hd__a221o_1 _11000_ (.A1(\cpuregs[1][18] ),
    .A2(net549),
    .B1(_05681_),
    .B2(net796),
    .C1(net823),
    .X(_05682_));
 sky130_fd_sc_hd__o21a_1 _11001_ (.A1(net838),
    .A2(_05680_),
    .B1(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(\cpuregs[12][18] ),
    .A1(\cpuregs[13][18] ),
    .S(net647),
    .X(_05684_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\cpuregs[14][18] ),
    .A1(\cpuregs[15][18] ),
    .S(net655),
    .X(_05685_));
 sky130_fd_sc_hd__or2_1 _11004_ (.A(net809),
    .B(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__o211a_1 _11005_ (.A1(net796),
    .A2(_05684_),
    .B1(_05686_),
    .C1(net823),
    .X(_05687_));
 sky130_fd_sc_hd__or2_1 _11006_ (.A(\cpuregs[8][18] ),
    .B(net648),
    .X(_05688_));
 sky130_fd_sc_hd__o211a_1 _11007_ (.A1(\cpuregs[9][18] ),
    .A2(net618),
    .B1(net603),
    .C1(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__or2_1 _11008_ (.A(\cpuregs[10][18] ),
    .B(net647),
    .X(_05690_));
 sky130_fd_sc_hd__o211a_1 _11009_ (.A1(\cpuregs[11][18] ),
    .A2(net618),
    .B1(net589),
    .C1(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__or4_1 _11010_ (.A(net787),
    .B(_05687_),
    .C(_05689_),
    .D(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__o211a_1 _11011_ (.A1(net779),
    .A2(_05683_),
    .B1(_05692_),
    .C1(net776),
    .X(_05693_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(\cpuregs[30][18] ),
    .A1(\cpuregs[31][18] ),
    .S(net648),
    .X(_05694_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(\cpuregs[28][18] ),
    .A1(\cpuregs[29][18] ),
    .S(net648),
    .X(_05695_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(_05694_),
    .A1(_05695_),
    .S(net809),
    .X(_05696_));
 sky130_fd_sc_hd__or2_1 _11015_ (.A(\cpuregs[24][18] ),
    .B(net648),
    .X(_05697_));
 sky130_fd_sc_hd__o211a_1 _11016_ (.A1(\cpuregs[25][18] ),
    .A2(net618),
    .B1(net603),
    .C1(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__or2_1 _11017_ (.A(\cpuregs[26][18] ),
    .B(net648),
    .X(_05699_));
 sky130_fd_sc_hd__o211a_1 _11018_ (.A1(\cpuregs[27][18] ),
    .A2(net618),
    .B1(net589),
    .C1(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__a2111o_1 _11019_ (.A1(net822),
    .A2(_05696_),
    .B1(_05698_),
    .C1(_05700_),
    .D1(net787),
    .X(_05701_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(\cpuregs[22][18] ),
    .A1(\cpuregs[23][18] ),
    .S(net647),
    .X(_05702_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(\cpuregs[20][18] ),
    .A1(\cpuregs[21][18] ),
    .S(net647),
    .X(_05703_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(_05702_),
    .A1(_05703_),
    .S(net809),
    .X(_05704_));
 sky130_fd_sc_hd__or2_1 _11023_ (.A(\cpuregs[16][18] ),
    .B(net647),
    .X(_05705_));
 sky130_fd_sc_hd__o211a_1 _11024_ (.A1(\cpuregs[17][18] ),
    .A2(net618),
    .B1(net603),
    .C1(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__o21a_1 _11025_ (.A1(\cpuregs[19][18] ),
    .A2(net618),
    .B1(net589),
    .X(_05707_));
 sky130_fd_sc_hd__o22a_1 _11026_ (.A1(\cpuregs[18][18] ),
    .A2(net552),
    .B1(_05707_),
    .B2(net779),
    .X(_05708_));
 sky130_fd_sc_hd__a211o_1 _11027_ (.A1(net822),
    .A2(_05704_),
    .B1(_05706_),
    .C1(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__a31oi_4 _11028_ (.A1(net772),
    .A2(_05701_),
    .A3(_05709_),
    .B1(_05693_),
    .Y(_05710_));
 sky130_fd_sc_hd__or2_1 _11029_ (.A(net1075),
    .B(\decoded_imm[18] ),
    .X(_05711_));
 sky130_fd_sc_hd__a21oi_1 _11030_ (.A1(net1075),
    .A2(_05710_),
    .B1(net855),
    .Y(_05712_));
 sky130_fd_sc_hd__a22o_1 _11031_ (.A1(net244),
    .A2(net855),
    .B1(_05711_),
    .B2(_05712_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(\cpuregs[6][19] ),
    .A1(\cpuregs[7][19] ),
    .S(net684),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(\cpuregs[4][19] ),
    .A1(\cpuregs[5][19] ),
    .S(net684),
    .X(_05714_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(_05713_),
    .A1(_05714_),
    .S(net816),
    .X(_05715_));
 sky130_fd_sc_hd__or2_1 _11035_ (.A(\cpuregs[0][19] ),
    .B(net681),
    .X(_05716_));
 sky130_fd_sc_hd__o211a_1 _11036_ (.A1(\cpuregs[1][19] ),
    .A2(net632),
    .B1(net610),
    .C1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__or2_1 _11037_ (.A(\cpuregs[2][19] ),
    .B(net681),
    .X(_05718_));
 sky130_fd_sc_hd__o211a_1 _11038_ (.A1(\cpuregs[3][19] ),
    .A2(net632),
    .B1(net597),
    .C1(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__a211o_1 _11039_ (.A1(net831),
    .A2(_05715_),
    .B1(_05719_),
    .C1(net784),
    .X(_05720_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(\cpuregs[12][19] ),
    .A1(\cpuregs[13][19] ),
    .S(net680),
    .X(_05721_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(\cpuregs[14][19] ),
    .A1(\cpuregs[15][19] ),
    .S(net680),
    .X(_05722_));
 sky130_fd_sc_hd__or2_1 _11042_ (.A(net816),
    .B(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__o211a_1 _11043_ (.A1(net804),
    .A2(_05721_),
    .B1(_05723_),
    .C1(net831),
    .X(_05724_));
 sky130_fd_sc_hd__or2_1 _11044_ (.A(\cpuregs[8][19] ),
    .B(net680),
    .X(_05725_));
 sky130_fd_sc_hd__o211a_1 _11045_ (.A1(\cpuregs[9][19] ),
    .A2(net632),
    .B1(net610),
    .C1(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__or2_1 _11046_ (.A(\cpuregs[10][19] ),
    .B(net680),
    .X(_05727_));
 sky130_fd_sc_hd__o211a_1 _11047_ (.A1(\cpuregs[11][19] ),
    .A2(net632),
    .B1(net597),
    .C1(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__or4_1 _11048_ (.A(net792),
    .B(_05724_),
    .C(_05726_),
    .D(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__o21a_1 _11049_ (.A1(_05717_),
    .A2(_05720_),
    .B1(_03171_),
    .X(_05730_));
 sky130_fd_sc_hd__mux2_1 _11050_ (.A0(\cpuregs[22][19] ),
    .A1(\cpuregs[23][19] ),
    .S(net680),
    .X(_05731_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(\cpuregs[20][19] ),
    .A1(\cpuregs[21][19] ),
    .S(net680),
    .X(_05732_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(_05731_),
    .A1(_05732_),
    .S(net816),
    .X(_05733_));
 sky130_fd_sc_hd__or2_1 _11053_ (.A(\cpuregs[16][19] ),
    .B(net680),
    .X(_05734_));
 sky130_fd_sc_hd__o211a_1 _11054_ (.A1(\cpuregs[17][19] ),
    .A2(net632),
    .B1(net610),
    .C1(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__o21a_1 _11055_ (.A1(\cpuregs[19][19] ),
    .A2(net632),
    .B1(net597),
    .X(_05736_));
 sky130_fd_sc_hd__o22a_1 _11056_ (.A1(\cpuregs[18][19] ),
    .A2(net554),
    .B1(_05736_),
    .B2(net784),
    .X(_05737_));
 sky130_fd_sc_hd__a211o_1 _11057_ (.A1(net831),
    .A2(_05733_),
    .B1(_05735_),
    .C1(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(\cpuregs[30][19] ),
    .A1(\cpuregs[31][19] ),
    .S(net681),
    .X(_05739_));
 sky130_fd_sc_hd__mux2_1 _11059_ (.A0(\cpuregs[28][19] ),
    .A1(\cpuregs[29][19] ),
    .S(net681),
    .X(_05740_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(_05739_),
    .A1(_05740_),
    .S(net816),
    .X(_05741_));
 sky130_fd_sc_hd__or2_1 _11061_ (.A(\cpuregs[24][19] ),
    .B(net681),
    .X(_05742_));
 sky130_fd_sc_hd__o211a_1 _11062_ (.A1(\cpuregs[25][19] ),
    .A2(net632),
    .B1(net610),
    .C1(_05742_),
    .X(_05743_));
 sky130_fd_sc_hd__or2_1 _11063_ (.A(\cpuregs[26][19] ),
    .B(net680),
    .X(_05744_));
 sky130_fd_sc_hd__o211a_1 _11064_ (.A1(\cpuregs[27][19] ),
    .A2(net632),
    .B1(net597),
    .C1(_05744_),
    .X(_05745_));
 sky130_fd_sc_hd__a2111o_1 _11065_ (.A1(net831),
    .A2(_05741_),
    .B1(_05743_),
    .C1(_05745_),
    .D1(net792),
    .X(_05746_));
 sky130_fd_sc_hd__and3_1 _11066_ (.A(net774),
    .B(_05738_),
    .C(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__a21oi_4 _11067_ (.A1(_05729_),
    .A2(_05730_),
    .B1(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__or2_1 _11068_ (.A(net1075),
    .B(\decoded_imm[19] ),
    .X(_05749_));
 sky130_fd_sc_hd__a21oi_1 _11069_ (.A1(\cpu_state[3] ),
    .A2(_05748_),
    .B1(net856),
    .Y(_05750_));
 sky130_fd_sc_hd__a22o_1 _11070_ (.A1(net1159),
    .A2(net856),
    .B1(_05749_),
    .B2(_05750_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _11071_ (.A0(\cpuregs[30][20] ),
    .A1(\cpuregs[31][20] ),
    .S(net661),
    .X(_05751_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(\cpuregs[28][20] ),
    .A1(\cpuregs[29][20] ),
    .S(net661),
    .X(_05752_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(_05751_),
    .A1(_05752_),
    .S(net810),
    .X(_05753_));
 sky130_fd_sc_hd__or2_1 _11074_ (.A(\cpuregs[24][20] ),
    .B(net658),
    .X(_05754_));
 sky130_fd_sc_hd__o211a_1 _11075_ (.A1(\cpuregs[25][20] ),
    .A2(net622),
    .B1(net605),
    .C1(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__or2_1 _11076_ (.A(\cpuregs[26][20] ),
    .B(net658),
    .X(_05756_));
 sky130_fd_sc_hd__o211a_1 _11077_ (.A1(\cpuregs[27][20] ),
    .A2(net622),
    .B1(net591),
    .C1(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__a2111o_1 _11078_ (.A1(net824),
    .A2(_05753_),
    .B1(_05755_),
    .C1(_05757_),
    .D1(net788),
    .X(_05758_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(\cpuregs[20][20] ),
    .A1(\cpuregs[21][20] ),
    .S(net657),
    .X(_05759_));
 sky130_fd_sc_hd__mux2_1 _11080_ (.A0(\cpuregs[22][20] ),
    .A1(\cpuregs[23][20] ),
    .S(net657),
    .X(_05760_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(_05759_),
    .A1(_05760_),
    .S(net798),
    .X(_05761_));
 sky130_fd_sc_hd__or2_1 _11082_ (.A(\cpuregs[16][20] ),
    .B(net657),
    .X(_05762_));
 sky130_fd_sc_hd__o211a_1 _11083_ (.A1(\cpuregs[17][20] ),
    .A2(net624),
    .B1(net605),
    .C1(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__o21a_1 _11084_ (.A1(\cpuregs[19][20] ),
    .A2(net622),
    .B1(net591),
    .X(_05764_));
 sky130_fd_sc_hd__o22a_1 _11085_ (.A1(\cpuregs[18][20] ),
    .A2(net552),
    .B1(_05764_),
    .B2(net782),
    .X(_05765_));
 sky130_fd_sc_hd__a211o_1 _11086_ (.A1(net824),
    .A2(_05761_),
    .B1(_05763_),
    .C1(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__and3_1 _11087_ (.A(net772),
    .B(_05758_),
    .C(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(\cpuregs[6][20] ),
    .A1(\cpuregs[7][20] ),
    .S(net661),
    .X(_05768_));
 sky130_fd_sc_hd__or2_1 _11089_ (.A(\cpuregs[4][20] ),
    .B(net661),
    .X(_05769_));
 sky130_fd_sc_hd__o211a_1 _11090_ (.A1(\cpuregs[5][20] ),
    .A2(net624),
    .B1(net811),
    .C1(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__a211o_1 _11091_ (.A1(net798),
    .A2(_05768_),
    .B1(_05770_),
    .C1(net838),
    .X(_05771_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(\cpuregs[2][20] ),
    .A1(\cpuregs[3][20] ),
    .S(net661),
    .X(_05772_));
 sky130_fd_sc_hd__a221o_1 _11093_ (.A1(\cpuregs[1][20] ),
    .A2(net549),
    .B1(_05772_),
    .B2(net799),
    .C1(net825),
    .X(_05773_));
 sky130_fd_sc_hd__a21o_1 _11094_ (.A1(_05771_),
    .A2(_05773_),
    .B1(net782),
    .X(_05774_));
 sky130_fd_sc_hd__mux2_1 _11095_ (.A0(\cpuregs[12][20] ),
    .A1(\cpuregs[13][20] ),
    .S(net657),
    .X(_05775_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(\cpuregs[14][20] ),
    .A1(\cpuregs[15][20] ),
    .S(net657),
    .X(_05776_));
 sky130_fd_sc_hd__or2_1 _11097_ (.A(net810),
    .B(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__o211a_1 _11098_ (.A1(net798),
    .A2(_05775_),
    .B1(_05777_),
    .C1(net824),
    .X(_05778_));
 sky130_fd_sc_hd__or2_1 _11099_ (.A(\cpuregs[8][20] ),
    .B(net657),
    .X(_05779_));
 sky130_fd_sc_hd__o211a_1 _11100_ (.A1(\cpuregs[9][20] ),
    .A2(net622),
    .B1(net605),
    .C1(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__or2_1 _11101_ (.A(\cpuregs[10][20] ),
    .B(net657),
    .X(_05781_));
 sky130_fd_sc_hd__o211a_1 _11102_ (.A1(\cpuregs[11][20] ),
    .A2(net622),
    .B1(net591),
    .C1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__o41a_1 _11103_ (.A1(net788),
    .A2(_05778_),
    .A3(_05780_),
    .A4(_05782_),
    .B1(net776),
    .X(_05783_));
 sky130_fd_sc_hd__a21oi_4 _11104_ (.A1(_05774_),
    .A2(_05783_),
    .B1(_05767_),
    .Y(_05784_));
 sky130_fd_sc_hd__or2_1 _11105_ (.A(net1081),
    .B(\decoded_imm[20] ),
    .X(_05785_));
 sky130_fd_sc_hd__a21oi_1 _11106_ (.A1(net1082),
    .A2(_05784_),
    .B1(net859),
    .Y(_05786_));
 sky130_fd_sc_hd__a22o_1 _11107_ (.A1(net247),
    .A2(net856),
    .B1(_05785_),
    .B2(_05786_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(\cpuregs[6][21] ),
    .A1(\cpuregs[7][21] ),
    .S(net685),
    .X(_05787_));
 sky130_fd_sc_hd__or2_1 _11109_ (.A(\cpuregs[4][21] ),
    .B(net684),
    .X(_05788_));
 sky130_fd_sc_hd__o211a_1 _11110_ (.A1(\cpuregs[5][21] ),
    .A2(net634),
    .B1(net818),
    .C1(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__a211o_1 _11111_ (.A1(net804),
    .A2(_05787_),
    .B1(_05789_),
    .C1(net840),
    .X(_05790_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(\cpuregs[2][21] ),
    .A1(\cpuregs[3][21] ),
    .S(net685),
    .X(_05791_));
 sky130_fd_sc_hd__a221o_1 _11113_ (.A1(\cpuregs[1][21] ),
    .A2(net549),
    .B1(_05791_),
    .B2(net804),
    .C1(net825),
    .X(_05792_));
 sky130_fd_sc_hd__a21o_1 _11114_ (.A1(_05790_),
    .A2(_05792_),
    .B1(net784),
    .X(_05793_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(\cpuregs[14][21] ),
    .A1(\cpuregs[15][21] ),
    .S(net661),
    .X(_05794_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(\cpuregs[12][21] ),
    .A1(\cpuregs[13][21] ),
    .S(net661),
    .X(_05795_));
 sky130_fd_sc_hd__or2_1 _11117_ (.A(net799),
    .B(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__o211a_1 _11118_ (.A1(net810),
    .A2(_05794_),
    .B1(_05796_),
    .C1(net825),
    .X(_05797_));
 sky130_fd_sc_hd__or2_1 _11119_ (.A(\cpuregs[8][21] ),
    .B(net661),
    .X(_05798_));
 sky130_fd_sc_hd__o211a_1 _11120_ (.A1(\cpuregs[9][21] ),
    .A2(net623),
    .B1(net606),
    .C1(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__or2_1 _11121_ (.A(\cpuregs[10][21] ),
    .B(net684),
    .X(_05800_));
 sky130_fd_sc_hd__o211a_1 _11122_ (.A1(\cpuregs[11][21] ),
    .A2(net634),
    .B1(net591),
    .C1(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__o41a_1 _11123_ (.A1(net791),
    .A2(_05797_),
    .A3(_05799_),
    .A4(_05801_),
    .B1(net776),
    .X(_05802_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(\cpuregs[30][21] ),
    .A1(\cpuregs[31][21] ),
    .S(net658),
    .X(_05803_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(\cpuregs[28][21] ),
    .A1(\cpuregs[29][21] ),
    .S(net658),
    .X(_05804_));
 sky130_fd_sc_hd__mux2_1 _11126_ (.A0(_05803_),
    .A1(_05804_),
    .S(net810),
    .X(_05805_));
 sky130_fd_sc_hd__or2_1 _11127_ (.A(\cpuregs[24][21] ),
    .B(net658),
    .X(_05806_));
 sky130_fd_sc_hd__o211a_1 _11128_ (.A1(\cpuregs[25][21] ),
    .A2(net622),
    .B1(net605),
    .C1(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__or2_1 _11129_ (.A(\cpuregs[26][21] ),
    .B(net681),
    .X(_05808_));
 sky130_fd_sc_hd__o211a_1 _11130_ (.A1(\cpuregs[27][21] ),
    .A2(net632),
    .B1(net591),
    .C1(_05808_),
    .X(_05809_));
 sky130_fd_sc_hd__a2111o_1 _11131_ (.A1(net824),
    .A2(_05805_),
    .B1(_05807_),
    .C1(_05809_),
    .D1(net788),
    .X(_05810_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(\cpuregs[20][21] ),
    .A1(\cpuregs[21][21] ),
    .S(net657),
    .X(_05811_));
 sky130_fd_sc_hd__mux2_1 _11133_ (.A0(\cpuregs[22][21] ),
    .A1(\cpuregs[23][21] ),
    .S(net680),
    .X(_05812_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(_05811_),
    .A1(_05812_),
    .S(net798),
    .X(_05813_));
 sky130_fd_sc_hd__or2_1 _11135_ (.A(\cpuregs[16][21] ),
    .B(net680),
    .X(_05814_));
 sky130_fd_sc_hd__o211a_1 _11136_ (.A1(\cpuregs[17][21] ),
    .A2(net622),
    .B1(net610),
    .C1(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__o21a_1 _11137_ (.A1(\cpuregs[19][21] ),
    .A2(net622),
    .B1(net591),
    .X(_05816_));
 sky130_fd_sc_hd__o22a_1 _11138_ (.A1(\cpuregs[18][21] ),
    .A2(net554),
    .B1(_05816_),
    .B2(net784),
    .X(_05817_));
 sky130_fd_sc_hd__a211o_1 _11139_ (.A1(net824),
    .A2(_05813_),
    .B1(_05815_),
    .C1(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__and3_1 _11140_ (.A(net774),
    .B(_05810_),
    .C(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__a21oi_4 _11141_ (.A1(_05793_),
    .A2(_05802_),
    .B1(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__or2_1 _11142_ (.A(net1080),
    .B(\decoded_imm[21] ),
    .X(_05821_));
 sky130_fd_sc_hd__a21oi_1 _11143_ (.A1(net1082),
    .A2(_05820_),
    .B1(net856),
    .Y(_05822_));
 sky130_fd_sc_hd__a22o_1 _11144_ (.A1(net248),
    .A2(net859),
    .B1(_05821_),
    .B2(_05822_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _11145_ (.A0(\cpuregs[6][22] ),
    .A1(\cpuregs[7][22] ),
    .S(net686),
    .X(_05823_));
 sky130_fd_sc_hd__mux2_1 _11146_ (.A0(\cpuregs[4][22] ),
    .A1(\cpuregs[5][22] ),
    .S(net686),
    .X(_05824_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(_05823_),
    .A1(_05824_),
    .S(net816),
    .X(_05825_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(\cpuregs[2][22] ),
    .A1(\cpuregs[3][22] ),
    .S(net683),
    .X(_05826_));
 sky130_fd_sc_hd__a221o_1 _11149_ (.A1(\cpuregs[1][22] ),
    .A2(net551),
    .B1(_05826_),
    .B2(net804),
    .C1(net831),
    .X(_05827_));
 sky130_fd_sc_hd__o21a_1 _11150_ (.A1(net840),
    .A2(_05825_),
    .B1(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__mux2_1 _11151_ (.A0(\cpuregs[12][22] ),
    .A1(\cpuregs[13][22] ),
    .S(net682),
    .X(_05829_));
 sky130_fd_sc_hd__mux2_1 _11152_ (.A0(\cpuregs[14][22] ),
    .A1(\cpuregs[15][22] ),
    .S(net682),
    .X(_05830_));
 sky130_fd_sc_hd__or2_1 _11153_ (.A(net816),
    .B(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__o211a_1 _11154_ (.A1(net804),
    .A2(_05829_),
    .B1(_05831_),
    .C1(net831),
    .X(_05832_));
 sky130_fd_sc_hd__or2_1 _11155_ (.A(\cpuregs[8][22] ),
    .B(net682),
    .X(_05833_));
 sky130_fd_sc_hd__o211a_1 _11156_ (.A1(\cpuregs[9][22] ),
    .A2(net633),
    .B1(net610),
    .C1(_05833_),
    .X(_05834_));
 sky130_fd_sc_hd__or2_1 _11157_ (.A(\cpuregs[10][22] ),
    .B(net682),
    .X(_05835_));
 sky130_fd_sc_hd__o211a_1 _11158_ (.A1(\cpuregs[11][22] ),
    .A2(net633),
    .B1(net597),
    .C1(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__or4_1 _11159_ (.A(net792),
    .B(_05832_),
    .C(_05834_),
    .D(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__o211a_1 _11160_ (.A1(net783),
    .A2(_05828_),
    .B1(_05837_),
    .C1(net778),
    .X(_05838_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(\cpuregs[30][22] ),
    .A1(\cpuregs[31][22] ),
    .S(net683),
    .X(_05839_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(\cpuregs[28][22] ),
    .A1(\cpuregs[29][22] ),
    .S(net683),
    .X(_05840_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(_05839_),
    .A1(_05840_),
    .S(net816),
    .X(_05841_));
 sky130_fd_sc_hd__or2_1 _11164_ (.A(\cpuregs[24][22] ),
    .B(net683),
    .X(_05842_));
 sky130_fd_sc_hd__o211a_1 _11165_ (.A1(\cpuregs[25][22] ),
    .A2(net633),
    .B1(net610),
    .C1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__or2_1 _11166_ (.A(\cpuregs[26][22] ),
    .B(net683),
    .X(_05844_));
 sky130_fd_sc_hd__o211a_1 _11167_ (.A1(\cpuregs[27][22] ),
    .A2(net633),
    .B1(net597),
    .C1(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__a2111o_1 _11168_ (.A1(net831),
    .A2(_05841_),
    .B1(_05843_),
    .C1(_05845_),
    .D1(net792),
    .X(_05846_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(\cpuregs[20][22] ),
    .A1(\cpuregs[21][22] ),
    .S(net682),
    .X(_05847_));
 sky130_fd_sc_hd__mux2_1 _11170_ (.A0(\cpuregs[22][22] ),
    .A1(\cpuregs[23][22] ),
    .S(net682),
    .X(_05848_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(_05847_),
    .A1(_05848_),
    .S(net804),
    .X(_05849_));
 sky130_fd_sc_hd__or2_1 _11172_ (.A(\cpuregs[16][22] ),
    .B(net682),
    .X(_05850_));
 sky130_fd_sc_hd__o211a_1 _11173_ (.A1(\cpuregs[17][22] ),
    .A2(net633),
    .B1(net610),
    .C1(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__o21a_1 _11174_ (.A1(\cpuregs[19][22] ),
    .A2(net633),
    .B1(net597),
    .X(_05852_));
 sky130_fd_sc_hd__o22a_1 _11175_ (.A1(\cpuregs[18][22] ),
    .A2(net554),
    .B1(_05852_),
    .B2(net783),
    .X(_05853_));
 sky130_fd_sc_hd__a211o_1 _11176_ (.A1(net831),
    .A2(_05849_),
    .B1(_05851_),
    .C1(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__a31oi_4 _11177_ (.A1(net774),
    .A2(_05846_),
    .A3(_05854_),
    .B1(_05838_),
    .Y(_05855_));
 sky130_fd_sc_hd__or2_1 _11178_ (.A(net1081),
    .B(\decoded_imm[22] ),
    .X(_05856_));
 sky130_fd_sc_hd__a21oi_1 _11179_ (.A1(net1081),
    .A2(_05855_),
    .B1(net856),
    .Y(_05857_));
 sky130_fd_sc_hd__a22o_1 _11180_ (.A1(net1158),
    .A2(net856),
    .B1(_05856_),
    .B2(_05857_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _11181_ (.A0(\cpuregs[30][23] ),
    .A1(\cpuregs[31][23] ),
    .S(net697),
    .X(_05858_));
 sky130_fd_sc_hd__mux2_1 _11182_ (.A0(\cpuregs[28][23] ),
    .A1(\cpuregs[29][23] ),
    .S(net697),
    .X(_05859_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(_05858_),
    .A1(_05859_),
    .S(net819),
    .X(_05860_));
 sky130_fd_sc_hd__or2_1 _11184_ (.A(\cpuregs[24][23] ),
    .B(net685),
    .X(_05861_));
 sky130_fd_sc_hd__o211a_1 _11185_ (.A1(\cpuregs[25][23] ),
    .A2(net634),
    .B1(net610),
    .C1(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__or2_1 _11186_ (.A(\cpuregs[26][23] ),
    .B(net685),
    .X(_05863_));
 sky130_fd_sc_hd__o211a_1 _11187_ (.A1(\cpuregs[27][23] ),
    .A2(net634),
    .B1(net600),
    .C1(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__a2111o_1 _11188_ (.A1(net835),
    .A2(_05860_),
    .B1(_05862_),
    .C1(_05864_),
    .D1(net792),
    .X(_05865_));
 sky130_fd_sc_hd__mux2_1 _11189_ (.A0(\cpuregs[22][23] ),
    .A1(\cpuregs[23][23] ),
    .S(net675),
    .X(_05866_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(\cpuregs[20][23] ),
    .A1(\cpuregs[21][23] ),
    .S(net697),
    .X(_05867_));
 sky130_fd_sc_hd__mux2_1 _11191_ (.A0(_05866_),
    .A1(_05867_),
    .S(net815),
    .X(_05868_));
 sky130_fd_sc_hd__or2_1 _11192_ (.A(\cpuregs[16][23] ),
    .B(net685),
    .X(_05869_));
 sky130_fd_sc_hd__o211a_1 _11193_ (.A1(\cpuregs[17][23] ),
    .A2(net624),
    .B1(net611),
    .C1(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__o21a_1 _11194_ (.A1(\cpuregs[19][23] ),
    .A2(net630),
    .B1(net595),
    .X(_05871_));
 sky130_fd_sc_hd__o22a_1 _11195_ (.A1(\cpuregs[18][23] ),
    .A2(net554),
    .B1(_05871_),
    .B2(net785),
    .X(_05872_));
 sky130_fd_sc_hd__a211o_1 _11196_ (.A1(net835),
    .A2(_05868_),
    .B1(_05870_),
    .C1(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__mux2_1 _11197_ (.A0(\cpuregs[6][23] ),
    .A1(\cpuregs[7][23] ),
    .S(net675),
    .X(_05874_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(\cpuregs[4][23] ),
    .A1(\cpuregs[5][23] ),
    .S(net675),
    .X(_05875_));
 sky130_fd_sc_hd__mux2_1 _11199_ (.A0(_05874_),
    .A1(_05875_),
    .S(net821),
    .X(_05876_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(\cpuregs[2][23] ),
    .A1(\cpuregs[3][23] ),
    .S(net675),
    .X(_05877_));
 sky130_fd_sc_hd__a221o_1 _11201_ (.A1(\cpuregs[1][23] ),
    .A2(net550),
    .B1(_05877_),
    .B2(net801),
    .C1(net829),
    .X(_05878_));
 sky130_fd_sc_hd__o21a_1 _11202_ (.A1(net838),
    .A2(_05876_),
    .B1(_05878_),
    .X(_05879_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(\cpuregs[12][23] ),
    .A1(\cpuregs[13][23] ),
    .S(net662),
    .X(_05880_));
 sky130_fd_sc_hd__mux2_1 _11204_ (.A0(\cpuregs[14][23] ),
    .A1(\cpuregs[15][23] ),
    .S(net661),
    .X(_05881_));
 sky130_fd_sc_hd__or2_1 _11205_ (.A(net810),
    .B(_05881_),
    .X(_05882_));
 sky130_fd_sc_hd__o211a_1 _11206_ (.A1(net798),
    .A2(_05880_),
    .B1(_05882_),
    .C1(net825),
    .X(_05883_));
 sky130_fd_sc_hd__or2_1 _11207_ (.A(\cpuregs[8][23] ),
    .B(net662),
    .X(_05884_));
 sky130_fd_sc_hd__o211a_1 _11208_ (.A1(\cpuregs[9][23] ),
    .A2(net623),
    .B1(net606),
    .C1(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__or2_1 _11209_ (.A(\cpuregs[10][23] ),
    .B(net662),
    .X(_05886_));
 sky130_fd_sc_hd__o211a_1 _11210_ (.A1(\cpuregs[11][23] ),
    .A2(net623),
    .B1(net592),
    .C1(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__or4_1 _11211_ (.A(net788),
    .B(_05883_),
    .C(_05885_),
    .D(_05887_),
    .X(_05888_));
 sky130_fd_sc_hd__o211a_1 _11212_ (.A1(net785),
    .A2(_05879_),
    .B1(_05888_),
    .C1(net776),
    .X(_05889_));
 sky130_fd_sc_hd__a31oi_4 _11213_ (.A1(net774),
    .A2(_05865_),
    .A3(_05873_),
    .B1(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__nand2_1 _11214_ (.A(net1082),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__o21a_1 _11215_ (.A1(net1082),
    .A2(\decoded_imm[23] ),
    .B1(_05133_),
    .X(_05892_));
 sky130_fd_sc_hd__a22o_1 _11216_ (.A1(net250),
    .A2(net859),
    .B1(_05891_),
    .B2(_05892_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(\cpuregs[30][24] ),
    .A1(\cpuregs[31][24] ),
    .S(net697),
    .X(_05893_));
 sky130_fd_sc_hd__mux2_1 _11218_ (.A0(\cpuregs[28][24] ),
    .A1(\cpuregs[29][24] ),
    .S(net697),
    .X(_05894_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(_05893_),
    .A1(_05894_),
    .S(net819),
    .X(_05895_));
 sky130_fd_sc_hd__or2_1 _11220_ (.A(\cpuregs[24][24] ),
    .B(net699),
    .X(_05896_));
 sky130_fd_sc_hd__o211a_1 _11221_ (.A1(\cpuregs[25][24] ),
    .A2(net640),
    .B1(net614),
    .C1(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__or2_1 _11222_ (.A(\cpuregs[26][24] ),
    .B(net699),
    .X(_05898_));
 sky130_fd_sc_hd__o211a_1 _11223_ (.A1(\cpuregs[27][24] ),
    .A2(net640),
    .B1(net601),
    .C1(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__a2111o_1 _11224_ (.A1(net835),
    .A2(_05895_),
    .B1(_05897_),
    .C1(_05899_),
    .D1(net794),
    .X(_05900_));
 sky130_fd_sc_hd__mux2_1 _11225_ (.A0(\cpuregs[22][24] ),
    .A1(\cpuregs[23][24] ),
    .S(net687),
    .X(_05901_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(\cpuregs[20][24] ),
    .A1(\cpuregs[21][24] ),
    .S(net687),
    .X(_05902_));
 sky130_fd_sc_hd__mux2_1 _11227_ (.A0(_05901_),
    .A1(_05902_),
    .S(net818),
    .X(_05903_));
 sky130_fd_sc_hd__or2_1 _11228_ (.A(\cpuregs[16][24] ),
    .B(net699),
    .X(_05904_));
 sky130_fd_sc_hd__o211a_1 _11229_ (.A1(\cpuregs[17][24] ),
    .A2(net640),
    .B1(net614),
    .C1(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__o21a_1 _11230_ (.A1(\cpuregs[19][24] ),
    .A2(net640),
    .B1(net601),
    .X(_05906_));
 sky130_fd_sc_hd__o22a_1 _11231_ (.A1(\cpuregs[18][24] ),
    .A2(net555),
    .B1(_05906_),
    .B2(net786),
    .X(_05907_));
 sky130_fd_sc_hd__a211o_1 _11232_ (.A1(net835),
    .A2(_05903_),
    .B1(_05905_),
    .C1(_05907_),
    .X(_05908_));
 sky130_fd_sc_hd__and3_1 _11233_ (.A(net775),
    .B(_05900_),
    .C(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(\cpuregs[6][24] ),
    .A1(\cpuregs[7][24] ),
    .S(net699),
    .X(_05910_));
 sky130_fd_sc_hd__or2_1 _11235_ (.A(\cpuregs[4][24] ),
    .B(net699),
    .X(_05911_));
 sky130_fd_sc_hd__o211a_1 _11236_ (.A1(\cpuregs[5][24] ),
    .A2(net642),
    .B1(net819),
    .C1(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__a211o_1 _11237_ (.A1(net808),
    .A2(_05910_),
    .B1(_05912_),
    .C1(net839),
    .X(_05913_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(\cpuregs[2][24] ),
    .A1(\cpuregs[3][24] ),
    .S(net699),
    .X(_05914_));
 sky130_fd_sc_hd__a221o_1 _11239_ (.A1(\cpuregs[1][24] ),
    .A2(net551),
    .B1(_05914_),
    .B2(net807),
    .C1(net836),
    .X(_05915_));
 sky130_fd_sc_hd__a21o_1 _11240_ (.A1(_05913_),
    .A2(_05915_),
    .B1(net785),
    .X(_05916_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(\cpuregs[14][24] ),
    .A1(\cpuregs[15][24] ),
    .S(net686),
    .X(_05917_));
 sky130_fd_sc_hd__mux2_1 _11242_ (.A0(\cpuregs[12][24] ),
    .A1(\cpuregs[13][24] ),
    .S(net686),
    .X(_05918_));
 sky130_fd_sc_hd__or2_1 _11243_ (.A(net804),
    .B(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__o211a_1 _11244_ (.A1(net818),
    .A2(_05917_),
    .B1(_05919_),
    .C1(net834),
    .X(_05920_));
 sky130_fd_sc_hd__or2_1 _11245_ (.A(\cpuregs[8][24] ),
    .B(net686),
    .X(_05921_));
 sky130_fd_sc_hd__o211a_1 _11246_ (.A1(\cpuregs[9][24] ),
    .A2(net634),
    .B1(net611),
    .C1(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__or2_1 _11247_ (.A(\cpuregs[10][24] ),
    .B(net686),
    .X(_05923_));
 sky130_fd_sc_hd__o211a_1 _11248_ (.A1(\cpuregs[11][24] ),
    .A2(net634),
    .B1(net597),
    .C1(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__o41a_1 _11249_ (.A1(net792),
    .A2(_05920_),
    .A3(_05922_),
    .A4(_05924_),
    .B1(net778),
    .X(_05925_));
 sky130_fd_sc_hd__a21oi_2 _11250_ (.A1(_05916_),
    .A2(_05925_),
    .B1(_05909_),
    .Y(_05926_));
 sky130_fd_sc_hd__nor2_1 _11251_ (.A(net1080),
    .B(\decoded_imm[24] ),
    .Y(_05927_));
 sky130_fd_sc_hd__a211o_1 _11252_ (.A1(net1081),
    .A2(_05926_),
    .B1(_05927_),
    .C1(net858),
    .X(_05928_));
 sky130_fd_sc_hd__o21ai_1 _11253_ (.A1(_02396_),
    .A2(_05133_),
    .B1(_05928_),
    .Y(_00803_));
 sky130_fd_sc_hd__mux2_1 _11254_ (.A0(\cpuregs[6][25] ),
    .A1(\cpuregs[7][25] ),
    .S(net706),
    .X(_05929_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(\cpuregs[4][25] ),
    .A1(\cpuregs[5][25] ),
    .S(net702),
    .X(_05930_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(_05929_),
    .A1(_05930_),
    .S(net820),
    .X(_05931_));
 sky130_fd_sc_hd__or2_1 _11257_ (.A(\cpuregs[0][25] ),
    .B(net702),
    .X(_05932_));
 sky130_fd_sc_hd__o211a_1 _11258_ (.A1(\cpuregs[1][25] ),
    .A2(net642),
    .B1(net615),
    .C1(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__or2_1 _11259_ (.A(\cpuregs[2][25] ),
    .B(net699),
    .X(_05934_));
 sky130_fd_sc_hd__o211a_1 _11260_ (.A1(\cpuregs[3][25] ),
    .A2(net642),
    .B1(net602),
    .C1(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__a211o_1 _11261_ (.A1(net836),
    .A2(_05931_),
    .B1(_05935_),
    .C1(net786),
    .X(_05936_));
 sky130_fd_sc_hd__mux2_1 _11262_ (.A0(\cpuregs[14][25] ),
    .A1(\cpuregs[15][25] ),
    .S(net703),
    .X(_05937_));
 sky130_fd_sc_hd__mux2_1 _11263_ (.A0(\cpuregs[12][25] ),
    .A1(\cpuregs[13][25] ),
    .S(net703),
    .X(_05938_));
 sky130_fd_sc_hd__or2_1 _11264_ (.A(net808),
    .B(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__o211a_1 _11265_ (.A1(net820),
    .A2(_05937_),
    .B1(_05939_),
    .C1(net836),
    .X(_05940_));
 sky130_fd_sc_hd__or2_1 _11266_ (.A(\cpuregs[8][25] ),
    .B(net703),
    .X(_05941_));
 sky130_fd_sc_hd__o211a_1 _11267_ (.A1(\cpuregs[9][25] ),
    .A2(net643),
    .B1(net615),
    .C1(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__or2_1 _11268_ (.A(\cpuregs[10][25] ),
    .B(net703),
    .X(_05943_));
 sky130_fd_sc_hd__o211a_1 _11269_ (.A1(\cpuregs[11][25] ),
    .A2(net643),
    .B1(net602),
    .C1(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__or4_1 _11270_ (.A(net794),
    .B(_05940_),
    .C(_05942_),
    .D(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__o21a_1 _11271_ (.A1(_05933_),
    .A2(_05936_),
    .B1(_03171_),
    .X(_05946_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(\cpuregs[22][25] ),
    .A1(\cpuregs[23][25] ),
    .S(net705),
    .X(_05947_));
 sky130_fd_sc_hd__mux2_1 _11273_ (.A0(\cpuregs[20][25] ),
    .A1(\cpuregs[21][25] ),
    .S(net702),
    .X(_05948_));
 sky130_fd_sc_hd__mux2_1 _11274_ (.A0(_05947_),
    .A1(_05948_),
    .S(net820),
    .X(_05949_));
 sky130_fd_sc_hd__or2_1 _11275_ (.A(\cpuregs[16][25] ),
    .B(net705),
    .X(_05950_));
 sky130_fd_sc_hd__o211a_1 _11276_ (.A1(\cpuregs[17][25] ),
    .A2(net642),
    .B1(net615),
    .C1(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__o21a_1 _11277_ (.A1(\cpuregs[19][25] ),
    .A2(net642),
    .B1(net602),
    .X(_05952_));
 sky130_fd_sc_hd__o22a_1 _11278_ (.A1(\cpuregs[18][25] ),
    .A2(net555),
    .B1(_05952_),
    .B2(net786),
    .X(_05953_));
 sky130_fd_sc_hd__a211o_1 _11279_ (.A1(net836),
    .A2(_05949_),
    .B1(_05951_),
    .C1(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__mux2_1 _11280_ (.A0(\cpuregs[28][25] ),
    .A1(\cpuregs[29][25] ),
    .S(net706),
    .X(_05955_));
 sky130_fd_sc_hd__mux2_1 _11281_ (.A0(\cpuregs[30][25] ),
    .A1(\cpuregs[31][25] ),
    .S(net704),
    .X(_05956_));
 sky130_fd_sc_hd__mux2_1 _11282_ (.A0(_05955_),
    .A1(_05956_),
    .S(net808),
    .X(_05957_));
 sky130_fd_sc_hd__or2_1 _11283_ (.A(\cpuregs[24][25] ),
    .B(net704),
    .X(_05958_));
 sky130_fd_sc_hd__o211a_1 _11284_ (.A1(\cpuregs[25][25] ),
    .A2(net644),
    .B1(net614),
    .C1(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__or2_1 _11285_ (.A(\cpuregs[26][25] ),
    .B(net704),
    .X(_05960_));
 sky130_fd_sc_hd__o211a_1 _11286_ (.A1(\cpuregs[27][25] ),
    .A2(net642),
    .B1(net602),
    .C1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__a2111o_1 _11287_ (.A1(net836),
    .A2(_05957_),
    .B1(_05959_),
    .C1(_05961_),
    .D1(net794),
    .X(_05962_));
 sky130_fd_sc_hd__and3_1 _11288_ (.A(net775),
    .B(_05954_),
    .C(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__a21oi_2 _11289_ (.A1(_05945_),
    .A2(_05946_),
    .B1(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__nand2_1 _11290_ (.A(net1083),
    .B(_05964_),
    .Y(_05965_));
 sky130_fd_sc_hd__o21a_1 _11291_ (.A1(net1083),
    .A2(\decoded_imm[25] ),
    .B1(_05133_),
    .X(_05966_));
 sky130_fd_sc_hd__a22o_1 _11292_ (.A1(net252),
    .A2(net858),
    .B1(_05965_),
    .B2(_05966_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(\cpuregs[6][26] ),
    .A1(\cpuregs[7][26] ),
    .S(net702),
    .X(_05967_));
 sky130_fd_sc_hd__mux2_1 _11294_ (.A0(\cpuregs[4][26] ),
    .A1(\cpuregs[5][26] ),
    .S(net702),
    .X(_05968_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(_05967_),
    .A1(_05968_),
    .S(net819),
    .X(_05969_));
 sky130_fd_sc_hd__mux2_1 _11296_ (.A0(\cpuregs[2][26] ),
    .A1(\cpuregs[3][26] ),
    .S(net702),
    .X(_05970_));
 sky130_fd_sc_hd__a221o_1 _11297_ (.A1(\cpuregs[1][26] ),
    .A2(net551),
    .B1(_05970_),
    .B2(net807),
    .C1(net836),
    .X(_05971_));
 sky130_fd_sc_hd__o21a_1 _11298_ (.A1(net840),
    .A2(_05969_),
    .B1(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(\cpuregs[12][26] ),
    .A1(\cpuregs[13][26] ),
    .S(net703),
    .X(_05973_));
 sky130_fd_sc_hd__mux2_1 _11300_ (.A0(\cpuregs[14][26] ),
    .A1(\cpuregs[15][26] ),
    .S(net704),
    .X(_05974_));
 sky130_fd_sc_hd__or2_1 _11301_ (.A(net820),
    .B(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__o211a_1 _11302_ (.A1(net807),
    .A2(_05973_),
    .B1(_05975_),
    .C1(net836),
    .X(_05976_));
 sky130_fd_sc_hd__or2_1 _11303_ (.A(\cpuregs[8][26] ),
    .B(net703),
    .X(_05977_));
 sky130_fd_sc_hd__o211a_1 _11304_ (.A1(\cpuregs[9][26] ),
    .A2(net643),
    .B1(net615),
    .C1(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__or2_1 _11305_ (.A(\cpuregs[10][26] ),
    .B(net694),
    .X(_05979_));
 sky130_fd_sc_hd__o211a_1 _11306_ (.A1(\cpuregs[11][26] ),
    .A2(net643),
    .B1(net601),
    .C1(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__or4_1 _11307_ (.A(net794),
    .B(_05976_),
    .C(_05978_),
    .D(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__o211a_1 _11308_ (.A1(net785),
    .A2(_05972_),
    .B1(_05981_),
    .C1(net778),
    .X(_05982_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(\cpuregs[28][26] ),
    .A1(\cpuregs[29][26] ),
    .S(net703),
    .X(_05983_));
 sky130_fd_sc_hd__mux2_1 _11310_ (.A0(\cpuregs[30][26] ),
    .A1(\cpuregs[31][26] ),
    .S(net703),
    .X(_05984_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(_05983_),
    .A1(_05984_),
    .S(net807),
    .X(_05985_));
 sky130_fd_sc_hd__or2_1 _11312_ (.A(\cpuregs[24][26] ),
    .B(net703),
    .X(_05986_));
 sky130_fd_sc_hd__o211a_1 _11313_ (.A1(\cpuregs[25][26] ),
    .A2(net643),
    .B1(net615),
    .C1(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__or2_1 _11314_ (.A(\cpuregs[26][26] ),
    .B(net703),
    .X(_05988_));
 sky130_fd_sc_hd__o211a_1 _11315_ (.A1(\cpuregs[27][26] ),
    .A2(net642),
    .B1(net601),
    .C1(_05988_),
    .X(_05989_));
 sky130_fd_sc_hd__a2111o_1 _11316_ (.A1(net836),
    .A2(_05985_),
    .B1(_05987_),
    .C1(_05989_),
    .D1(net794),
    .X(_05990_));
 sky130_fd_sc_hd__mux2_1 _11317_ (.A0(\cpuregs[22][26] ),
    .A1(\cpuregs[23][26] ),
    .S(net702),
    .X(_05991_));
 sky130_fd_sc_hd__mux2_1 _11318_ (.A0(\cpuregs[20][26] ),
    .A1(\cpuregs[21][26] ),
    .S(net702),
    .X(_05992_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(_05991_),
    .A1(_05992_),
    .S(net820),
    .X(_05993_));
 sky130_fd_sc_hd__or2_1 _11320_ (.A(\cpuregs[16][26] ),
    .B(net702),
    .X(_05994_));
 sky130_fd_sc_hd__o211a_1 _11321_ (.A1(\cpuregs[17][26] ),
    .A2(net642),
    .B1(net615),
    .C1(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__o21a_1 _11322_ (.A1(\cpuregs[19][26] ),
    .A2(net642),
    .B1(net602),
    .X(_05996_));
 sky130_fd_sc_hd__o22a_1 _11323_ (.A1(\cpuregs[18][26] ),
    .A2(net555),
    .B1(_05996_),
    .B2(net786),
    .X(_05997_));
 sky130_fd_sc_hd__a211o_1 _11324_ (.A1(net836),
    .A2(_05993_),
    .B1(_05995_),
    .C1(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__a31oi_4 _11325_ (.A1(net775),
    .A2(_05990_),
    .A3(_05998_),
    .B1(_05982_),
    .Y(_05999_));
 sky130_fd_sc_hd__or2_1 _11326_ (.A(net1083),
    .B(\decoded_imm[26] ),
    .X(_06000_));
 sky130_fd_sc_hd__a21oi_1 _11327_ (.A1(net1083),
    .A2(_05999_),
    .B1(net857),
    .Y(_06001_));
 sky130_fd_sc_hd__a22o_1 _11328_ (.A1(net253),
    .A2(net857),
    .B1(_06000_),
    .B2(_06001_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _11329_ (.A0(\cpuregs[6][27] ),
    .A1(\cpuregs[7][27] ),
    .S(net695),
    .X(_06002_));
 sky130_fd_sc_hd__mux2_1 _11330_ (.A0(\cpuregs[4][27] ),
    .A1(\cpuregs[5][27] ),
    .S(net695),
    .X(_06003_));
 sky130_fd_sc_hd__mux2_1 _11331_ (.A0(_06002_),
    .A1(_06003_),
    .S(net817),
    .X(_06004_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(\cpuregs[2][27] ),
    .A1(\cpuregs[3][27] ),
    .S(net692),
    .X(_06005_));
 sky130_fd_sc_hd__a221o_1 _11333_ (.A1(\cpuregs[1][27] ),
    .A2(net551),
    .B1(_06005_),
    .B2(net806),
    .C1(net833),
    .X(_06006_));
 sky130_fd_sc_hd__o21a_1 _11334_ (.A1(net840),
    .A2(_06004_),
    .B1(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__mux2_1 _11335_ (.A0(\cpuregs[14][27] ),
    .A1(\cpuregs[15][27] ),
    .S(net693),
    .X(_06008_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(\cpuregs[12][27] ),
    .A1(\cpuregs[13][27] ),
    .S(net693),
    .X(_06009_));
 sky130_fd_sc_hd__or2_1 _11337_ (.A(net805),
    .B(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__o211a_1 _11338_ (.A1(net817),
    .A2(_06008_),
    .B1(_06010_),
    .C1(net833),
    .X(_06011_));
 sky130_fd_sc_hd__or2_1 _11339_ (.A(\cpuregs[8][27] ),
    .B(net693),
    .X(_06012_));
 sky130_fd_sc_hd__o211a_1 _11340_ (.A1(\cpuregs[9][27] ),
    .A2(net638),
    .B1(net613),
    .C1(_06012_),
    .X(_06013_));
 sky130_fd_sc_hd__or2_1 _11341_ (.A(\cpuregs[10][27] ),
    .B(net693),
    .X(_06014_));
 sky130_fd_sc_hd__o211a_1 _11342_ (.A1(\cpuregs[11][27] ),
    .A2(net639),
    .B1(net598),
    .C1(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__or4_1 _11343_ (.A(net793),
    .B(_06011_),
    .C(_06013_),
    .D(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__o211a_1 _11344_ (.A1(net783),
    .A2(_06007_),
    .B1(_06016_),
    .C1(net778),
    .X(_06017_));
 sky130_fd_sc_hd__mux2_1 _11345_ (.A0(\cpuregs[28][27] ),
    .A1(\cpuregs[29][27] ),
    .S(net694),
    .X(_06018_));
 sky130_fd_sc_hd__mux2_1 _11346_ (.A0(\cpuregs[30][27] ),
    .A1(\cpuregs[31][27] ),
    .S(net694),
    .X(_06019_));
 sky130_fd_sc_hd__mux2_1 _11347_ (.A0(_06018_),
    .A1(_06019_),
    .S(net806),
    .X(_06020_));
 sky130_fd_sc_hd__or2_1 _11348_ (.A(\cpuregs[24][27] ),
    .B(net693),
    .X(_06021_));
 sky130_fd_sc_hd__o211a_1 _11349_ (.A1(\cpuregs[25][27] ),
    .A2(net639),
    .B1(net613),
    .C1(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__or2_1 _11350_ (.A(\cpuregs[26][27] ),
    .B(net693),
    .X(_06023_));
 sky130_fd_sc_hd__o211a_1 _11351_ (.A1(\cpuregs[27][27] ),
    .A2(net639),
    .B1(net599),
    .C1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__a2111o_1 _11352_ (.A1(net833),
    .A2(_06020_),
    .B1(_06022_),
    .C1(_06024_),
    .D1(net793),
    .X(_06025_));
 sky130_fd_sc_hd__mux2_1 _11353_ (.A0(\cpuregs[20][27] ),
    .A1(\cpuregs[21][27] ),
    .S(net692),
    .X(_06026_));
 sky130_fd_sc_hd__mux2_1 _11354_ (.A0(\cpuregs[22][27] ),
    .A1(\cpuregs[23][27] ),
    .S(net692),
    .X(_06027_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(_06026_),
    .A1(_06027_),
    .S(net805),
    .X(_06028_));
 sky130_fd_sc_hd__or2_1 _11356_ (.A(\cpuregs[16][27] ),
    .B(net692),
    .X(_06029_));
 sky130_fd_sc_hd__o211a_1 _11357_ (.A1(\cpuregs[17][27] ),
    .A2(net638),
    .B1(net613),
    .C1(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__o21a_1 _11358_ (.A1(\cpuregs[19][27] ),
    .A2(net638),
    .B1(net599),
    .X(_06031_));
 sky130_fd_sc_hd__o22a_1 _11359_ (.A1(\cpuregs[18][27] ),
    .A2(net554),
    .B1(_06031_),
    .B2(net784),
    .X(_06032_));
 sky130_fd_sc_hd__a211o_1 _11360_ (.A1(net833),
    .A2(_06028_),
    .B1(_06030_),
    .C1(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__a31oi_4 _11361_ (.A1(net774),
    .A2(_06025_),
    .A3(_06033_),
    .B1(_06017_),
    .Y(_06034_));
 sky130_fd_sc_hd__nor2_1 _11362_ (.A(net1081),
    .B(\decoded_imm[27] ),
    .Y(_06035_));
 sky130_fd_sc_hd__a211o_1 _11363_ (.A1(net1081),
    .A2(_06034_),
    .B1(_06035_),
    .C1(net858),
    .X(_06036_));
 sky130_fd_sc_hd__o21ai_1 _11364_ (.A1(_02397_),
    .A2(net860),
    .B1(_06036_),
    .Y(_00806_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(\cpuregs[6][28] ),
    .A1(\cpuregs[7][28] ),
    .S(net692),
    .X(_06037_));
 sky130_fd_sc_hd__mux2_1 _11366_ (.A0(\cpuregs[4][28] ),
    .A1(\cpuregs[5][28] ),
    .S(net692),
    .X(_06038_));
 sky130_fd_sc_hd__mux2_1 _11367_ (.A0(_06037_),
    .A1(_06038_),
    .S(net817),
    .X(_06039_));
 sky130_fd_sc_hd__mux2_1 _11368_ (.A0(\cpuregs[2][28] ),
    .A1(\cpuregs[3][28] ),
    .S(net691),
    .X(_06040_));
 sky130_fd_sc_hd__a221o_1 _11369_ (.A1(\cpuregs[1][28] ),
    .A2(net551),
    .B1(_06040_),
    .B2(net805),
    .C1(net832),
    .X(_06041_));
 sky130_fd_sc_hd__o21a_1 _11370_ (.A1(net840),
    .A2(_06039_),
    .B1(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__mux2_1 _11371_ (.A0(\cpuregs[14][28] ),
    .A1(\cpuregs[15][28] ),
    .S(net689),
    .X(_06043_));
 sky130_fd_sc_hd__mux2_1 _11372_ (.A0(\cpuregs[12][28] ),
    .A1(\cpuregs[13][28] ),
    .S(net689),
    .X(_06044_));
 sky130_fd_sc_hd__or2_1 _11373_ (.A(net805),
    .B(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__o211a_1 _11374_ (.A1(net817),
    .A2(_06043_),
    .B1(_06045_),
    .C1(net832),
    .X(_06046_));
 sky130_fd_sc_hd__or2_1 _11375_ (.A(\cpuregs[8][28] ),
    .B(net689),
    .X(_06047_));
 sky130_fd_sc_hd__o211a_1 _11376_ (.A1(\cpuregs[9][28] ),
    .A2(net637),
    .B1(net612),
    .C1(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__or2_1 _11377_ (.A(\cpuregs[10][28] ),
    .B(net689),
    .X(_06049_));
 sky130_fd_sc_hd__o211a_1 _11378_ (.A1(\cpuregs[11][28] ),
    .A2(net637),
    .B1(net598),
    .C1(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__or4_1 _11379_ (.A(net793),
    .B(_06046_),
    .C(_06048_),
    .D(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__o211a_1 _11380_ (.A1(net783),
    .A2(_06042_),
    .B1(_06051_),
    .C1(net778),
    .X(_06052_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(\cpuregs[28][28] ),
    .A1(\cpuregs[29][28] ),
    .S(net690),
    .X(_06053_));
 sky130_fd_sc_hd__mux2_1 _11382_ (.A0(\cpuregs[30][28] ),
    .A1(\cpuregs[31][28] ),
    .S(net690),
    .X(_06054_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(_06053_),
    .A1(_06054_),
    .S(net805),
    .X(_06055_));
 sky130_fd_sc_hd__or2_1 _11384_ (.A(\cpuregs[24][28] ),
    .B(net689),
    .X(_06056_));
 sky130_fd_sc_hd__o211a_1 _11385_ (.A1(\cpuregs[25][28] ),
    .A2(net637),
    .B1(net612),
    .C1(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__or2_1 _11386_ (.A(\cpuregs[26][28] ),
    .B(net690),
    .X(_06058_));
 sky130_fd_sc_hd__o211a_1 _11387_ (.A1(\cpuregs[27][28] ),
    .A2(net637),
    .B1(net598),
    .C1(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__a2111o_1 _11388_ (.A1(net832),
    .A2(_06055_),
    .B1(_06057_),
    .C1(_06059_),
    .D1(net793),
    .X(_06060_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(\cpuregs[22][28] ),
    .A1(\cpuregs[23][28] ),
    .S(net688),
    .X(_06061_));
 sky130_fd_sc_hd__mux2_1 _11390_ (.A0(\cpuregs[20][28] ),
    .A1(\cpuregs[21][28] ),
    .S(net688),
    .X(_06062_));
 sky130_fd_sc_hd__mux2_1 _11391_ (.A0(_06061_),
    .A1(_06062_),
    .S(net817),
    .X(_06063_));
 sky130_fd_sc_hd__or2_1 _11392_ (.A(\cpuregs[16][28] ),
    .B(net688),
    .X(_06064_));
 sky130_fd_sc_hd__o211a_1 _11393_ (.A1(\cpuregs[17][28] ),
    .A2(net636),
    .B1(net612),
    .C1(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__o21a_1 _11394_ (.A1(\cpuregs[19][28] ),
    .A2(net636),
    .B1(net598),
    .X(_06066_));
 sky130_fd_sc_hd__o22a_1 _11395_ (.A1(\cpuregs[18][28] ),
    .A2(net554),
    .B1(_06066_),
    .B2(net783),
    .X(_06067_));
 sky130_fd_sc_hd__a211o_1 _11396_ (.A1(net832),
    .A2(_06063_),
    .B1(_06065_),
    .C1(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__a31oi_4 _11397_ (.A1(net774),
    .A2(_06060_),
    .A3(_06068_),
    .B1(_06052_),
    .Y(_06069_));
 sky130_fd_sc_hd__or2_1 _11398_ (.A(net1081),
    .B(\decoded_imm[28] ),
    .X(_06070_));
 sky130_fd_sc_hd__a21oi_1 _11399_ (.A1(net1083),
    .A2(_06069_),
    .B1(net857),
    .Y(_06071_));
 sky130_fd_sc_hd__a22o_1 _11400_ (.A1(net255),
    .A2(net857),
    .B1(_06070_),
    .B2(_06071_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _11401_ (.A0(\cpuregs[6][29] ),
    .A1(\cpuregs[7][29] ),
    .S(net706),
    .X(_06072_));
 sky130_fd_sc_hd__or2_1 _11402_ (.A(\cpuregs[4][29] ),
    .B(net706),
    .X(_06073_));
 sky130_fd_sc_hd__o211a_1 _11403_ (.A1(\cpuregs[5][29] ),
    .A2(net644),
    .B1(net820),
    .C1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__a211o_1 _11404_ (.A1(net808),
    .A2(_06072_),
    .B1(_06074_),
    .C1(net839),
    .X(_06075_));
 sky130_fd_sc_hd__mux2_1 _11405_ (.A0(\cpuregs[2][29] ),
    .A1(\cpuregs[3][29] ),
    .S(net705),
    .X(_06076_));
 sky130_fd_sc_hd__a221o_1 _11406_ (.A1(\cpuregs[1][29] ),
    .A2(net551),
    .B1(_06076_),
    .B2(net808),
    .C1(net837),
    .X(_06077_));
 sky130_fd_sc_hd__a21o_1 _11407_ (.A1(_06075_),
    .A2(_06077_),
    .B1(net786),
    .X(_06078_));
 sky130_fd_sc_hd__mux2_1 _11408_ (.A0(\cpuregs[14][29] ),
    .A1(\cpuregs[15][29] ),
    .S(net704),
    .X(_06079_));
 sky130_fd_sc_hd__mux2_1 _11409_ (.A0(\cpuregs[12][29] ),
    .A1(\cpuregs[13][29] ),
    .S(net704),
    .X(_06080_));
 sky130_fd_sc_hd__or2_1 _11410_ (.A(net808),
    .B(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__o211a_1 _11411_ (.A1(net819),
    .A2(_06079_),
    .B1(_06081_),
    .C1(net836),
    .X(_06082_));
 sky130_fd_sc_hd__or2_1 _11412_ (.A(\cpuregs[8][29] ),
    .B(net704),
    .X(_06083_));
 sky130_fd_sc_hd__o211a_1 _11413_ (.A1(\cpuregs[9][29] ),
    .A2(net643),
    .B1(net615),
    .C1(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__or2_1 _11414_ (.A(\cpuregs[10][29] ),
    .B(net702),
    .X(_06085_));
 sky130_fd_sc_hd__o211a_1 _11415_ (.A1(\cpuregs[11][29] ),
    .A2(net642),
    .B1(net602),
    .C1(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__o41a_1 _11416_ (.A1(net795),
    .A2(_06082_),
    .A3(_06084_),
    .A4(_06086_),
    .B1(net778),
    .X(_06087_));
 sky130_fd_sc_hd__mux2_1 _11417_ (.A0(\cpuregs[30][29] ),
    .A1(\cpuregs[31][29] ),
    .S(net706),
    .X(_06088_));
 sky130_fd_sc_hd__mux2_1 _11418_ (.A0(\cpuregs[28][29] ),
    .A1(\cpuregs[29][29] ),
    .S(net706),
    .X(_06089_));
 sky130_fd_sc_hd__mux2_1 _11419_ (.A0(_06088_),
    .A1(_06089_),
    .S(net820),
    .X(_06090_));
 sky130_fd_sc_hd__or2_1 _11420_ (.A(\cpuregs[24][29] ),
    .B(net706),
    .X(_06091_));
 sky130_fd_sc_hd__o211a_1 _11421_ (.A1(\cpuregs[25][29] ),
    .A2(net644),
    .B1(net615),
    .C1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__or2_1 _11422_ (.A(\cpuregs[26][29] ),
    .B(net707),
    .X(_06093_));
 sky130_fd_sc_hd__o211a_1 _11423_ (.A1(\cpuregs[27][29] ),
    .A2(net644),
    .B1(net602),
    .C1(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__a2111o_1 _11424_ (.A1(net837),
    .A2(_06090_),
    .B1(_06092_),
    .C1(_06094_),
    .D1(net794),
    .X(_06095_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(\cpuregs[20][29] ),
    .A1(\cpuregs[21][29] ),
    .S(net706),
    .X(_06096_));
 sky130_fd_sc_hd__mux2_1 _11426_ (.A0(\cpuregs[22][29] ),
    .A1(\cpuregs[23][29] ),
    .S(net706),
    .X(_06097_));
 sky130_fd_sc_hd__mux2_1 _11427_ (.A0(_06096_),
    .A1(_06097_),
    .S(net808),
    .X(_06098_));
 sky130_fd_sc_hd__or2_1 _11428_ (.A(\cpuregs[16][29] ),
    .B(net706),
    .X(_06099_));
 sky130_fd_sc_hd__o211a_1 _11429_ (.A1(\cpuregs[17][29] ),
    .A2(net644),
    .B1(net615),
    .C1(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__o21a_1 _11430_ (.A1(\cpuregs[19][29] ),
    .A2(net644),
    .B1(net602),
    .X(_06101_));
 sky130_fd_sc_hd__o22a_1 _11431_ (.A1(\cpuregs[18][29] ),
    .A2(net555),
    .B1(_06101_),
    .B2(net786),
    .X(_06102_));
 sky130_fd_sc_hd__a211o_1 _11432_ (.A1(net837),
    .A2(_06098_),
    .B1(_06100_),
    .C1(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__and3_1 _11433_ (.A(net775),
    .B(_06095_),
    .C(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__a21oi_2 _11434_ (.A1(_06078_),
    .A2(_06087_),
    .B1(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__or2_1 _11435_ (.A(net1081),
    .B(\decoded_imm[29] ),
    .X(_06106_));
 sky130_fd_sc_hd__a21oi_1 _11436_ (.A1(net1083),
    .A2(_06105_),
    .B1(net857),
    .Y(_06107_));
 sky130_fd_sc_hd__a22o_1 _11437_ (.A1(net256),
    .A2(net857),
    .B1(_06106_),
    .B2(_06107_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _11438_ (.A0(\cpuregs[6][30] ),
    .A1(\cpuregs[7][30] ),
    .S(net692),
    .X(_06108_));
 sky130_fd_sc_hd__mux2_1 _11439_ (.A0(\cpuregs[4][30] ),
    .A1(\cpuregs[5][30] ),
    .S(net688),
    .X(_06109_));
 sky130_fd_sc_hd__mux2_1 _11440_ (.A0(_06108_),
    .A1(_06109_),
    .S(net817),
    .X(_06110_));
 sky130_fd_sc_hd__or2_1 _11441_ (.A(\cpuregs[0][30] ),
    .B(net691),
    .X(_06111_));
 sky130_fd_sc_hd__o211a_1 _11442_ (.A1(\cpuregs[1][30] ),
    .A2(net637),
    .B1(net612),
    .C1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__or2_1 _11443_ (.A(\cpuregs[2][30] ),
    .B(net691),
    .X(_06113_));
 sky130_fd_sc_hd__o211a_1 _11444_ (.A1(\cpuregs[3][30] ),
    .A2(net636),
    .B1(net598),
    .C1(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__a211o_1 _11445_ (.A1(net832),
    .A2(_06110_),
    .B1(_06114_),
    .C1(net783),
    .X(_06115_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(\cpuregs[12][30] ),
    .A1(\cpuregs[13][30] ),
    .S(net689),
    .X(_06116_));
 sky130_fd_sc_hd__mux2_1 _11447_ (.A0(\cpuregs[14][30] ),
    .A1(\cpuregs[15][30] ),
    .S(net689),
    .X(_06117_));
 sky130_fd_sc_hd__or2_1 _11448_ (.A(net817),
    .B(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__o211a_1 _11449_ (.A1(net805),
    .A2(_06116_),
    .B1(_06118_),
    .C1(net833),
    .X(_06119_));
 sky130_fd_sc_hd__or2_1 _11450_ (.A(\cpuregs[8][30] ),
    .B(net689),
    .X(_06120_));
 sky130_fd_sc_hd__o211a_1 _11451_ (.A1(\cpuregs[9][30] ),
    .A2(net637),
    .B1(net612),
    .C1(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__or2_1 _11452_ (.A(\cpuregs[10][30] ),
    .B(net689),
    .X(_06122_));
 sky130_fd_sc_hd__o211a_1 _11453_ (.A1(\cpuregs[11][30] ),
    .A2(net637),
    .B1(net598),
    .C1(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__or4_2 _11454_ (.A(net793),
    .B(_06119_),
    .C(_06121_),
    .D(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__o21a_1 _11455_ (.A1(_06112_),
    .A2(_06115_),
    .B1(_03171_),
    .X(_06125_));
 sky130_fd_sc_hd__mux2_1 _11456_ (.A0(\cpuregs[20][30] ),
    .A1(\cpuregs[21][30] ),
    .S(net688),
    .X(_06126_));
 sky130_fd_sc_hd__mux2_1 _11457_ (.A0(\cpuregs[22][30] ),
    .A1(\cpuregs[23][30] ),
    .S(net689),
    .X(_06127_));
 sky130_fd_sc_hd__mux2_1 _11458_ (.A0(_06126_),
    .A1(_06127_),
    .S(net805),
    .X(_06128_));
 sky130_fd_sc_hd__or2_1 _11459_ (.A(\cpuregs[16][30] ),
    .B(net688),
    .X(_06129_));
 sky130_fd_sc_hd__o211a_1 _11460_ (.A1(\cpuregs[17][30] ),
    .A2(net636),
    .B1(net612),
    .C1(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__o21a_1 _11461_ (.A1(\cpuregs[19][30] ),
    .A2(net636),
    .B1(net598),
    .X(_06131_));
 sky130_fd_sc_hd__o22a_1 _11462_ (.A1(\cpuregs[18][30] ),
    .A2(net554),
    .B1(_06131_),
    .B2(net783),
    .X(_06132_));
 sky130_fd_sc_hd__a211o_1 _11463_ (.A1(net832),
    .A2(_06128_),
    .B1(_06130_),
    .C1(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__mux2_1 _11464_ (.A0(\cpuregs[28][30] ),
    .A1(\cpuregs[29][30] ),
    .S(net690),
    .X(_06134_));
 sky130_fd_sc_hd__mux2_1 _11465_ (.A0(\cpuregs[30][30] ),
    .A1(\cpuregs[31][30] ),
    .S(net690),
    .X(_06135_));
 sky130_fd_sc_hd__mux2_1 _11466_ (.A0(_06134_),
    .A1(_06135_),
    .S(net805),
    .X(_06136_));
 sky130_fd_sc_hd__or2_1 _11467_ (.A(\cpuregs[24][30] ),
    .B(net690),
    .X(_06137_));
 sky130_fd_sc_hd__o211a_1 _11468_ (.A1(\cpuregs[25][30] ),
    .A2(net637),
    .B1(net612),
    .C1(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__or2_1 _11469_ (.A(\cpuregs[26][30] ),
    .B(net690),
    .X(_06139_));
 sky130_fd_sc_hd__o211a_1 _11470_ (.A1(\cpuregs[27][30] ),
    .A2(net637),
    .B1(net598),
    .C1(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__a2111o_1 _11471_ (.A1(net832),
    .A2(_06136_),
    .B1(_06138_),
    .C1(_06140_),
    .D1(net793),
    .X(_06141_));
 sky130_fd_sc_hd__and3_1 _11472_ (.A(net774),
    .B(_06133_),
    .C(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__a21oi_4 _11473_ (.A1(_06124_),
    .A2(_06125_),
    .B1(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__or2_1 _11474_ (.A(net1083),
    .B(\decoded_imm[30] ),
    .X(_06144_));
 sky130_fd_sc_hd__a21oi_1 _11475_ (.A1(net1083),
    .A2(_06143_),
    .B1(net857),
    .Y(_06145_));
 sky130_fd_sc_hd__a22o_1 _11476_ (.A1(net258),
    .A2(net857),
    .B1(_06144_),
    .B2(_06145_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _11477_ (.A(net1084),
    .B(\decoded_imm[31] ),
    .X(_06146_));
 sky130_fd_sc_hd__a21oi_1 _11478_ (.A1(net1084),
    .A2(_05076_),
    .B1(net857),
    .Y(_06147_));
 sky130_fd_sc_hd__a22o_1 _11479_ (.A1(net1157),
    .A2(net857),
    .B1(_06146_),
    .B2(_06147_),
    .X(_00810_));
 sky130_fd_sc_hd__o21a_1 _11480_ (.A1(_02436_),
    .A2(_02438_),
    .B1(net1084),
    .X(_06148_));
 sky130_fd_sc_hd__nor2_1 _11481_ (.A(net1072),
    .B(net1089),
    .Y(_06149_));
 sky130_fd_sc_hd__or2_1 _11482_ (.A(net1072),
    .B(net1089),
    .X(_06150_));
 sky130_fd_sc_hd__and3b_1 _11483_ (.A_N(_05125_),
    .B(_06149_),
    .C(_02387_),
    .X(_06151_));
 sky130_fd_sc_hd__a211o_1 _11484_ (.A1(\cpu_state[2] ),
    .A2(_02471_),
    .B1(_06148_),
    .C1(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__or4_1 _11485_ (.A(net1061),
    .B(_02487_),
    .C(_05125_),
    .D(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__a21oi_1 _11486_ (.A1(_02368_),
    .A2(_06152_),
    .B1(net1208),
    .Y(_06154_));
 sky130_fd_sc_hd__o21a_1 _11487_ (.A1(_03739_),
    .A2(_06153_),
    .B1(_06154_),
    .X(_00811_));
 sky130_fd_sc_hd__o221a_1 _11488_ (.A1(net1072),
    .A2(_02370_),
    .B1(_02487_),
    .B2(net1156),
    .C1(net1232),
    .X(_00812_));
 sky130_fd_sc_hd__a221o_1 _11489_ (.A1(net991),
    .A2(_02480_),
    .B1(_02487_),
    .B2(instr_jalr),
    .C1(_06149_),
    .X(_06155_));
 sky130_fd_sc_hd__o221a_1 _11490_ (.A1(latched_branch),
    .A2(_06150_),
    .B1(_06155_),
    .B2(_03740_),
    .C1(net1232),
    .X(_00813_));
 sky130_fd_sc_hd__o221a_1 _11491_ (.A1(_02370_),
    .A2(net1061),
    .B1(_02454_),
    .B2(mem_do_rdata),
    .C1(net1232),
    .X(_06156_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(instr_lh),
    .A2(_02455_),
    .B1(_06156_),
    .B2(net3026),
    .X(_00815_));
 sky130_fd_sc_hd__a22o_1 _11493_ (.A1(net3036),
    .A2(_02455_),
    .B1(_06156_),
    .B2(latched_is_lb),
    .X(_00816_));
 sky130_fd_sc_hd__or4bb_1 _11494_ (.A(\genblk2.pcpi_div.pcpi_wait ),
    .B(\genblk1.genblk1.pcpi_mul.pcpi_wait ),
    .C_N(net267),
    .D_N(net1237),
    .X(_06157_));
 sky130_fd_sc_hd__or3_1 _11495_ (.A(\pcpi_timeout_counter[2] ),
    .B(\pcpi_timeout_counter[1] ),
    .C(\pcpi_timeout_counter[0] ),
    .X(_06158_));
 sky130_fd_sc_hd__inv_2 _11496_ (.A(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__nor2_1 _11497_ (.A(net2542),
    .B(_06158_),
    .Y(_06160_));
 sky130_fd_sc_hd__o21bai_1 _11498_ (.A1(net2850),
    .A2(_06160_),
    .B1_N(_06157_),
    .Y(_00817_));
 sky130_fd_sc_hd__nor3_1 _11499_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .C(_06160_),
    .Y(_06161_));
 sky130_fd_sc_hd__a211o_1 _11500_ (.A1(net2861),
    .A2(net2850),
    .B1(_06157_),
    .C1(_06161_),
    .X(_00818_));
 sky130_fd_sc_hd__o21a_1 _11501_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(net2606),
    .X(_06162_));
 sky130_fd_sc_hd__a211o_1 _11502_ (.A1(net2542),
    .A2(_06159_),
    .B1(_06162_),
    .C1(_06157_),
    .X(_00819_));
 sky130_fd_sc_hd__a21o_1 _11503_ (.A1(net2542),
    .A2(_06158_),
    .B1(_06157_),
    .X(_00820_));
 sky130_fd_sc_hd__and2_1 _11504_ (.A(net1240),
    .B(_06160_),
    .X(_00821_));
 sky130_fd_sc_hd__nor2_1 _11505_ (.A(_02380_),
    .B(decoder_pseudo_trigger),
    .Y(_06163_));
 sky130_fd_sc_hd__or2_1 _11506_ (.A(_02380_),
    .B(decoder_pseudo_trigger),
    .X(_06164_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(net2554),
    .A1(\mem_rdata_q[0] ),
    .S(net746),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _11508_ (.A0(net2648),
    .A1(net2645),
    .S(net747),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(net193),
    .A1(net3048),
    .S(net746),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _11510_ (.A0(net2612),
    .A1(\mem_rdata_q[3] ),
    .S(net746),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _11511_ (.A0(net2636),
    .A1(\mem_rdata_q[4] ),
    .S(net746),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _11512_ (.A0(net2980),
    .A1(\mem_rdata_q[5] ),
    .S(net746),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(net2737),
    .A1(\mem_rdata_q[6] ),
    .S(net746),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _11514_ (.A0(\mem_rdata_q[7] ),
    .A1(net2055),
    .S(net736),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(\mem_rdata_q[8] ),
    .A1(net1924),
    .S(net736),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _11516_ (.A0(\mem_rdata_q[9] ),
    .A1(net1863),
    .S(net738),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(\mem_rdata_q[10] ),
    .A1(net2042),
    .S(net737),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _11518_ (.A0(\mem_rdata_q[11] ),
    .A1(net1782),
    .S(net738),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _11519_ (.A0(\mem_rdata_q[12] ),
    .A1(net174),
    .S(net740),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _11520_ (.A0(\mem_rdata_q[13] ),
    .A1(net175),
    .S(net740),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _11521_ (.A0(\mem_rdata_q[14] ),
    .A1(net3049),
    .S(net740),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _11522_ (.A0(\mem_rdata_q[15] ),
    .A1(net2238),
    .S(net742),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _11523_ (.A0(\mem_rdata_q[16] ),
    .A1(net1973),
    .S(net742),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _11524_ (.A0(\mem_rdata_q[17] ),
    .A1(net2109),
    .S(net742),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _11525_ (.A0(\mem_rdata_q[18] ),
    .A1(net2611),
    .S(net742),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _11526_ (.A0(\mem_rdata_q[19] ),
    .A1(net2101),
    .S(net742),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _11527_ (.A0(\mem_rdata_q[20] ),
    .A1(net2349),
    .S(net736),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _11528_ (.A0(\mem_rdata_q[21] ),
    .A1(net1896),
    .S(net742),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _11529_ (.A0(\mem_rdata_q[22] ),
    .A1(net2423),
    .S(net742),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _11530_ (.A0(\mem_rdata_q[23] ),
    .A1(net2053),
    .S(net737),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _11531_ (.A0(\mem_rdata_q[24] ),
    .A1(net1589),
    .S(net737),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _11532_ (.A0(\mem_rdata_q[25] ),
    .A1(net2680),
    .S(net736),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _11533_ (.A0(\mem_rdata_q[26] ),
    .A1(net2684),
    .S(net736),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _11534_ (.A0(\mem_rdata_q[27] ),
    .A1(net2875),
    .S(net736),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _11535_ (.A0(\mem_rdata_q[28] ),
    .A1(net2729),
    .S(net736),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _11536_ (.A0(\mem_rdata_q[29] ),
    .A1(net2643),
    .S(net736),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _11537_ (.A0(\mem_rdata_q[30] ),
    .A1(net194),
    .S(net736),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _11538_ (.A0(\mem_rdata_q[31] ),
    .A1(net2588),
    .S(net736),
    .X(_00853_));
 sky130_fd_sc_hd__nand2_1 _11539_ (.A(net1),
    .B(net12),
    .Y(_06165_));
 sky130_fd_sc_hd__or3b_1 _11540_ (.A(_06165_),
    .B(net26),
    .C_N(net23),
    .X(_06166_));
 sky130_fd_sc_hd__inv_2 _11541_ (.A(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__and4b_1 _11542_ (.A_N(net29),
    .B(net27),
    .C(net28),
    .D(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__mux2_1 _11543_ (.A0(net2557),
    .A1(_06168_),
    .S(net547),
    .X(_00854_));
 sky130_fd_sc_hd__or3b_1 _11544_ (.A(net29),
    .B(net28),
    .C_N(net27),
    .X(_06169_));
 sky130_fd_sc_hd__nor2_1 _11545_ (.A(_06166_),
    .B(_06169_),
    .Y(_06170_));
 sky130_fd_sc_hd__mux2_1 _11546_ (.A0(net1414),
    .A1(_06170_),
    .S(net547),
    .X(_00855_));
 sky130_fd_sc_hd__nand3b_1 _11547_ (.A_N(net27),
    .B(net28),
    .C(net29),
    .Y(_06171_));
 sky130_fd_sc_hd__nand2_1 _11548_ (.A(net26),
    .B(net23),
    .Y(_06172_));
 sky130_fd_sc_hd__o31a_1 _11549_ (.A1(_06165_),
    .A2(_06171_),
    .A3(_06172_),
    .B1(net547),
    .X(_06173_));
 sky130_fd_sc_hd__o21ba_1 _11550_ (.A1(net1152),
    .A2(net547),
    .B1_N(_06173_),
    .X(_00856_));
 sky130_fd_sc_hd__nor2_1 _11551_ (.A(net1209),
    .B(net746),
    .Y(_06174_));
 sky130_fd_sc_hd__nor3_2 _11552_ (.A(\mem_rdata_q[14] ),
    .B(\mem_rdata_q[13] ),
    .C(\mem_rdata_q[12] ),
    .Y(_06175_));
 sky130_fd_sc_hd__and2_1 _11553_ (.A(net746),
    .B(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__inv_2 _11554_ (.A(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__and3_2 _11555_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(net1233),
    .C(net747),
    .X(_06178_));
 sky130_fd_sc_hd__a22o_1 _11556_ (.A1(net1998),
    .A2(net563),
    .B1(_06175_),
    .B2(_06178_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2b_1 _11557_ (.A_N(\mem_rdata_q[13] ),
    .B(\mem_rdata_q[12] ),
    .Y(_06179_));
 sky130_fd_sc_hd__nor2_1 _11558_ (.A(\mem_rdata_q[14] ),
    .B(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__and2_1 _11559_ (.A(net747),
    .B(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__a22o_1 _11560_ (.A1(net3018),
    .A2(net561),
    .B1(_06178_),
    .B2(_06180_),
    .X(_00858_));
 sky130_fd_sc_hd__nor3_1 _11561_ (.A(_02388_),
    .B(\mem_rdata_q[13] ),
    .C(\mem_rdata_q[12] ),
    .Y(_06182_));
 sky130_fd_sc_hd__a22o_1 _11562_ (.A1(net2609),
    .A2(net561),
    .B1(_06178_),
    .B2(_06182_),
    .X(_00859_));
 sky130_fd_sc_hd__nor2_2 _11563_ (.A(_02388_),
    .B(_06179_),
    .Y(_06183_));
 sky130_fd_sc_hd__a22o_1 _11564_ (.A1(net2778),
    .A2(net561),
    .B1(_06178_),
    .B2(_06183_),
    .X(_00860_));
 sky130_fd_sc_hd__and3b_1 _11565_ (.A_N(\mem_rdata_q[12] ),
    .B(\mem_rdata_q[13] ),
    .C(\mem_rdata_q[14] ),
    .X(_06184_));
 sky130_fd_sc_hd__a22o_1 _11566_ (.A1(net1649),
    .A2(net562),
    .B1(_06178_),
    .B2(_06184_),
    .X(_00861_));
 sky130_fd_sc_hd__and3_1 _11567_ (.A(\mem_rdata_q[14] ),
    .B(\mem_rdata_q[13] ),
    .C(\mem_rdata_q[12] ),
    .X(_06185_));
 sky130_fd_sc_hd__a22o_1 _11568_ (.A1(net2994),
    .A2(net563),
    .B1(_06178_),
    .B2(_06185_),
    .X(_00862_));
 sky130_fd_sc_hd__or4_1 _11569_ (.A(net5),
    .B(net4),
    .C(_06166_),
    .D(_06171_),
    .X(_06186_));
 sky130_fd_sc_hd__or4_1 _11570_ (.A(_02369_),
    .B(net6),
    .C(_02452_),
    .D(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__o21ai_1 _11571_ (.A1(_02382_),
    .A2(net547),
    .B1(_06187_),
    .Y(_00863_));
 sky130_fd_sc_hd__a22o_1 _11572_ (.A1(net3036),
    .A2(net740),
    .B1(_06176_),
    .B2(is_lb_lh_lw_lbu_lhu),
    .X(_00864_));
 sky130_fd_sc_hd__a22o_1 _11573_ (.A1(instr_lh),
    .A2(net741),
    .B1(_06181_),
    .B2(is_lb_lh_lw_lbu_lhu),
    .X(_00865_));
 sky130_fd_sc_hd__or3b_2 _11574_ (.A(\mem_rdata_q[14] ),
    .B(\mem_rdata_q[12] ),
    .C_N(\mem_rdata_q[13] ),
    .X(_06188_));
 sky130_fd_sc_hd__inv_2 _11575_ (.A(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nor2_1 _11576_ (.A(net741),
    .B(_06188_),
    .Y(_06190_));
 sky130_fd_sc_hd__a22o_1 _11577_ (.A1(net2904),
    .A2(net740),
    .B1(_06190_),
    .B2(is_lb_lh_lw_lbu_lhu),
    .X(_00866_));
 sky130_fd_sc_hd__and2_1 _11578_ (.A(is_lb_lh_lw_lbu_lhu),
    .B(net747),
    .X(_06191_));
 sky130_fd_sc_hd__a22o_1 _11579_ (.A1(net2930),
    .A2(net740),
    .B1(net732),
    .B2(_06191_),
    .X(_00867_));
 sky130_fd_sc_hd__a22o_1 _11580_ (.A1(net2849),
    .A2(net740),
    .B1(_06183_),
    .B2(_06191_),
    .X(_00868_));
 sky130_fd_sc_hd__a22o_1 _11581_ (.A1(net2912),
    .A2(net740),
    .B1(_06176_),
    .B2(is_sb_sh_sw),
    .X(_00869_));
 sky130_fd_sc_hd__a22o_1 _11582_ (.A1(net2932),
    .A2(net741),
    .B1(_06181_),
    .B2(is_sb_sh_sw),
    .X(_00870_));
 sky130_fd_sc_hd__and3_2 _11583_ (.A(net1234),
    .B(is_alu_reg_imm),
    .C(net746),
    .X(_06192_));
 sky130_fd_sc_hd__a22o_1 _11584_ (.A1(net2281),
    .A2(net563),
    .B1(_06175_),
    .B2(_06192_),
    .X(_00871_));
 sky130_fd_sc_hd__a22o_1 _11585_ (.A1(net2802),
    .A2(net562),
    .B1(_06189_),
    .B2(_06192_),
    .X(_00872_));
 sky130_fd_sc_hd__and3_1 _11586_ (.A(_02388_),
    .B(\mem_rdata_q[13] ),
    .C(\mem_rdata_q[12] ),
    .X(_06193_));
 sky130_fd_sc_hd__a22o_1 _11587_ (.A1(net2550),
    .A2(net561),
    .B1(_06192_),
    .B2(_06193_),
    .X(_00873_));
 sky130_fd_sc_hd__a22o_1 _11588_ (.A1(net3024),
    .A2(net561),
    .B1(net732),
    .B2(_06192_),
    .X(_00874_));
 sky130_fd_sc_hd__a22o_1 _11589_ (.A1(net2864),
    .A2(net562),
    .B1(_06184_),
    .B2(_06192_),
    .X(_00875_));
 sky130_fd_sc_hd__a22o_1 _11590_ (.A1(net2922),
    .A2(net563),
    .B1(_06185_),
    .B2(_06192_),
    .X(_00876_));
 sky130_fd_sc_hd__a22o_1 _11591_ (.A1(net2896),
    .A2(net740),
    .B1(_06190_),
    .B2(is_sb_sh_sw),
    .X(_00877_));
 sky130_fd_sc_hd__nor2_1 _11592_ (.A(\mem_rdata_q[29] ),
    .B(\mem_rdata_q[28] ),
    .Y(_06194_));
 sky130_fd_sc_hd__or4_1 _11593_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[27] ),
    .C(\mem_rdata_q[26] ),
    .D(\mem_rdata_q[25] ),
    .X(_06195_));
 sky130_fd_sc_hd__or3_2 _11594_ (.A(\mem_rdata_q[31] ),
    .B(\mem_rdata_q[29] ),
    .C(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__nor2_1 _11595_ (.A(\mem_rdata_q[30] ),
    .B(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__or2_1 _11596_ (.A(\mem_rdata_q[30] ),
    .B(_06196_),
    .X(_06198_));
 sky130_fd_sc_hd__a32o_1 _11597_ (.A1(is_alu_reg_imm),
    .A2(_06181_),
    .A3(_06197_),
    .B1(net740),
    .B2(net2362),
    .X(_00878_));
 sky130_fd_sc_hd__nor2_1 _11598_ (.A(net741),
    .B(_06196_),
    .Y(_06199_));
 sky130_fd_sc_hd__nor2_1 _11599_ (.A(net741),
    .B(_06198_),
    .Y(_06200_));
 sky130_fd_sc_hd__a32o_1 _11600_ (.A1(is_alu_reg_imm),
    .A2(_06183_),
    .A3(_06200_),
    .B1(net741),
    .B2(instr_srli),
    .X(_00879_));
 sky130_fd_sc_hd__and3_2 _11601_ (.A(net1234),
    .B(is_alu_reg_reg),
    .C(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__a22o_1 _11602_ (.A1(net2400),
    .A2(net563),
    .B1(_06175_),
    .B2(_06201_),
    .X(_00880_));
 sky130_fd_sc_hd__and4_1 _11603_ (.A(net1234),
    .B(\mem_rdata_q[30] ),
    .C(is_alu_reg_reg),
    .D(_06199_),
    .X(_06202_));
 sky130_fd_sc_hd__a22o_1 _11604_ (.A1(net1145),
    .A2(net563),
    .B1(_06175_),
    .B2(_06202_),
    .X(_00881_));
 sky130_fd_sc_hd__a22o_1 _11605_ (.A1(net2800),
    .A2(net561),
    .B1(_06180_),
    .B2(_06201_),
    .X(_00882_));
 sky130_fd_sc_hd__a22o_1 _11606_ (.A1(net2654),
    .A2(net562),
    .B1(_06189_),
    .B2(_06201_),
    .X(_00883_));
 sky130_fd_sc_hd__a22o_1 _11607_ (.A1(net2572),
    .A2(net561),
    .B1(_06193_),
    .B2(_06201_),
    .X(_00884_));
 sky130_fd_sc_hd__a22o_1 _11608_ (.A1(net3032),
    .A2(net561),
    .B1(net732),
    .B2(_06201_),
    .X(_00885_));
 sky130_fd_sc_hd__a22o_1 _11609_ (.A1(instr_srl),
    .A2(net561),
    .B1(_06183_),
    .B2(_06201_),
    .X(_00886_));
 sky130_fd_sc_hd__a22o_1 _11610_ (.A1(net2608),
    .A2(net563),
    .B1(_06183_),
    .B2(_06202_),
    .X(_00887_));
 sky130_fd_sc_hd__a22o_1 _11611_ (.A1(net2727),
    .A2(net562),
    .B1(_06184_),
    .B2(_06201_),
    .X(_00888_));
 sky130_fd_sc_hd__a22o_1 _11612_ (.A1(net3005),
    .A2(net563),
    .B1(_06185_),
    .B2(_06201_),
    .X(_00889_));
 sky130_fd_sc_hd__and4_1 _11613_ (.A(is_alu_reg_imm),
    .B(\mem_rdata_q[30] ),
    .C(_06183_),
    .D(_06199_),
    .X(_06203_));
 sky130_fd_sc_hd__a21o_1 _11614_ (.A1(net1862),
    .A2(net741),
    .B1(_06203_),
    .X(_00890_));
 sky130_fd_sc_hd__and4_1 _11615_ (.A(\mem_rdata_q[31] ),
    .B(\mem_rdata_q[30] ),
    .C(net746),
    .D(_06194_),
    .X(_06204_));
 sky130_fd_sc_hd__nor2_1 _11616_ (.A(\mem_rdata_q[25] ),
    .B(\mem_rdata_q[24] ),
    .Y(_06205_));
 sky130_fd_sc_hd__and4bb_1 _11617_ (.A_N(\mem_rdata_q[27] ),
    .B_N(\mem_rdata_q[26] ),
    .C(_06204_),
    .D(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__or3_1 _11618_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .C(\mem_rdata_q[21] ),
    .X(_06207_));
 sky130_fd_sc_hd__nand2_1 _11619_ (.A(\mem_rdata_q[4] ),
    .B(\mem_rdata_q[6] ),
    .Y(_06208_));
 sky130_fd_sc_hd__or4_1 _11620_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .D(\mem_rdata_q[2] ),
    .X(_06209_));
 sky130_fd_sc_hd__nand2_1 _11621_ (.A(\mem_rdata_q[0] ),
    .B(\mem_rdata_q[1] ),
    .Y(_06210_));
 sky130_fd_sc_hd__or4_1 _11622_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .C(_06209_),
    .D(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__or4_1 _11623_ (.A(\mem_rdata_q[3] ),
    .B(_02401_),
    .C(_06208_),
    .D(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__or2_1 _11624_ (.A(_06188_),
    .B(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__nor2_1 _11625_ (.A(_06207_),
    .B(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__a22o_1 _11626_ (.A1(net3057),
    .A2(net737),
    .B1(_06206_),
    .B2(_06214_),
    .X(_00891_));
 sky130_fd_sc_hd__and4b_1 _11627_ (.A_N(\mem_rdata_q[26] ),
    .B(_06204_),
    .C(_06205_),
    .D(\mem_rdata_q[27] ),
    .X(_06215_));
 sky130_fd_sc_hd__a22o_1 _11628_ (.A1(instr_rdcycleh),
    .A2(net738),
    .B1(_06214_),
    .B2(_06215_),
    .X(_00892_));
 sky130_fd_sc_hd__or4b_1 _11629_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .C(\mem_rdata_q[20] ),
    .D_N(\mem_rdata_q[21] ),
    .X(_06216_));
 sky130_fd_sc_hd__nor2_1 _11630_ (.A(_06213_),
    .B(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__a22o_1 _11631_ (.A1(net3029),
    .A2(net737),
    .B1(_06206_),
    .B2(_06217_),
    .X(_00893_));
 sky130_fd_sc_hd__a22o_1 _11632_ (.A1(net1134),
    .A2(net737),
    .B1(_06215_),
    .B2(_06217_),
    .X(_00894_));
 sky130_fd_sc_hd__or4b_1 _11633_ (.A(\mem_rdata_q[4] ),
    .B(\mem_rdata_q[5] ),
    .C(\mem_rdata_q[6] ),
    .D_N(\mem_rdata_q[3] ),
    .X(_06218_));
 sky130_fd_sc_hd__nor4_1 _11634_ (.A(net1208),
    .B(_02400_),
    .C(_06210_),
    .D(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__a22o_1 _11635_ (.A1(net2398),
    .A2(_06174_),
    .B1(_06176_),
    .B2(net731),
    .X(_00895_));
 sky130_fd_sc_hd__or4_1 _11636_ (.A(\mem_rdata_q[11] ),
    .B(\mem_rdata_q[10] ),
    .C(\mem_rdata_q[9] ),
    .D(\mem_rdata_q[8] ),
    .X(_06220_));
 sky130_fd_sc_hd__or4_1 _11637_ (.A(\mem_rdata_q[24] ),
    .B(\mem_rdata_q[7] ),
    .C(_06207_),
    .D(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__or4_1 _11638_ (.A(_06177_),
    .B(_06198_),
    .C(_06212_),
    .D(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__a21bo_1 _11639_ (.A1(net1353),
    .A2(net741),
    .B1_N(_06222_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _11640_ (.A0(\decoded_imm_j[4] ),
    .A1(net17),
    .S(net546),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(net3064),
    .A1(net18),
    .S(net545),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _11642_ (.A0(\decoded_imm_j[6] ),
    .A1(net19),
    .S(net545),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _11643_ (.A0(\decoded_imm_j[7] ),
    .A1(net20),
    .S(net545),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _11644_ (.A0(net2984),
    .A1(net21),
    .S(net545),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _11645_ (.A0(\decoded_imm_j[9] ),
    .A1(net22),
    .S(net545),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(\decoded_imm_j[10] ),
    .A1(net24),
    .S(net545),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(\decoded_imm_j[12] ),
    .A1(net4),
    .S(net545),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _11648_ (.A0(\decoded_imm_j[13] ),
    .A1(net5),
    .S(net545),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _11649_ (.A0(\decoded_imm_j[14] ),
    .A1(net6),
    .S(net545),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _11650_ (.A0(net3044),
    .A1(net11),
    .S(net546),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _11651_ (.A0(\decoded_imm_j[20] ),
    .A1(net25),
    .S(net547),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _11652_ (.A0(net1740),
    .A1(net30),
    .S(net548),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _11653_ (.A0(net1465),
    .A1(net31),
    .S(net548),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(net1406),
    .A1(net32),
    .S(net548),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _11655_ (.A0(net1613),
    .A1(net2),
    .S(net548),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _11656_ (.A0(net1405),
    .A1(net3),
    .S(net548),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _11657_ (.A0(\decoded_imm_j[15] ),
    .A1(net7),
    .S(net546),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _11658_ (.A0(\decoded_imm_j[16] ),
    .A1(net8),
    .S(net546),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _11659_ (.A0(\decoded_imm_j[17] ),
    .A1(net9),
    .S(net546),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(\decoded_imm_j[18] ),
    .A1(net10),
    .S(net546),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(\decoded_imm_j[11] ),
    .A1(net13),
    .S(net545),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(\decoded_imm_j[1] ),
    .A1(net14),
    .S(net546),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _11663_ (.A0(\decoded_imm_j[2] ),
    .A1(net15),
    .S(net546),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(\decoded_imm_j[3] ),
    .A1(net16),
    .S(net546),
    .X(_00921_));
 sky130_fd_sc_hd__or3_2 _11665_ (.A(instr_jalr),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(is_alu_reg_imm),
    .X(_06223_));
 sky130_fd_sc_hd__and3_1 _11666_ (.A(\mem_rdata_q[20] ),
    .B(net745),
    .C(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__and3_1 _11667_ (.A(is_sb_sh_sw),
    .B(\mem_rdata_q[7] ),
    .C(net745),
    .X(_06225_));
 sky130_fd_sc_hd__a211o_1 _11668_ (.A1(\decoded_imm[0] ),
    .A2(net734),
    .B1(_06224_),
    .C1(_06225_),
    .X(_00922_));
 sky130_fd_sc_hd__or3_2 _11669_ (.A(net26),
    .B(net23),
    .C(_06165_),
    .X(_06226_));
 sky130_fd_sc_hd__inv_2 _11670_ (.A(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__nor4_1 _11671_ (.A(net29),
    .B(net27),
    .C(net28),
    .D(_06226_),
    .Y(_06228_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(is_lb_lh_lw_lbu_lhu),
    .A1(_06228_),
    .S(net547),
    .X(_00923_));
 sky130_fd_sc_hd__a2111oi_1 _11673_ (.A1(\mem_rdata_q[30] ),
    .A2(_02388_),
    .B1(net737),
    .C1(_06179_),
    .D1(_06196_),
    .Y(_06229_));
 sky130_fd_sc_hd__a22o_1 _11674_ (.A1(net2671),
    .A2(net737),
    .B1(_06229_),
    .B2(is_alu_reg_imm),
    .X(_00924_));
 sky130_fd_sc_hd__a211o_1 _11675_ (.A1(is_alu_reg_imm),
    .A2(_06179_),
    .B1(net737),
    .C1(instr_jalr),
    .X(_06230_));
 sky130_fd_sc_hd__o21a_1 _11676_ (.A1(net2658),
    .A2(net747),
    .B1(_06230_),
    .X(_00925_));
 sky130_fd_sc_hd__or4b_1 _11677_ (.A(net29),
    .B(_06226_),
    .C(net27),
    .D_N(net28),
    .X(_06231_));
 sky130_fd_sc_hd__inv_2 _11678_ (.A(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__mux2_1 _11679_ (.A0(is_sb_sh_sw),
    .A1(_06232_),
    .S(net548),
    .X(_00926_));
 sky130_fd_sc_hd__a22o_1 _11680_ (.A1(net2688),
    .A2(net737),
    .B1(net560),
    .B2(net2710),
    .X(_00927_));
 sky130_fd_sc_hd__o21ai_1 _11681_ (.A1(_06171_),
    .A2(_06226_),
    .B1(net547),
    .Y(_06233_));
 sky130_fd_sc_hd__o211a_1 _11682_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(net548),
    .B1(_06233_),
    .C1(net1233),
    .X(_00928_));
 sky130_fd_sc_hd__and3_1 _11683_ (.A(\latched_rd[1] ),
    .B(\latched_rd[0] ),
    .C(_04290_),
    .X(_06234_));
 sky130_fd_sc_hd__mux2_1 _11684_ (.A0(net1937),
    .A1(net586),
    .S(net375),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(net2079),
    .A1(net584),
    .S(net375),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _11686_ (.A0(net1696),
    .A1(net582),
    .S(net375),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _11687_ (.A0(net1853),
    .A1(net578),
    .S(net374),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _11688_ (.A0(net2193),
    .A1(net573),
    .S(net374),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _11689_ (.A0(net1854),
    .A1(net542),
    .S(net374),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _11690_ (.A0(net1982),
    .A1(net540),
    .S(net374),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _11691_ (.A0(net1796),
    .A1(net524),
    .S(net373),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(net1858),
    .A1(net522),
    .S(net373),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _11693_ (.A0(net1859),
    .A1(net409),
    .S(net373),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(net1747),
    .A1(net406),
    .S(net373),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _11695_ (.A0(net2033),
    .A1(net355),
    .S(net373),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(net2029),
    .A1(net351),
    .S(net373),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _11697_ (.A0(net1978),
    .A1(net348),
    .S(net373),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(net1663),
    .A1(net345),
    .S(net374),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _11699_ (.A0(net1769),
    .A1(net340),
    .S(net373),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(net1991),
    .A1(net337),
    .S(net374),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _11701_ (.A0(net1988),
    .A1(net332),
    .S(net373),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(net1909),
    .A1(net330),
    .S(net373),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _11703_ (.A0(net2149),
    .A1(net326),
    .S(net375),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(net1888),
    .A1(net322),
    .S(net374),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _11705_ (.A0(net1906),
    .A1(net319),
    .S(net374),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(net2052),
    .A1(net314),
    .S(net375),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(net2066),
    .A1(net310),
    .S(net375),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(net1925),
    .A1(net307),
    .S(net375),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _11709_ (.A0(net2442),
    .A1(net304),
    .S(net375),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _11710_ (.A0(net2011),
    .A1(net300),
    .S(net375),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(net1968),
    .A1(net295),
    .S(net376),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _11712_ (.A0(net2040),
    .A1(net292),
    .S(net376),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _11713_ (.A0(net2163),
    .A1(net288),
    .S(net375),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(net2096),
    .A1(net282),
    .S(net376),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _11715_ (.A0(net2118),
    .A1(net280),
    .S(net376),
    .X(_00960_));
 sky130_fd_sc_hd__nor2_1 _11716_ (.A(_06169_),
    .B(_06226_),
    .Y(_06235_));
 sky130_fd_sc_hd__mux2_1 _11717_ (.A0(is_alu_reg_imm),
    .A1(_06235_),
    .S(net547),
    .X(_00961_));
 sky130_fd_sc_hd__and4b_1 _11718_ (.A_N(net29),
    .B(net27),
    .C(net28),
    .D(_06227_),
    .X(_06236_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(net2710),
    .A1(_06236_),
    .S(net547),
    .X(_00962_));
 sky130_fd_sc_hd__or4_1 _11720_ (.A(instr_sltu),
    .B(instr_slt),
    .C(instr_sltiu),
    .D(instr_slti),
    .X(_06237_));
 sky130_fd_sc_hd__o21a_1 _11721_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(_06237_),
    .B1(net561),
    .X(_00963_));
 sky130_fd_sc_hd__nor2_1 _11722_ (.A(net1208),
    .B(net268),
    .Y(_06238_));
 sky130_fd_sc_hd__or2_1 _11723_ (.A(net1209),
    .B(net268),
    .X(_06239_));
 sky130_fd_sc_hd__o21a_4 _11724_ (.A1(net96),
    .A2(net129),
    .B1(_06238_),
    .X(_06240_));
 sky130_fd_sc_hd__and2b_1 _11725_ (.A_N(mem_do_wdata),
    .B(net982),
    .X(_06241_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(net1834),
    .A1(_06241_),
    .S(net536),
    .X(_00964_));
 sky130_fd_sc_hd__or3_2 _11727_ (.A(net1208),
    .B(_02487_),
    .C(_06149_),
    .X(_06242_));
 sky130_fd_sc_hd__and3_2 _11728_ (.A(_02363_),
    .B(net1089),
    .C(net1232),
    .X(_06243_));
 sky130_fd_sc_hd__a22o_1 _11729_ (.A1(\latched_rd[0] ),
    .A2(_06242_),
    .B1(_06243_),
    .B2(net1740),
    .X(_00965_));
 sky130_fd_sc_hd__a22o_1 _11730_ (.A1(\latched_rd[1] ),
    .A2(_06242_),
    .B1(_06243_),
    .B2(net1465),
    .X(_00966_));
 sky130_fd_sc_hd__a22o_1 _11731_ (.A1(\latched_rd[2] ),
    .A2(_06242_),
    .B1(_06243_),
    .B2(net1406),
    .X(_00967_));
 sky130_fd_sc_hd__a22o_1 _11732_ (.A1(\latched_rd[3] ),
    .A2(_06242_),
    .B1(_06243_),
    .B2(net1613),
    .X(_00968_));
 sky130_fd_sc_hd__a22o_1 _11733_ (.A1(\latched_rd[4] ),
    .A2(_06242_),
    .B1(_06243_),
    .B2(net1405),
    .X(_00969_));
 sky130_fd_sc_hd__and3_2 _11734_ (.A(mem_do_wdata),
    .B(_02418_),
    .C(_06238_),
    .X(_06244_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(net1426),
    .A1(net1181),
    .S(net727),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(net1468),
    .A1(net1179),
    .S(net729),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _11737_ (.A0(net1736),
    .A1(net119),
    .S(net727),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _11738_ (.A0(net1876),
    .A1(net122),
    .S(net727),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _11739_ (.A0(net1735),
    .A1(net1175),
    .S(net729),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(net1575),
    .A1(net1173),
    .S(net729),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _11741_ (.A0(net1462),
    .A1(net1171),
    .S(net729),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(net1700),
    .A1(net1170),
    .S(net729),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _11743_ (.A0(net1495),
    .A1(net127),
    .S(net730),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _11744_ (.A0(net1635),
    .A1(net128),
    .S(net730),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _11745_ (.A0(net1447),
    .A1(net98),
    .S(net727),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(net1642),
    .A1(net99),
    .S(net730),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _11747_ (.A0(net1965),
    .A1(net100),
    .S(net730),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(net1482),
    .A1(net101),
    .S(net727),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _11749_ (.A0(net1890),
    .A1(net102),
    .S(net727),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(net1508),
    .A1(net103),
    .S(net728),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _11751_ (.A0(net1718),
    .A1(net104),
    .S(net727),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _11752_ (.A0(net2647),
    .A1(net105),
    .S(net730),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(net1512),
    .A1(net106),
    .S(net730),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(net1398),
    .A1(net107),
    .S(net727),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(net1546),
    .A1(net109),
    .S(net727),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _11756_ (.A0(net1437),
    .A1(net110),
    .S(net727),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(net1644),
    .A1(net111),
    .S(net730),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _11758_ (.A0(net1520),
    .A1(net112),
    .S(net728),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _11759_ (.A0(net2548),
    .A1(net113),
    .S(net729),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(net1669),
    .A1(net114),
    .S(net729),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _11761_ (.A0(net1807),
    .A1(net115),
    .S(net729),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(net2698),
    .A1(net116),
    .S(net729),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _11763_ (.A0(net1761),
    .A1(net117),
    .S(net730),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(net1673),
    .A1(net118),
    .S(net729),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _11765_ (.A0(net1791),
    .A1(net120),
    .S(net728),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(net1479),
    .A1(net121),
    .S(net728),
    .X(_01001_));
 sky130_fd_sc_hd__nand2b_4 _11767_ (.A_N(net268),
    .B(net96),
    .Y(_06245_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(net167),
    .A1(net130),
    .S(net536),
    .X(_06246_));
 sky130_fd_sc_hd__and2_1 _11769_ (.A(_06245_),
    .B(_06246_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(net168),
    .A1(net131),
    .S(net536),
    .X(_06247_));
 sky130_fd_sc_hd__and2_1 _11771_ (.A(_06245_),
    .B(_06247_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(net169),
    .A1(net132),
    .S(net536),
    .X(_06248_));
 sky130_fd_sc_hd__and2_1 _11773_ (.A(_06245_),
    .B(_06248_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _11774_ (.A0(net170),
    .A1(net133),
    .S(net536),
    .X(_06249_));
 sky130_fd_sc_hd__and2_1 _11775_ (.A(_06245_),
    .B(_06249_),
    .X(_01005_));
 sky130_fd_sc_hd__or2_1 _11776_ (.A(mem_do_wdata),
    .B(_02419_),
    .X(_06250_));
 sky130_fd_sc_hd__or4_1 _11777_ (.A(_02418_),
    .B(_02448_),
    .C(net964),
    .D(_06239_),
    .X(_06251_));
 sky130_fd_sc_hd__o31ai_1 _11778_ (.A1(_02417_),
    .A2(_06239_),
    .A3(_06250_),
    .B1(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__and3b_1 _11779_ (.A_N(net33),
    .B(net268),
    .C(net1234),
    .X(_06253_));
 sky130_fd_sc_hd__a211o_1 _11780_ (.A1(_02448_),
    .A2(_06238_),
    .B1(_06252_),
    .C1(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__a21o_1 _11781_ (.A1(net2817),
    .A2(_06254_),
    .B1(net536),
    .X(_01006_));
 sky130_fd_sc_hd__nor2_1 _11782_ (.A(net175),
    .B(net174),
    .Y(_06255_));
 sky130_fd_sc_hd__and2_1 _11783_ (.A(_04299_),
    .B(_06255_),
    .X(_01007_));
 sky130_fd_sc_hd__o311a_1 _11784_ (.A1(net1157),
    .A2(net258),
    .A3(_05118_),
    .B1(_03368_),
    .C1(\genblk2.pcpi_div.instr_div ),
    .X(_06256_));
 sky130_fd_sc_hd__a211o_1 _11785_ (.A1(net1189),
    .A2(\genblk2.pcpi_div.instr_rem ),
    .B1(net866),
    .C1(net1216),
    .X(_06257_));
 sky130_fd_sc_hd__o22a_1 _11786_ (.A1(\genblk2.pcpi_div.outsign ),
    .A2(_05120_),
    .B1(_06256_),
    .B2(_06257_),
    .X(_01008_));
 sky130_fd_sc_hd__nor2_1 _11787_ (.A(net867),
    .B(_05095_),
    .Y(_06258_));
 sky130_fd_sc_hd__and2b_1 _11788_ (.A_N(\genblk2.pcpi_div.divisor[31] ),
    .B(\genblk2.pcpi_div.dividend[31] ),
    .X(_06259_));
 sky130_fd_sc_hd__xor2_1 _11789_ (.A(\genblk2.pcpi_div.divisor[30] ),
    .B(\genblk2.pcpi_div.dividend[30] ),
    .X(_06260_));
 sky130_fd_sc_hd__nand2b_1 _11790_ (.A_N(\genblk2.pcpi_div.dividend[29] ),
    .B(\genblk2.pcpi_div.divisor[29] ),
    .Y(_06261_));
 sky130_fd_sc_hd__inv_2 _11791_ (.A(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__nand2b_1 _11792_ (.A_N(\genblk2.pcpi_div.divisor[29] ),
    .B(\genblk2.pcpi_div.dividend[29] ),
    .Y(_06263_));
 sky130_fd_sc_hd__and2b_1 _11793_ (.A_N(\genblk2.pcpi_div.divisor[28] ),
    .B(\genblk2.pcpi_div.dividend[28] ),
    .X(_06264_));
 sky130_fd_sc_hd__and2b_1 _11794_ (.A_N(\genblk2.pcpi_div.dividend[28] ),
    .B(\genblk2.pcpi_div.divisor[28] ),
    .X(_06265_));
 sky130_fd_sc_hd__or2_1 _11795_ (.A(_06264_),
    .B(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__and2b_1 _11796_ (.A_N(\genblk2.pcpi_div.divisor[24] ),
    .B(\genblk2.pcpi_div.dividend[24] ),
    .X(_06267_));
 sky130_fd_sc_hd__and2b_1 _11797_ (.A_N(\genblk2.pcpi_div.dividend[24] ),
    .B(\genblk2.pcpi_div.divisor[24] ),
    .X(_06268_));
 sky130_fd_sc_hd__nor2_1 _11798_ (.A(_06267_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__and2b_1 _11799_ (.A_N(\genblk2.pcpi_div.divisor[23] ),
    .B(\genblk2.pcpi_div.dividend[23] ),
    .X(_06270_));
 sky130_fd_sc_hd__and2b_1 _11800_ (.A_N(\genblk2.pcpi_div.dividend[23] ),
    .B(\genblk2.pcpi_div.divisor[23] ),
    .X(_06271_));
 sky130_fd_sc_hd__nand2b_1 _11801_ (.A_N(\genblk2.pcpi_div.divisor[22] ),
    .B(\genblk2.pcpi_div.dividend[22] ),
    .Y(_06272_));
 sky130_fd_sc_hd__xnor2_1 _11802_ (.A(\genblk2.pcpi_div.divisor[22] ),
    .B(\genblk2.pcpi_div.dividend[22] ),
    .Y(_06273_));
 sky130_fd_sc_hd__or3b_1 _11803_ (.A(_06270_),
    .B(_06271_),
    .C_N(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__and2b_1 _11804_ (.A_N(\genblk2.pcpi_div.divisor[21] ),
    .B(\genblk2.pcpi_div.dividend[21] ),
    .X(_06275_));
 sky130_fd_sc_hd__and2b_1 _11805_ (.A_N(\genblk2.pcpi_div.dividend[21] ),
    .B(\genblk2.pcpi_div.divisor[21] ),
    .X(_06276_));
 sky130_fd_sc_hd__or2_1 _11806_ (.A(_06275_),
    .B(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__xnor2_1 _11807_ (.A(\genblk2.pcpi_div.divisor[20] ),
    .B(\genblk2.pcpi_div.dividend[20] ),
    .Y(_06278_));
 sky130_fd_sc_hd__and2b_1 _11808_ (.A_N(\genblk2.pcpi_div.dividend[19] ),
    .B(\genblk2.pcpi_div.divisor[19] ),
    .X(_06279_));
 sky130_fd_sc_hd__nand2b_1 _11809_ (.A_N(\genblk2.pcpi_div.divisor[18] ),
    .B(\genblk2.pcpi_div.dividend[18] ),
    .Y(_06280_));
 sky130_fd_sc_hd__and2b_1 _11810_ (.A_N(\genblk2.pcpi_div.divisor[19] ),
    .B(\genblk2.pcpi_div.dividend[19] ),
    .X(_06281_));
 sky130_fd_sc_hd__o21ba_1 _11811_ (.A1(_06279_),
    .A2(_06280_),
    .B1_N(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__or2_1 _11812_ (.A(_06279_),
    .B(_06281_),
    .X(_06283_));
 sky130_fd_sc_hd__nand2b_1 _11813_ (.A_N(\genblk2.pcpi_div.dividend[18] ),
    .B(\genblk2.pcpi_div.divisor[18] ),
    .Y(_06284_));
 sky130_fd_sc_hd__nand2_1 _11814_ (.A(_06280_),
    .B(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__nor2_1 _11815_ (.A(_06283_),
    .B(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__and2b_1 _11816_ (.A_N(\genblk2.pcpi_div.dividend[17] ),
    .B(\genblk2.pcpi_div.divisor[17] ),
    .X(_06287_));
 sky130_fd_sc_hd__and2b_1 _11817_ (.A_N(\genblk2.pcpi_div.divisor[17] ),
    .B(\genblk2.pcpi_div.dividend[17] ),
    .X(_06288_));
 sky130_fd_sc_hd__a21oi_1 _11818_ (.A1(_02360_),
    .A2(\genblk2.pcpi_div.dividend[16] ),
    .B1(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__nor2_1 _11819_ (.A(_06287_),
    .B(_06288_),
    .Y(_06290_));
 sky130_fd_sc_hd__xor2_1 _11820_ (.A(\genblk2.pcpi_div.divisor[16] ),
    .B(\genblk2.pcpi_div.dividend[16] ),
    .X(_06291_));
 sky130_fd_sc_hd__and2b_1 _11821_ (.A_N(\genblk2.pcpi_div.dividend[15] ),
    .B(\genblk2.pcpi_div.divisor[15] ),
    .X(_06292_));
 sky130_fd_sc_hd__nand2b_1 _11822_ (.A_N(\genblk2.pcpi_div.divisor[15] ),
    .B(\genblk2.pcpi_div.dividend[15] ),
    .Y(_06293_));
 sky130_fd_sc_hd__xor2_1 _11823_ (.A(\genblk2.pcpi_div.divisor[14] ),
    .B(\genblk2.pcpi_div.dividend[14] ),
    .X(_06294_));
 sky130_fd_sc_hd__and2b_1 _11824_ (.A_N(\genblk2.pcpi_div.dividend[13] ),
    .B(\genblk2.pcpi_div.divisor[13] ),
    .X(_06295_));
 sky130_fd_sc_hd__nand2b_1 _11825_ (.A_N(\genblk2.pcpi_div.divisor[13] ),
    .B(\genblk2.pcpi_div.dividend[13] ),
    .Y(_06296_));
 sky130_fd_sc_hd__nand2b_1 _11826_ (.A_N(\genblk2.pcpi_div.divisor[12] ),
    .B(\genblk2.pcpi_div.dividend[12] ),
    .Y(_06297_));
 sky130_fd_sc_hd__nand2b_1 _11827_ (.A_N(\genblk2.pcpi_div.dividend[12] ),
    .B(\genblk2.pcpi_div.divisor[12] ),
    .Y(_06298_));
 sky130_fd_sc_hd__nand2_1 _11828_ (.A(_06297_),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__and2b_1 _11829_ (.A_N(\genblk2.pcpi_div.divisor[11] ),
    .B(\genblk2.pcpi_div.dividend[11] ),
    .X(_06300_));
 sky130_fd_sc_hd__nand2b_1 _11830_ (.A_N(\genblk2.pcpi_div.divisor[11] ),
    .B(\genblk2.pcpi_div.dividend[11] ),
    .Y(_06301_));
 sky130_fd_sc_hd__and2b_1 _11831_ (.A_N(\genblk2.pcpi_div.dividend[11] ),
    .B(\genblk2.pcpi_div.divisor[11] ),
    .X(_06302_));
 sky130_fd_sc_hd__nand2b_1 _11832_ (.A_N(\genblk2.pcpi_div.divisor[10] ),
    .B(\genblk2.pcpi_div.dividend[10] ),
    .Y(_06303_));
 sky130_fd_sc_hd__xnor2_1 _11833_ (.A(\genblk2.pcpi_div.divisor[10] ),
    .B(\genblk2.pcpi_div.dividend[10] ),
    .Y(_06304_));
 sky130_fd_sc_hd__and2b_1 _11834_ (.A_N(\genblk2.pcpi_div.dividend[9] ),
    .B(\genblk2.pcpi_div.divisor[9] ),
    .X(_06305_));
 sky130_fd_sc_hd__and2b_1 _11835_ (.A_N(\genblk2.pcpi_div.divisor[9] ),
    .B(\genblk2.pcpi_div.dividend[9] ),
    .X(_06306_));
 sky130_fd_sc_hd__and2b_1 _11836_ (.A_N(\genblk2.pcpi_div.divisor[7] ),
    .B(\genblk2.pcpi_div.dividend[7] ),
    .X(_06307_));
 sky130_fd_sc_hd__xor2_1 _11837_ (.A(\genblk2.pcpi_div.divisor[6] ),
    .B(\genblk2.pcpi_div.dividend[6] ),
    .X(_06308_));
 sky130_fd_sc_hd__and2b_1 _11838_ (.A_N(\genblk2.pcpi_div.divisor[5] ),
    .B(\genblk2.pcpi_div.dividend[5] ),
    .X(_06309_));
 sky130_fd_sc_hd__inv_2 _11839_ (.A(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__and2b_1 _11840_ (.A_N(\genblk2.pcpi_div.dividend[5] ),
    .B(\genblk2.pcpi_div.divisor[5] ),
    .X(_06311_));
 sky130_fd_sc_hd__nand2b_1 _11841_ (.A_N(\genblk2.pcpi_div.divisor[4] ),
    .B(\genblk2.pcpi_div.dividend[4] ),
    .Y(_06312_));
 sky130_fd_sc_hd__nand2b_1 _11842_ (.A_N(\genblk2.pcpi_div.dividend[4] ),
    .B(\genblk2.pcpi_div.divisor[4] ),
    .Y(_06313_));
 sky130_fd_sc_hd__and2b_1 _11843_ (.A_N(\genblk2.pcpi_div.divisor[3] ),
    .B(\genblk2.pcpi_div.dividend[3] ),
    .X(_06314_));
 sky130_fd_sc_hd__nand2b_1 _11844_ (.A_N(\genblk2.pcpi_div.divisor[3] ),
    .B(\genblk2.pcpi_div.dividend[3] ),
    .Y(_06315_));
 sky130_fd_sc_hd__and2b_1 _11845_ (.A_N(\genblk2.pcpi_div.divisor[2] ),
    .B(\genblk2.pcpi_div.dividend[2] ),
    .X(_06316_));
 sky130_fd_sc_hd__nand2b_1 _11846_ (.A_N(\genblk2.pcpi_div.divisor[2] ),
    .B(\genblk2.pcpi_div.dividend[2] ),
    .Y(_06317_));
 sky130_fd_sc_hd__nand2b_1 _11847_ (.A_N(\genblk2.pcpi_div.dividend[2] ),
    .B(\genblk2.pcpi_div.divisor[2] ),
    .Y(_06318_));
 sky130_fd_sc_hd__and2b_1 _11848_ (.A_N(\genblk2.pcpi_div.divisor[1] ),
    .B(\genblk2.pcpi_div.dividend[1] ),
    .X(_06319_));
 sky130_fd_sc_hd__nand2b_1 _11849_ (.A_N(\genblk2.pcpi_div.dividend[0] ),
    .B(\genblk2.pcpi_div.divisor[0] ),
    .Y(_06320_));
 sky130_fd_sc_hd__xnor2_1 _11850_ (.A(\genblk2.pcpi_div.divisor[1] ),
    .B(\genblk2.pcpi_div.dividend[1] ),
    .Y(_06321_));
 sky130_fd_sc_hd__and2_1 _11851_ (.A(_06320_),
    .B(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__o211a_1 _11852_ (.A1(_06319_),
    .A2(_06322_),
    .B1(_06317_),
    .C1(_06318_),
    .X(_06323_));
 sky130_fd_sc_hd__nand2b_1 _11853_ (.A_N(\genblk2.pcpi_div.dividend[3] ),
    .B(\genblk2.pcpi_div.divisor[3] ),
    .Y(_06324_));
 sky130_fd_sc_hd__o211a_1 _11854_ (.A1(_06316_),
    .A2(_06323_),
    .B1(_06324_),
    .C1(_06315_),
    .X(_06325_));
 sky130_fd_sc_hd__o211ai_2 _11855_ (.A1(_06314_),
    .A2(_06325_),
    .B1(_06312_),
    .C1(_06313_),
    .Y(_06326_));
 sky130_fd_sc_hd__and2_1 _11856_ (.A(_06312_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__a311o_1 _11857_ (.A1(_06310_),
    .A2(_06312_),
    .A3(_06326_),
    .B1(_06311_),
    .C1(_06308_),
    .X(_06328_));
 sky130_fd_sc_hd__o21ai_1 _11858_ (.A1(\genblk2.pcpi_div.divisor[6] ),
    .A2(_02391_),
    .B1(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__nand2b_1 _11859_ (.A_N(\genblk2.pcpi_div.dividend[7] ),
    .B(\genblk2.pcpi_div.divisor[7] ),
    .Y(_06330_));
 sky130_fd_sc_hd__nand2b_1 _11860_ (.A_N(_06307_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__a21o_1 _11861_ (.A1(_06329_),
    .A2(_06330_),
    .B1(_06307_),
    .X(_06332_));
 sky130_fd_sc_hd__xnor2_1 _11862_ (.A(\genblk2.pcpi_div.divisor[8] ),
    .B(\genblk2.pcpi_div.dividend[8] ),
    .Y(_06333_));
 sky130_fd_sc_hd__and2_1 _11863_ (.A(_06332_),
    .B(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__a21o_1 _11864_ (.A1(_02361_),
    .A2(\genblk2.pcpi_div.dividend[8] ),
    .B1(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__or3b_1 _11865_ (.A(\genblk2.pcpi_div.divisor[8] ),
    .B(_06305_),
    .C_N(\genblk2.pcpi_div.dividend[8] ),
    .X(_06336_));
 sky130_fd_sc_hd__and2b_1 _11866_ (.A_N(_06306_),
    .B(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__nor2_1 _11867_ (.A(_06305_),
    .B(_06306_),
    .Y(_06338_));
 sky130_fd_sc_hd__a21bo_1 _11868_ (.A1(_06334_),
    .A2(_06338_),
    .B1_N(_06337_),
    .X(_06339_));
 sky130_fd_sc_hd__a21boi_1 _11869_ (.A1(_06304_),
    .A2(_06339_),
    .B1_N(_06303_),
    .Y(_06340_));
 sky130_fd_sc_hd__nor2_1 _11870_ (.A(_06300_),
    .B(_06302_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand2_1 _11871_ (.A(_06304_),
    .B(_06341_),
    .Y(_06342_));
 sky130_fd_sc_hd__o221a_1 _11872_ (.A1(_06302_),
    .A2(_06303_),
    .B1(_06337_),
    .B2(_06342_),
    .C1(_06301_),
    .X(_06343_));
 sky130_fd_sc_hd__or4b_1 _11873_ (.A(_06305_),
    .B(_06342_),
    .C(_06306_),
    .D_N(_06333_),
    .X(_06344_));
 sky130_fd_sc_hd__nand2b_1 _11874_ (.A_N(_06344_),
    .B(_06332_),
    .Y(_06345_));
 sky130_fd_sc_hd__a21o_1 _11875_ (.A1(_06343_),
    .A2(_06345_),
    .B1(_06299_),
    .X(_06346_));
 sky130_fd_sc_hd__a31o_1 _11876_ (.A1(_06296_),
    .A2(_06297_),
    .A3(_06346_),
    .B1(_06295_),
    .X(_06347_));
 sky130_fd_sc_hd__or2_1 _11877_ (.A(_06294_),
    .B(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__o21ai_1 _11878_ (.A1(\genblk2.pcpi_div.divisor[14] ),
    .A2(_02390_),
    .B1(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__nand2b_1 _11879_ (.A_N(_06292_),
    .B(_06293_),
    .Y(_06350_));
 sky130_fd_sc_hd__or2_1 _11880_ (.A(_06294_),
    .B(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__nand2b_1 _11881_ (.A_N(_06295_),
    .B(_06296_),
    .Y(_06352_));
 sky130_fd_sc_hd__or3_1 _11882_ (.A(_06299_),
    .B(_06351_),
    .C(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__nor2_1 _11883_ (.A(_06344_),
    .B(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__o2bb2a_1 _11884_ (.A1_N(_06332_),
    .A2_N(_06354_),
    .B1(_06343_),
    .B2(_06353_),
    .X(_06355_));
 sky130_fd_sc_hd__a211o_1 _11885_ (.A1(_06296_),
    .A2(_06297_),
    .B1(_06351_),
    .C1(_06295_),
    .X(_06356_));
 sky130_fd_sc_hd__o311a_1 _11886_ (.A1(\genblk2.pcpi_div.divisor[14] ),
    .A2(_02390_),
    .A3(_06292_),
    .B1(_06293_),
    .C1(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__a21o_1 _11887_ (.A1(_06355_),
    .A2(_06357_),
    .B1(_06291_),
    .X(_06358_));
 sky130_fd_sc_hd__a21oi_1 _11888_ (.A1(_06289_),
    .A2(_06358_),
    .B1(_06287_),
    .Y(_06359_));
 sky130_fd_sc_hd__or4_1 _11889_ (.A(_06283_),
    .B(_06285_),
    .C(_06287_),
    .D(_06289_),
    .X(_06360_));
 sky130_fd_sc_hd__nand2_1 _11890_ (.A(_06286_),
    .B(_06290_),
    .Y(_06361_));
 sky130_fd_sc_hd__o211ai_2 _11891_ (.A1(_06358_),
    .A2(_06361_),
    .B1(_06360_),
    .C1(_06282_),
    .Y(_06362_));
 sky130_fd_sc_hd__nand2_1 _11892_ (.A(_06278_),
    .B(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__or4bb_1 _11893_ (.A(_06274_),
    .B(_06277_),
    .C_N(_06278_),
    .D_N(_06362_),
    .X(_06364_));
 sky130_fd_sc_hd__o21ba_1 _11894_ (.A1(_06271_),
    .A2(_06272_),
    .B1_N(_06270_),
    .X(_06365_));
 sky130_fd_sc_hd__a21oi_1 _11895_ (.A1(_02359_),
    .A2(\genblk2.pcpi_div.dividend[20] ),
    .B1(_06275_),
    .Y(_06366_));
 sky130_fd_sc_hd__o31a_1 _11896_ (.A1(_06274_),
    .A2(_06276_),
    .A3(_06366_),
    .B1(_06365_),
    .X(_06367_));
 sky130_fd_sc_hd__and2_1 _11897_ (.A(_06364_),
    .B(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__a21bo_1 _11898_ (.A1(_06364_),
    .A2(_06367_),
    .B1_N(_06269_),
    .X(_06369_));
 sky130_fd_sc_hd__and2b_1 _11899_ (.A_N(\genblk2.pcpi_div.dividend[27] ),
    .B(\genblk2.pcpi_div.divisor[27] ),
    .X(_06370_));
 sky130_fd_sc_hd__nand2b_1 _11900_ (.A_N(\genblk2.pcpi_div.divisor[27] ),
    .B(\genblk2.pcpi_div.dividend[27] ),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2b_1 _11901_ (.A_N(_06370_),
    .B(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__nand2b_1 _11902_ (.A_N(\genblk2.pcpi_div.divisor[26] ),
    .B(\genblk2.pcpi_div.dividend[26] ),
    .Y(_06373_));
 sky130_fd_sc_hd__nand2b_1 _11903_ (.A_N(\genblk2.pcpi_div.dividend[26] ),
    .B(\genblk2.pcpi_div.divisor[26] ),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_1 _11904_ (.A(_06373_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__or2_1 _11905_ (.A(_06372_),
    .B(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__and2b_1 _11906_ (.A_N(\genblk2.pcpi_div.dividend[25] ),
    .B(\genblk2.pcpi_div.divisor[25] ),
    .X(_06377_));
 sky130_fd_sc_hd__and2b_1 _11907_ (.A_N(\genblk2.pcpi_div.divisor[25] ),
    .B(\genblk2.pcpi_div.dividend[25] ),
    .X(_06378_));
 sky130_fd_sc_hd__or2_1 _11908_ (.A(_06377_),
    .B(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__nor2_1 _11909_ (.A(_06267_),
    .B(_06378_),
    .Y(_06380_));
 sky130_fd_sc_hd__a21o_1 _11910_ (.A1(_06371_),
    .A2(_06373_),
    .B1(_06370_),
    .X(_06381_));
 sky130_fd_sc_hd__o31a_1 _11911_ (.A1(_06376_),
    .A2(_06377_),
    .A3(_06380_),
    .B1(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__o31a_1 _11912_ (.A1(_06369_),
    .A2(_06376_),
    .A3(_06379_),
    .B1(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__o21ba_1 _11913_ (.A1(_06265_),
    .A2(_06383_),
    .B1_N(_06264_),
    .X(_06384_));
 sky130_fd_sc_hd__nand2_1 _11914_ (.A(_06261_),
    .B(_06263_),
    .Y(_06385_));
 sky130_fd_sc_hd__a21o_1 _11915_ (.A1(_06263_),
    .A2(_06384_),
    .B1(_06262_),
    .X(_06386_));
 sky130_fd_sc_hd__a211o_1 _11916_ (.A1(_06263_),
    .A2(_06384_),
    .B1(_06260_),
    .C1(_06262_),
    .X(_06387_));
 sky130_fd_sc_hd__o21ai_1 _11917_ (.A1(\genblk2.pcpi_div.divisor[30] ),
    .A2(_02389_),
    .B1(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__or3_1 _11918_ (.A(\genblk2.pcpi_div.divisor[61] ),
    .B(\genblk2.pcpi_div.divisor[60] ),
    .C(\genblk2.pcpi_div.divisor[62] ),
    .X(_06389_));
 sky130_fd_sc_hd__or4_1 _11919_ (.A(\genblk2.pcpi_div.divisor[59] ),
    .B(\genblk2.pcpi_div.divisor[58] ),
    .C(\genblk2.pcpi_div.divisor[57] ),
    .D(\genblk2.pcpi_div.divisor[56] ),
    .X(_06390_));
 sky130_fd_sc_hd__or4_1 _11920_ (.A(\genblk2.pcpi_div.divisor[51] ),
    .B(\genblk2.pcpi_div.divisor[50] ),
    .C(\genblk2.pcpi_div.divisor[49] ),
    .D(\genblk2.pcpi_div.divisor[48] ),
    .X(_06391_));
 sky130_fd_sc_hd__or4_1 _11921_ (.A(\genblk2.pcpi_div.divisor[47] ),
    .B(\genblk2.pcpi_div.divisor[46] ),
    .C(\genblk2.pcpi_div.divisor[45] ),
    .D(\genblk2.pcpi_div.divisor[44] ),
    .X(_06392_));
 sky130_fd_sc_hd__and2b_1 _11922_ (.A_N(\genblk2.pcpi_div.dividend[31] ),
    .B(\genblk2.pcpi_div.divisor[31] ),
    .X(_06393_));
 sky130_fd_sc_hd__or4_1 _11923_ (.A(\genblk2.pcpi_div.divisor[39] ),
    .B(\genblk2.pcpi_div.divisor[38] ),
    .C(\genblk2.pcpi_div.divisor[37] ),
    .D(\genblk2.pcpi_div.divisor[36] ),
    .X(_06394_));
 sky130_fd_sc_hd__or4_1 _11924_ (.A(\genblk2.pcpi_div.divisor[43] ),
    .B(\genblk2.pcpi_div.divisor[42] ),
    .C(\genblk2.pcpi_div.divisor[41] ),
    .D(\genblk2.pcpi_div.divisor[40] ),
    .X(_06395_));
 sky130_fd_sc_hd__or4_1 _11925_ (.A(\genblk2.pcpi_div.divisor[55] ),
    .B(\genblk2.pcpi_div.divisor[54] ),
    .C(\genblk2.pcpi_div.divisor[53] ),
    .D(\genblk2.pcpi_div.divisor[52] ),
    .X(_06396_));
 sky130_fd_sc_hd__or4_1 _11926_ (.A(\genblk2.pcpi_div.divisor[35] ),
    .B(\genblk2.pcpi_div.divisor[34] ),
    .C(\genblk2.pcpi_div.divisor[33] ),
    .D(\genblk2.pcpi_div.divisor[32] ),
    .X(_06397_));
 sky130_fd_sc_hd__or4_2 _11927_ (.A(_06389_),
    .B(_06390_),
    .C(_06391_),
    .D(_06396_),
    .X(_06398_));
 sky130_fd_sc_hd__or4_1 _11928_ (.A(_06392_),
    .B(_06394_),
    .C(_06395_),
    .D(_06397_),
    .X(_06399_));
 sky130_fd_sc_hd__nor3_1 _11929_ (.A(_06393_),
    .B(_06398_),
    .C(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__nor2_1 _11930_ (.A(_06259_),
    .B(_06393_),
    .Y(_06401_));
 sky130_fd_sc_hd__o21ai_1 _11931_ (.A1(_06259_),
    .A2(_06388_),
    .B1(_06400_),
    .Y(_06402_));
 sky130_fd_sc_hd__a21oi_2 _11932_ (.A1(_06258_),
    .A2(_06402_),
    .B1(net384),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2b_1 _11933_ (.A_N(\genblk2.pcpi_div.divisor[0] ),
    .B(\genblk2.pcpi_div.dividend[0] ),
    .Y(_06404_));
 sky130_fd_sc_hd__and3_1 _11934_ (.A(net866),
    .B(_06320_),
    .C(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__a21oi_1 _11935_ (.A1(_02384_),
    .A2(net873),
    .B1(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(\genblk2.pcpi_div.dividend[0] ),
    .A1(_06406_),
    .S(net276),
    .X(_01009_));
 sky130_fd_sc_hd__nor2_1 _11937_ (.A(_06320_),
    .B(_06321_),
    .Y(_06407_));
 sky130_fd_sc_hd__nor2_1 _11938_ (.A(_06322_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__and2_2 _11939_ (.A(net1189),
    .B(_02507_),
    .X(_06409_));
 sky130_fd_sc_hd__a21oi_1 _11940_ (.A1(net1052),
    .A2(net726),
    .B1(net1049),
    .Y(_06410_));
 sky130_fd_sc_hd__a31o_1 _11941_ (.A1(net1049),
    .A2(net1052),
    .A3(net726),
    .B1(net866),
    .X(_06411_));
 sky130_fd_sc_hd__a2bb2o_1 _11942_ (.A1_N(_06411_),
    .A2_N(_06410_),
    .B1(_06408_),
    .B2(net866),
    .X(_06412_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(\genblk2.pcpi_div.dividend[1] ),
    .A1(_06412_),
    .S(net276),
    .X(_01010_));
 sky130_fd_sc_hd__a21oi_1 _11944_ (.A1(_02443_),
    .A2(net726),
    .B1(net1046),
    .Y(_06413_));
 sky130_fd_sc_hd__a31o_1 _11945_ (.A1(net1046),
    .A2(_02443_),
    .A3(net726),
    .B1(net866),
    .X(_06414_));
 sky130_fd_sc_hd__a211o_1 _11946_ (.A1(_06317_),
    .A2(_06318_),
    .B1(_06319_),
    .C1(_06322_),
    .X(_06415_));
 sky130_fd_sc_hd__or3b_1 _11947_ (.A(net873),
    .B(_06323_),
    .C_N(_06415_),
    .X(_06416_));
 sky130_fd_sc_hd__o21ai_1 _11948_ (.A1(_06413_),
    .A2(_06414_),
    .B1(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(\genblk2.pcpi_div.dividend[2] ),
    .A1(_06417_),
    .S(net277),
    .X(_01011_));
 sky130_fd_sc_hd__a211o_1 _11950_ (.A1(_06315_),
    .A2(_06324_),
    .B1(_06323_),
    .C1(_06316_),
    .X(_06418_));
 sky130_fd_sc_hd__nor2_1 _11951_ (.A(net873),
    .B(_06325_),
    .Y(_06419_));
 sky130_fd_sc_hd__o21a_1 _11952_ (.A1(net1046),
    .A2(_02443_),
    .B1(_06409_),
    .X(_06420_));
 sky130_fd_sc_hd__xnor2_1 _11953_ (.A(_02402_),
    .B(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__a22o_1 _11954_ (.A1(_06418_),
    .A2(_06419_),
    .B1(_06421_),
    .B2(net873),
    .X(_06422_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(\genblk2.pcpi_div.dividend[3] ),
    .A1(_06422_),
    .S(net277),
    .X(_01012_));
 sky130_fd_sc_hd__or3_2 _11956_ (.A(net1046),
    .B(net228),
    .C(_02443_),
    .X(_06423_));
 sky130_fd_sc_hd__a21o_1 _11957_ (.A1(net726),
    .A2(_06423_),
    .B1(net1043),
    .X(_06424_));
 sky130_fd_sc_hd__a31oi_1 _11958_ (.A1(net1043),
    .A2(net726),
    .A3(_06423_),
    .B1(net866),
    .Y(_06425_));
 sky130_fd_sc_hd__a211o_1 _11959_ (.A1(_06312_),
    .A2(_06313_),
    .B1(_06314_),
    .C1(_06325_),
    .X(_06426_));
 sky130_fd_sc_hd__a32o_1 _11960_ (.A1(net866),
    .A2(_06326_),
    .A3(_06426_),
    .B1(_06425_),
    .B2(_06424_),
    .X(_06427_));
 sky130_fd_sc_hd__mux2_1 _11961_ (.A0(\genblk2.pcpi_div.dividend[4] ),
    .A1(_06427_),
    .S(net276),
    .X(_01013_));
 sky130_fd_sc_hd__nor2_1 _11962_ (.A(_06309_),
    .B(_06311_),
    .Y(_06428_));
 sky130_fd_sc_hd__xnor2_1 _11963_ (.A(_06327_),
    .B(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__o21ai_1 _11964_ (.A1(net1043),
    .A2(_06423_),
    .B1(net726),
    .Y(_06430_));
 sky130_fd_sc_hd__xnor2_1 _11965_ (.A(net1041),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__mux2_1 _11966_ (.A0(_06429_),
    .A1(_06431_),
    .S(net868),
    .X(_06432_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(net3010),
    .A1(_06432_),
    .S(net276),
    .X(_01014_));
 sky130_fd_sc_hd__o211ai_1 _11968_ (.A1(_06311_),
    .A2(_06327_),
    .B1(_06308_),
    .C1(_06310_),
    .Y(_06433_));
 sky130_fd_sc_hd__or3_2 _11969_ (.A(net1043),
    .B(net1041),
    .C(_06423_),
    .X(_06434_));
 sky130_fd_sc_hd__a21o_1 _11970_ (.A1(net726),
    .A2(_06434_),
    .B1(net1039),
    .X(_06435_));
 sky130_fd_sc_hd__nand3_1 _11971_ (.A(net1039),
    .B(net726),
    .C(_06434_),
    .Y(_06436_));
 sky130_fd_sc_hd__and3_1 _11972_ (.A(net868),
    .B(_06435_),
    .C(_06436_),
    .X(_06437_));
 sky130_fd_sc_hd__a31o_1 _11973_ (.A1(net865),
    .A2(_06328_),
    .A3(_06433_),
    .B1(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__mux2_1 _11974_ (.A0(\genblk2.pcpi_div.dividend[6] ),
    .A1(_06438_),
    .S(net276),
    .X(_01015_));
 sky130_fd_sc_hd__xnor2_1 _11975_ (.A(_06329_),
    .B(_06331_),
    .Y(_06439_));
 sky130_fd_sc_hd__o21a_1 _11976_ (.A1(net1039),
    .A2(_06434_),
    .B1(net726),
    .X(_06440_));
 sky130_fd_sc_hd__nand2_1 _11977_ (.A(net1036),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__o21a_1 _11978_ (.A1(net1036),
    .A2(_06440_),
    .B1(net868),
    .X(_06442_));
 sky130_fd_sc_hd__a22o_1 _11979_ (.A1(net865),
    .A2(_06439_),
    .B1(_06441_),
    .B2(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__mux2_1 _11980_ (.A0(\genblk2.pcpi_div.dividend[7] ),
    .A1(_06443_),
    .S(net271),
    .X(_01016_));
 sky130_fd_sc_hd__o31a_1 _11981_ (.A1(net1039),
    .A2(net1036),
    .A3(_06434_),
    .B1(net723),
    .X(_06444_));
 sky130_fd_sc_hd__xor2_1 _11982_ (.A(net1034),
    .B(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__o21ai_1 _11983_ (.A1(_06332_),
    .A2(_06333_),
    .B1(net862),
    .Y(_06446_));
 sky130_fd_sc_hd__a2bb2o_1 _11984_ (.A1_N(_06334_),
    .A2_N(_06446_),
    .B1(_06445_),
    .B2(net867),
    .X(_06447_));
 sky130_fd_sc_hd__mux2_1 _11985_ (.A0(\genblk2.pcpi_div.dividend[8] ),
    .A1(_06447_),
    .S(net271),
    .X(_01017_));
 sky130_fd_sc_hd__or4_2 _11986_ (.A(net1039),
    .B(net1036),
    .C(net1034),
    .D(_06434_),
    .X(_06448_));
 sky130_fd_sc_hd__a21oi_1 _11987_ (.A1(net723),
    .A2(_06448_),
    .B1(net1031),
    .Y(_06449_));
 sky130_fd_sc_hd__a31o_1 _11988_ (.A1(net1032),
    .A2(net723),
    .A3(_06448_),
    .B1(net862),
    .X(_06450_));
 sky130_fd_sc_hd__xnor2_1 _11989_ (.A(_06335_),
    .B(_06338_),
    .Y(_06451_));
 sky130_fd_sc_hd__o221a_1 _11990_ (.A1(_06449_),
    .A2(_06450_),
    .B1(_06451_),
    .B2(net867),
    .C1(net271),
    .X(_06452_));
 sky130_fd_sc_hd__o21ba_1 _11991_ (.A1(\genblk2.pcpi_div.dividend[9] ),
    .A2(net271),
    .B1_N(_06452_),
    .X(_01018_));
 sky130_fd_sc_hd__o21a_1 _11992_ (.A1(net1032),
    .A2(_06448_),
    .B1(net723),
    .X(_06453_));
 sky130_fd_sc_hd__xnor2_1 _11993_ (.A(net1030),
    .B(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__nor2_1 _11994_ (.A(net862),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__xnor2_1 _11995_ (.A(_06304_),
    .B(_06339_),
    .Y(_06456_));
 sky130_fd_sc_hd__o21ai_1 _11996_ (.A1(net867),
    .A2(_06456_),
    .B1(net271),
    .Y(_06457_));
 sky130_fd_sc_hd__o22a_1 _11997_ (.A1(\genblk2.pcpi_div.dividend[10] ),
    .A2(net271),
    .B1(_06455_),
    .B2(_06457_),
    .X(_01019_));
 sky130_fd_sc_hd__xnor2_1 _11998_ (.A(_06340_),
    .B(_06341_),
    .Y(_06458_));
 sky130_fd_sc_hd__or3_1 _11999_ (.A(net1032),
    .B(net1030),
    .C(_06448_),
    .X(_06459_));
 sky130_fd_sc_hd__a21oi_1 _12000_ (.A1(net723),
    .A2(_06459_),
    .B1(net1028),
    .Y(_06460_));
 sky130_fd_sc_hd__a31o_1 _12001_ (.A1(net1028),
    .A2(net723),
    .A3(_06459_),
    .B1(net862),
    .X(_06461_));
 sky130_fd_sc_hd__a2bb2o_1 _12002_ (.A1_N(_06461_),
    .A2_N(_06460_),
    .B1(_06458_),
    .B2(net862),
    .X(_06462_));
 sky130_fd_sc_hd__mux2_1 _12003_ (.A0(\genblk2.pcpi_div.dividend[11] ),
    .A1(_06462_),
    .S(net271),
    .X(_01020_));
 sky130_fd_sc_hd__nand3_1 _12004_ (.A(_06299_),
    .B(_06343_),
    .C(_06345_),
    .Y(_06463_));
 sky130_fd_sc_hd__or2_1 _12005_ (.A(net205),
    .B(_06459_),
    .X(_06464_));
 sky130_fd_sc_hd__a21o_1 _12006_ (.A1(net723),
    .A2(_06464_),
    .B1(net1026),
    .X(_06465_));
 sky130_fd_sc_hd__a31oi_1 _12007_ (.A1(net1027),
    .A2(net723),
    .A3(_06464_),
    .B1(net862),
    .Y(_06466_));
 sky130_fd_sc_hd__a32o_1 _12008_ (.A1(net862),
    .A2(_06346_),
    .A3(_06463_),
    .B1(_06465_),
    .B2(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__mux2_1 _12009_ (.A0(\genblk2.pcpi_div.dividend[12] ),
    .A1(_06467_),
    .S(net271),
    .X(_01021_));
 sky130_fd_sc_hd__a21oi_1 _12010_ (.A1(_06297_),
    .A2(_06346_),
    .B1(_06352_),
    .Y(_06468_));
 sky130_fd_sc_hd__and3_1 _12011_ (.A(_06297_),
    .B(_06346_),
    .C(_06352_),
    .X(_06469_));
 sky130_fd_sc_hd__or2_1 _12012_ (.A(net1027),
    .B(_06464_),
    .X(_06470_));
 sky130_fd_sc_hd__a21oi_1 _12013_ (.A1(net721),
    .A2(_06470_),
    .B1(net1024),
    .Y(_06471_));
 sky130_fd_sc_hd__a311o_1 _12014_ (.A1(net1025),
    .A2(net721),
    .A3(_06470_),
    .B1(_06471_),
    .C1(net862),
    .X(_06472_));
 sky130_fd_sc_hd__o31ai_1 _12015_ (.A1(net867),
    .A2(_06468_),
    .A3(_06469_),
    .B1(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__mux2_1 _12016_ (.A0(net3020),
    .A1(_06473_),
    .S(net269),
    .X(_01022_));
 sky130_fd_sc_hd__o21a_1 _12017_ (.A1(net1025),
    .A2(_06470_),
    .B1(net721),
    .X(_06474_));
 sky130_fd_sc_hd__o21ai_1 _12018_ (.A1(net1023),
    .A2(_06474_),
    .B1(net867),
    .Y(_06475_));
 sky130_fd_sc_hd__a21oi_1 _12019_ (.A1(net1023),
    .A2(_06474_),
    .B1(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__nand2_1 _12020_ (.A(_06294_),
    .B(_06347_),
    .Y(_06477_));
 sky130_fd_sc_hd__a31o_1 _12021_ (.A1(net861),
    .A2(_06348_),
    .A3(_06477_),
    .B1(_06476_),
    .X(_06478_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(net3043),
    .A1(_06478_),
    .S(net269),
    .X(_01023_));
 sky130_fd_sc_hd__xnor2_1 _12023_ (.A(_06349_),
    .B(_06350_),
    .Y(_06479_));
 sky130_fd_sc_hd__or3_1 _12024_ (.A(net1025),
    .B(net1023),
    .C(_06470_),
    .X(_06480_));
 sky130_fd_sc_hd__a21oi_1 _12025_ (.A1(net721),
    .A2(_06480_),
    .B1(net1021),
    .Y(_06481_));
 sky130_fd_sc_hd__a31o_1 _12026_ (.A1(net1021),
    .A2(net721),
    .A3(_06480_),
    .B1(net861),
    .X(_06482_));
 sky130_fd_sc_hd__a2bb2o_1 _12027_ (.A1_N(_06482_),
    .A2_N(_06481_),
    .B1(_06479_),
    .B2(net861),
    .X(_06483_));
 sky130_fd_sc_hd__mux2_1 _12028_ (.A0(\genblk2.pcpi_div.dividend[15] ),
    .A1(_06483_),
    .S(net269),
    .X(_01024_));
 sky130_fd_sc_hd__or2_1 _12029_ (.A(net1021),
    .B(_06480_),
    .X(_06484_));
 sky130_fd_sc_hd__a21oi_1 _12030_ (.A1(net722),
    .A2(_06484_),
    .B1(net1019),
    .Y(_06485_));
 sky130_fd_sc_hd__a31o_1 _12031_ (.A1(net1019),
    .A2(net722),
    .A3(_06484_),
    .B1(net862),
    .X(_06486_));
 sky130_fd_sc_hd__nor2_1 _12032_ (.A(_06485_),
    .B(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nand3_1 _12033_ (.A(_06291_),
    .B(_06355_),
    .C(_06357_),
    .Y(_06488_));
 sky130_fd_sc_hd__a31o_1 _12034_ (.A1(net861),
    .A2(_06358_),
    .A3(_06488_),
    .B1(_06487_),
    .X(_06489_));
 sky130_fd_sc_hd__mux2_1 _12035_ (.A0(\genblk2.pcpi_div.dividend[16] ),
    .A1(_06489_),
    .S(net269),
    .X(_01025_));
 sky130_fd_sc_hd__a21bo_1 _12036_ (.A1(_02360_),
    .A2(\genblk2.pcpi_div.dividend[16] ),
    .B1_N(_06358_),
    .X(_06490_));
 sky130_fd_sc_hd__xor2_1 _12037_ (.A(_06290_),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__or2_1 _12038_ (.A(net1019),
    .B(_06484_),
    .X(_06492_));
 sky130_fd_sc_hd__a21oi_1 _12039_ (.A1(net721),
    .A2(_06492_),
    .B1(net1016),
    .Y(_06493_));
 sky130_fd_sc_hd__a31o_1 _12040_ (.A1(net1016),
    .A2(net721),
    .A3(_06492_),
    .B1(net861),
    .X(_06494_));
 sky130_fd_sc_hd__a2bb2o_1 _12041_ (.A1_N(_06494_),
    .A2_N(_06493_),
    .B1(_06491_),
    .B2(net861),
    .X(_06495_));
 sky130_fd_sc_hd__mux2_1 _12042_ (.A0(\genblk2.pcpi_div.dividend[17] ),
    .A1(_06495_),
    .S(net269),
    .X(_01026_));
 sky130_fd_sc_hd__o21ai_1 _12043_ (.A1(net1016),
    .A2(_06492_),
    .B1(net721),
    .Y(_06496_));
 sky130_fd_sc_hd__xnor2_1 _12044_ (.A(net1015),
    .B(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__nand2b_1 _12045_ (.A_N(_06285_),
    .B(_06359_),
    .Y(_06498_));
 sky130_fd_sc_hd__xnor2_1 _12046_ (.A(_06285_),
    .B(_06359_),
    .Y(_06499_));
 sky130_fd_sc_hd__mux2_1 _12047_ (.A0(_06497_),
    .A1(_06499_),
    .S(net861),
    .X(_06500_));
 sky130_fd_sc_hd__mux2_1 _12048_ (.A0(net3021),
    .A1(_06500_),
    .S(net269),
    .X(_01027_));
 sky130_fd_sc_hd__or4_1 _12049_ (.A(net1019),
    .B(net1016),
    .C(net1015),
    .D(_06484_),
    .X(_06501_));
 sky130_fd_sc_hd__and3_1 _12050_ (.A(net1013),
    .B(net722),
    .C(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__a21oi_1 _12051_ (.A1(net722),
    .A2(_06501_),
    .B1(net1013),
    .Y(_06503_));
 sky130_fd_sc_hd__or3_1 _12052_ (.A(net861),
    .B(_06502_),
    .C(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__a21oi_1 _12053_ (.A1(_06280_),
    .A2(_06498_),
    .B1(_06283_),
    .Y(_06505_));
 sky130_fd_sc_hd__a31o_1 _12054_ (.A1(_06280_),
    .A2(_06283_),
    .A3(_06498_),
    .B1(net867),
    .X(_06506_));
 sky130_fd_sc_hd__o211a_1 _12055_ (.A1(_06505_),
    .A2(_06506_),
    .B1(net269),
    .C1(_06504_),
    .X(_06507_));
 sky130_fd_sc_hd__o21ba_1 _12056_ (.A1(\genblk2.pcpi_div.dividend[19] ),
    .A2(net269),
    .B1_N(_06507_),
    .X(_01028_));
 sky130_fd_sc_hd__or2_1 _12057_ (.A(net1013),
    .B(_06501_),
    .X(_06508_));
 sky130_fd_sc_hd__nand3_1 _12058_ (.A(net1011),
    .B(net721),
    .C(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__a21o_1 _12059_ (.A1(net721),
    .A2(_06508_),
    .B1(net1011),
    .X(_06510_));
 sky130_fd_sc_hd__and3_1 _12060_ (.A(net867),
    .B(_06509_),
    .C(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__or2_1 _12061_ (.A(_06278_),
    .B(_06362_),
    .X(_06512_));
 sky130_fd_sc_hd__a31o_1 _12062_ (.A1(net863),
    .A2(_06363_),
    .A3(_06512_),
    .B1(_06511_),
    .X(_06513_));
 sky130_fd_sc_hd__mux2_1 _12063_ (.A0(\genblk2.pcpi_div.dividend[20] ),
    .A1(_06513_),
    .S(net269),
    .X(_01029_));
 sky130_fd_sc_hd__a21bo_1 _12064_ (.A1(_02359_),
    .A2(\genblk2.pcpi_div.dividend[20] ),
    .B1_N(_06363_),
    .X(_06514_));
 sky130_fd_sc_hd__xnor2_1 _12065_ (.A(_06277_),
    .B(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__or2_1 _12066_ (.A(net1011),
    .B(_06508_),
    .X(_06516_));
 sky130_fd_sc_hd__a21oi_1 _12067_ (.A1(net722),
    .A2(_06516_),
    .B1(net1009),
    .Y(_06517_));
 sky130_fd_sc_hd__a31o_1 _12068_ (.A1(net1009),
    .A2(net722),
    .A3(_06516_),
    .B1(net861),
    .X(_06518_));
 sky130_fd_sc_hd__a2bb2o_1 _12069_ (.A1_N(_06518_),
    .A2_N(_06517_),
    .B1(_06515_),
    .B2(net861),
    .X(_06519_));
 sky130_fd_sc_hd__mux2_1 _12070_ (.A0(\genblk2.pcpi_div.dividend[21] ),
    .A1(_06519_),
    .S(net270),
    .X(_01030_));
 sky130_fd_sc_hd__and2b_1 _12071_ (.A_N(_06276_),
    .B(_06514_),
    .X(_06520_));
 sky130_fd_sc_hd__o21ai_1 _12072_ (.A1(_06275_),
    .A2(_06520_),
    .B1(_06273_),
    .Y(_06521_));
 sky130_fd_sc_hd__or3_1 _12073_ (.A(_06273_),
    .B(_06275_),
    .C(_06520_),
    .X(_06522_));
 sky130_fd_sc_hd__or3_1 _12074_ (.A(net1011),
    .B(net1009),
    .C(_06508_),
    .X(_06523_));
 sky130_fd_sc_hd__a21oi_1 _12075_ (.A1(net724),
    .A2(_06523_),
    .B1(net1008),
    .Y(_06524_));
 sky130_fd_sc_hd__a31o_1 _12076_ (.A1(net1008),
    .A2(net724),
    .A3(_06523_),
    .B1(net863),
    .X(_06525_));
 sky130_fd_sc_hd__nor2_1 _12077_ (.A(_06524_),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__a31o_1 _12078_ (.A1(net863),
    .A2(_06521_),
    .A3(_06522_),
    .B1(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__mux2_1 _12079_ (.A0(\genblk2.pcpi_div.dividend[22] ),
    .A1(_06527_),
    .S(net273),
    .X(_01031_));
 sky130_fd_sc_hd__or2_1 _12080_ (.A(net1008),
    .B(_06523_),
    .X(_06528_));
 sky130_fd_sc_hd__a21oi_1 _12081_ (.A1(net724),
    .A2(_06528_),
    .B1(net1006),
    .Y(_06529_));
 sky130_fd_sc_hd__a31o_1 _12082_ (.A1(net1006),
    .A2(net724),
    .A3(_06528_),
    .B1(net863),
    .X(_06530_));
 sky130_fd_sc_hd__nor2_1 _12083_ (.A(_06529_),
    .B(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__o211ai_1 _12084_ (.A1(_06270_),
    .A2(_06271_),
    .B1(_06272_),
    .C1(_06521_),
    .Y(_06532_));
 sky130_fd_sc_hd__a211o_1 _12085_ (.A1(_06272_),
    .A2(_06521_),
    .B1(_06270_),
    .C1(_06271_),
    .X(_06533_));
 sky130_fd_sc_hd__a31o_1 _12086_ (.A1(net863),
    .A2(_06532_),
    .A3(_06533_),
    .B1(_06531_),
    .X(_06534_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(net3050),
    .A1(_06534_),
    .S(net273),
    .X(_01032_));
 sky130_fd_sc_hd__xnor2_1 _12088_ (.A(_06269_),
    .B(_06368_),
    .Y(_06535_));
 sky130_fd_sc_hd__or2_1 _12089_ (.A(net1006),
    .B(_06528_),
    .X(_06536_));
 sky130_fd_sc_hd__a21oi_1 _12090_ (.A1(net724),
    .A2(_06536_),
    .B1(net1005),
    .Y(_06537_));
 sky130_fd_sc_hd__a31o_1 _12091_ (.A1(net1005),
    .A2(net724),
    .A3(_06536_),
    .B1(net863),
    .X(_06538_));
 sky130_fd_sc_hd__a2bb2o_1 _12092_ (.A1_N(_06538_),
    .A2_N(_06537_),
    .B1(_06535_),
    .B2(net863),
    .X(_06539_));
 sky130_fd_sc_hd__mux2_1 _12093_ (.A0(\genblk2.pcpi_div.dividend[24] ),
    .A1(_06539_),
    .S(net273),
    .X(_01033_));
 sky130_fd_sc_hd__and2b_1 _12094_ (.A_N(_06267_),
    .B(_06369_),
    .X(_06540_));
 sky130_fd_sc_hd__xnor2_1 _12095_ (.A(_06379_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__or2_1 _12096_ (.A(net1005),
    .B(_06536_),
    .X(_06542_));
 sky130_fd_sc_hd__a21oi_1 _12097_ (.A1(net724),
    .A2(_06542_),
    .B1(net1003),
    .Y(_06543_));
 sky130_fd_sc_hd__a31o_1 _12098_ (.A1(net1003),
    .A2(net724),
    .A3(_06542_),
    .B1(net863),
    .X(_06544_));
 sky130_fd_sc_hd__o221a_1 _12099_ (.A1(net867),
    .A2(_06541_),
    .B1(_06543_),
    .B2(_06544_),
    .C1(net275),
    .X(_06545_));
 sky130_fd_sc_hd__o21ba_1 _12100_ (.A1(\genblk2.pcpi_div.dividend[25] ),
    .A2(net273),
    .B1_N(_06545_),
    .X(_01034_));
 sky130_fd_sc_hd__a21o_1 _12101_ (.A1(_06369_),
    .A2(_06380_),
    .B1(_06377_),
    .X(_06546_));
 sky130_fd_sc_hd__nand2_1 _12102_ (.A(_06375_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__or2_1 _12103_ (.A(_06375_),
    .B(_06546_),
    .X(_06548_));
 sky130_fd_sc_hd__or2_1 _12104_ (.A(net1003),
    .B(_06542_),
    .X(_06549_));
 sky130_fd_sc_hd__a21o_1 _12105_ (.A1(net724),
    .A2(_06549_),
    .B1(net1001),
    .X(_06550_));
 sky130_fd_sc_hd__a31oi_1 _12106_ (.A1(net1001),
    .A2(net725),
    .A3(_06549_),
    .B1(net863),
    .Y(_06551_));
 sky130_fd_sc_hd__a32o_1 _12107_ (.A1(net863),
    .A2(_06547_),
    .A3(_06548_),
    .B1(_06550_),
    .B2(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__mux2_1 _12108_ (.A0(\genblk2.pcpi_div.dividend[26] ),
    .A1(_06552_),
    .S(net273),
    .X(_01035_));
 sky130_fd_sc_hd__a21oi_1 _12109_ (.A1(_06373_),
    .A2(_06548_),
    .B1(_06372_),
    .Y(_06553_));
 sky130_fd_sc_hd__a31o_1 _12110_ (.A1(_06372_),
    .A2(_06373_),
    .A3(_06548_),
    .B1(net869),
    .X(_06554_));
 sky130_fd_sc_hd__o21ai_1 _12111_ (.A1(net1001),
    .A2(_06549_),
    .B1(net724),
    .Y(_06555_));
 sky130_fd_sc_hd__xnor2_1 _12112_ (.A(net999),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__a2bb2o_1 _12113_ (.A1_N(_06553_),
    .A2_N(_06554_),
    .B1(_06556_),
    .B2(net869),
    .X(_06557_));
 sky130_fd_sc_hd__mux2_1 _12114_ (.A0(\genblk2.pcpi_div.dividend[27] ),
    .A1(_06557_),
    .S(net275),
    .X(_01036_));
 sky130_fd_sc_hd__or3_2 _12115_ (.A(net1001),
    .B(net999),
    .C(_06549_),
    .X(_06558_));
 sky130_fd_sc_hd__a21oi_1 _12116_ (.A1(net725),
    .A2(_06558_),
    .B1(net997),
    .Y(_06559_));
 sky130_fd_sc_hd__a31o_1 _12117_ (.A1(net997),
    .A2(net725),
    .A3(_06558_),
    .B1(net864),
    .X(_06560_));
 sky130_fd_sc_hd__xnor2_1 _12118_ (.A(_06266_),
    .B(_06383_),
    .Y(_06561_));
 sky130_fd_sc_hd__o221a_1 _12119_ (.A1(_06559_),
    .A2(_06560_),
    .B1(_06561_),
    .B2(net869),
    .C1(net275),
    .X(_06562_));
 sky130_fd_sc_hd__o21ba_1 _12120_ (.A1(net3033),
    .A2(net274),
    .B1_N(_06562_),
    .X(_01037_));
 sky130_fd_sc_hd__xor2_1 _12121_ (.A(_06384_),
    .B(_06385_),
    .X(_06563_));
 sky130_fd_sc_hd__o21ai_1 _12122_ (.A1(net997),
    .A2(_06558_),
    .B1(net725),
    .Y(_06564_));
 sky130_fd_sc_hd__xnor2_1 _12123_ (.A(net995),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(_06563_),
    .A1(_06565_),
    .S(net869),
    .X(_06566_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(\genblk2.pcpi_div.dividend[29] ),
    .A1(_06566_),
    .S(net274),
    .X(_01038_));
 sky130_fd_sc_hd__or3_1 _12126_ (.A(net997),
    .B(net995),
    .C(_06558_),
    .X(_06567_));
 sky130_fd_sc_hd__a21oi_1 _12127_ (.A1(net725),
    .A2(_06567_),
    .B1(net993),
    .Y(_06568_));
 sky130_fd_sc_hd__a31o_1 _12128_ (.A1(net993),
    .A2(net725),
    .A3(_06567_),
    .B1(net864),
    .X(_06569_));
 sky130_fd_sc_hd__and2_1 _12129_ (.A(_06260_),
    .B(_06386_),
    .X(_06570_));
 sky130_fd_sc_hd__nand2_1 _12130_ (.A(net864),
    .B(_06387_),
    .Y(_06571_));
 sky130_fd_sc_hd__o221a_1 _12131_ (.A1(_06568_),
    .A2(_06569_),
    .B1(_06570_),
    .B2(_06571_),
    .C1(net274),
    .X(_06572_));
 sky130_fd_sc_hd__o21ba_1 _12132_ (.A1(\genblk2.pcpi_div.dividend[30] ),
    .A2(net275),
    .B1_N(_06572_),
    .X(_01039_));
 sky130_fd_sc_hd__o21ai_1 _12133_ (.A1(net993),
    .A2(_06567_),
    .B1(_02507_),
    .Y(_06573_));
 sky130_fd_sc_hd__or2_1 _12134_ (.A(_06388_),
    .B(_06401_),
    .X(_06574_));
 sky130_fd_sc_hd__nand2_1 _12135_ (.A(_06388_),
    .B(_06401_),
    .Y(_06575_));
 sky130_fd_sc_hd__and3_1 _12136_ (.A(net864),
    .B(_06574_),
    .C(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__a31o_1 _12137_ (.A1(net1189),
    .A2(net867),
    .A3(_06573_),
    .B1(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__mux2_1 _12138_ (.A0(net2989),
    .A1(_06577_),
    .S(net274),
    .X(_01040_));
 sky130_fd_sc_hd__a31o_1 _12139_ (.A1(net2663),
    .A2(net1223),
    .A3(_05094_),
    .B1(net749),
    .X(_01041_));
 sky130_fd_sc_hd__and2_1 _12140_ (.A(net1223),
    .B(_06258_),
    .X(_06578_));
 sky130_fd_sc_hd__a22o_1 _12141_ (.A1(net2602),
    .A2(net385),
    .B1(net372),
    .B2(\genblk2.pcpi_div.quotient_msk[1] ),
    .X(_01042_));
 sky130_fd_sc_hd__a22o_1 _12142_ (.A1(\genblk2.pcpi_div.quotient_msk[1] ),
    .A2(net382),
    .B1(net372),
    .B2(net2750),
    .X(_01043_));
 sky130_fd_sc_hd__a22o_1 _12143_ (.A1(net2750),
    .A2(net382),
    .B1(net372),
    .B2(net2858),
    .X(_01044_));
 sky130_fd_sc_hd__a22o_1 _12144_ (.A1(net2858),
    .A2(net383),
    .B1(net371),
    .B2(net2966),
    .X(_01045_));
 sky130_fd_sc_hd__a22o_1 _12145_ (.A1(\genblk2.pcpi_div.quotient_msk[4] ),
    .A2(net382),
    .B1(net371),
    .B2(net2529),
    .X(_01046_));
 sky130_fd_sc_hd__a22o_1 _12146_ (.A1(net2529),
    .A2(net382),
    .B1(net371),
    .B2(net2833),
    .X(_01047_));
 sky130_fd_sc_hd__a22o_1 _12147_ (.A1(net2833),
    .A2(net382),
    .B1(net371),
    .B2(net2909),
    .X(_01048_));
 sky130_fd_sc_hd__a22o_1 _12148_ (.A1(net2909),
    .A2(net382),
    .B1(net366),
    .B2(net2920),
    .X(_01049_));
 sky130_fd_sc_hd__a22o_1 _12149_ (.A1(\genblk2.pcpi_div.quotient_msk[8] ),
    .A2(net382),
    .B1(net367),
    .B2(net2756),
    .X(_01050_));
 sky130_fd_sc_hd__a22o_1 _12150_ (.A1(net2756),
    .A2(net378),
    .B1(net367),
    .B2(net2798),
    .X(_01051_));
 sky130_fd_sc_hd__a22o_1 _12151_ (.A1(net2798),
    .A2(net378),
    .B1(net367),
    .B2(net2866),
    .X(_01052_));
 sky130_fd_sc_hd__a22o_1 _12152_ (.A1(\genblk2.pcpi_div.quotient_msk[11] ),
    .A2(net379),
    .B1(net367),
    .B2(net2803),
    .X(_01053_));
 sky130_fd_sc_hd__a22o_1 _12153_ (.A1(net2803),
    .A2(net378),
    .B1(net366),
    .B2(net2859),
    .X(_01054_));
 sky130_fd_sc_hd__a22o_1 _12154_ (.A1(net2859),
    .A2(net378),
    .B1(net366),
    .B2(net2863),
    .X(_01055_));
 sky130_fd_sc_hd__a22o_1 _12155_ (.A1(\genblk2.pcpi_div.quotient_msk[14] ),
    .A2(net378),
    .B1(net367),
    .B2(net2785),
    .X(_01056_));
 sky130_fd_sc_hd__a22o_1 _12156_ (.A1(\genblk2.pcpi_div.quotient_msk[15] ),
    .A2(net378),
    .B1(net367),
    .B2(net2776),
    .X(_01057_));
 sky130_fd_sc_hd__a22o_1 _12157_ (.A1(net2776),
    .A2(net378),
    .B1(net366),
    .B2(net2856),
    .X(_01058_));
 sky130_fd_sc_hd__a22o_1 _12158_ (.A1(net2856),
    .A2(net378),
    .B1(net365),
    .B2(net2893),
    .X(_01059_));
 sky130_fd_sc_hd__a22o_1 _12159_ (.A1(\genblk2.pcpi_div.quotient_msk[18] ),
    .A2(net377),
    .B1(net365),
    .B2(net2839),
    .X(_01060_));
 sky130_fd_sc_hd__a22o_1 _12160_ (.A1(\genblk2.pcpi_div.quotient_msk[19] ),
    .A2(net377),
    .B1(net365),
    .B2(net2794),
    .X(_01061_));
 sky130_fd_sc_hd__a22o_1 _12161_ (.A1(net2794),
    .A2(net384),
    .B1(net365),
    .B2(net2810),
    .X(_01062_));
 sky130_fd_sc_hd__a22o_1 _12162_ (.A1(net2810),
    .A2(net378),
    .B1(net365),
    .B2(net2828),
    .X(_01063_));
 sky130_fd_sc_hd__a22o_1 _12163_ (.A1(net2828),
    .A2(net378),
    .B1(net364),
    .B2(net2886),
    .X(_01064_));
 sky130_fd_sc_hd__a22o_1 _12164_ (.A1(\genblk2.pcpi_div.quotient_msk[23] ),
    .A2(net380),
    .B1(net369),
    .B2(net2867),
    .X(_01065_));
 sky130_fd_sc_hd__a22o_1 _12165_ (.A1(\genblk2.pcpi_div.quotient_msk[24] ),
    .A2(net380),
    .B1(net368),
    .B2(net2791),
    .X(_01066_));
 sky130_fd_sc_hd__a22o_1 _12166_ (.A1(net2791),
    .A2(net380),
    .B1(net368),
    .B2(net2882),
    .X(_01067_));
 sky130_fd_sc_hd__a22o_1 _12167_ (.A1(net2882),
    .A2(net380),
    .B1(net368),
    .B2(net2986),
    .X(_01068_));
 sky130_fd_sc_hd__a22o_1 _12168_ (.A1(\genblk2.pcpi_div.quotient_msk[27] ),
    .A2(net380),
    .B1(net368),
    .B2(net2843),
    .X(_01069_));
 sky130_fd_sc_hd__a22o_1 _12169_ (.A1(\genblk2.pcpi_div.quotient_msk[28] ),
    .A2(net380),
    .B1(net368),
    .B2(net2732),
    .X(_01070_));
 sky130_fd_sc_hd__a22o_1 _12170_ (.A1(net2732),
    .A2(net380),
    .B1(net368),
    .B2(net2847),
    .X(_01071_));
 sky130_fd_sc_hd__a22o_1 _12171_ (.A1(net2847),
    .A2(net380),
    .B1(net368),
    .B2(net2879),
    .X(_01072_));
 sky130_fd_sc_hd__o21ba_1 _12172_ (.A1(net2879),
    .A2(net750),
    .B1_N(net368),
    .X(_01073_));
 sky130_fd_sc_hd__a21oi_1 _12173_ (.A1(net2602),
    .A2(net277),
    .B1(net2746),
    .Y(_06579_));
 sky130_fd_sc_hd__nor2_1 _12174_ (.A(net751),
    .B(_06579_),
    .Y(_01074_));
 sky130_fd_sc_hd__a21oi_1 _12175_ (.A1(\genblk2.pcpi_div.quotient_msk[1] ),
    .A2(net277),
    .B1(net2999),
    .Y(_06580_));
 sky130_fd_sc_hd__nor2_1 _12176_ (.A(net751),
    .B(net3000),
    .Y(_01075_));
 sky130_fd_sc_hd__a21oi_1 _12177_ (.A1(net2750),
    .A2(net276),
    .B1(net2908),
    .Y(_06581_));
 sky130_fd_sc_hd__nor2_1 _12178_ (.A(net751),
    .B(_06581_),
    .Y(_01076_));
 sky130_fd_sc_hd__a21oi_1 _12179_ (.A1(\genblk2.pcpi_div.quotient_msk[3] ),
    .A2(net276),
    .B1(net2694),
    .Y(_06582_));
 sky130_fd_sc_hd__nor2_1 _12180_ (.A(net751),
    .B(net2695),
    .Y(_01077_));
 sky130_fd_sc_hd__a21oi_1 _12181_ (.A1(\genblk2.pcpi_div.quotient_msk[4] ),
    .A2(net276),
    .B1(net3011),
    .Y(_06583_));
 sky130_fd_sc_hd__nor2_1 _12182_ (.A(net751),
    .B(_06583_),
    .Y(_01078_));
 sky130_fd_sc_hd__a21oi_1 _12183_ (.A1(net2529),
    .A2(net276),
    .B1(net2925),
    .Y(_06584_));
 sky130_fd_sc_hd__nor2_1 _12184_ (.A(net751),
    .B(_06584_),
    .Y(_01079_));
 sky130_fd_sc_hd__a21oi_1 _12185_ (.A1(\genblk2.pcpi_div.quotient_msk[6] ),
    .A2(net276),
    .B1(net2685),
    .Y(_06585_));
 sky130_fd_sc_hd__nor2_1 _12186_ (.A(net751),
    .B(net2686),
    .Y(_01080_));
 sky130_fd_sc_hd__a21oi_1 _12187_ (.A1(net2909),
    .A2(net274),
    .B1(net2937),
    .Y(_06586_));
 sky130_fd_sc_hd__nor2_1 _12188_ (.A(net749),
    .B(_06586_),
    .Y(_01081_));
 sky130_fd_sc_hd__a21oi_1 _12189_ (.A1(\genblk2.pcpi_div.quotient_msk[8] ),
    .A2(net274),
    .B1(net2933),
    .Y(_06587_));
 sky130_fd_sc_hd__nor2_1 _12190_ (.A(net749),
    .B(net2934),
    .Y(_01082_));
 sky130_fd_sc_hd__a21oi_1 _12191_ (.A1(net2756),
    .A2(net274),
    .B1(net2877),
    .Y(_06588_));
 sky130_fd_sc_hd__nor2_1 _12192_ (.A(net749),
    .B(_06588_),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_1 _12193_ (.A1(net2798),
    .A2(net272),
    .B1(net2801),
    .Y(_06589_));
 sky130_fd_sc_hd__nor2_1 _12194_ (.A(net749),
    .B(_06589_),
    .Y(_01084_));
 sky130_fd_sc_hd__a21oi_1 _12195_ (.A1(\genblk2.pcpi_div.quotient_msk[11] ),
    .A2(net272),
    .B1(net2713),
    .Y(_06590_));
 sky130_fd_sc_hd__nor2_1 _12196_ (.A(net749),
    .B(net2714),
    .Y(_01085_));
 sky130_fd_sc_hd__a21oi_1 _12197_ (.A1(\genblk2.pcpi_div.quotient_msk[12] ),
    .A2(net271),
    .B1(net2961),
    .Y(_06591_));
 sky130_fd_sc_hd__nor2_1 _12198_ (.A(net748),
    .B(net2962),
    .Y(_01086_));
 sky130_fd_sc_hd__a21oi_1 _12199_ (.A1(\genblk2.pcpi_div.quotient_msk[13] ),
    .A2(net271),
    .B1(net2834),
    .Y(_06592_));
 sky130_fd_sc_hd__nor2_1 _12200_ (.A(net748),
    .B(net2835),
    .Y(_01087_));
 sky130_fd_sc_hd__a21oi_1 _12201_ (.A1(net2863),
    .A2(net274),
    .B1(net2944),
    .Y(_06593_));
 sky130_fd_sc_hd__nor2_1 _12202_ (.A(net749),
    .B(_06593_),
    .Y(_01088_));
 sky130_fd_sc_hd__a21oi_1 _12203_ (.A1(net2785),
    .A2(net272),
    .B1(net2829),
    .Y(_06594_));
 sky130_fd_sc_hd__nor2_1 _12204_ (.A(net748),
    .B(_06594_),
    .Y(_01089_));
 sky130_fd_sc_hd__a21oi_1 _12205_ (.A1(net2776),
    .A2(net270),
    .B1(net2819),
    .Y(_06595_));
 sky130_fd_sc_hd__nor2_1 _12206_ (.A(net748),
    .B(_06595_),
    .Y(_01090_));
 sky130_fd_sc_hd__a21oi_1 _12207_ (.A1(\genblk2.pcpi_div.quotient_msk[17] ),
    .A2(net269),
    .B1(net2735),
    .Y(_06596_));
 sky130_fd_sc_hd__nor2_1 _12208_ (.A(net748),
    .B(net2736),
    .Y(_01091_));
 sky130_fd_sc_hd__a21oi_1 _12209_ (.A1(net2893),
    .A2(net270),
    .B1(net2926),
    .Y(_06597_));
 sky130_fd_sc_hd__nor2_1 _12210_ (.A(net748),
    .B(_06597_),
    .Y(_01092_));
 sky130_fd_sc_hd__a21oi_1 _12211_ (.A1(\genblk2.pcpi_div.quotient_msk[19] ),
    .A2(net270),
    .B1(net2812),
    .Y(_06598_));
 sky130_fd_sc_hd__nor2_1 _12212_ (.A(net748),
    .B(net2813),
    .Y(_01093_));
 sky130_fd_sc_hd__a21oi_1 _12213_ (.A1(\genblk2.pcpi_div.quotient_msk[20] ),
    .A2(net270),
    .B1(net2761),
    .Y(_06599_));
 sky130_fd_sc_hd__nor2_1 _12214_ (.A(net748),
    .B(net2762),
    .Y(_01094_));
 sky130_fd_sc_hd__a21oi_1 _12215_ (.A1(net2810),
    .A2(net273),
    .B1(net2881),
    .Y(_06600_));
 sky130_fd_sc_hd__nor2_1 _12216_ (.A(net748),
    .B(_06600_),
    .Y(_01095_));
 sky130_fd_sc_hd__a21oi_1 _12217_ (.A1(\genblk2.pcpi_div.quotient_msk[22] ),
    .A2(net273),
    .B1(net2808),
    .Y(_06601_));
 sky130_fd_sc_hd__nor2_1 _12218_ (.A(net748),
    .B(net2809),
    .Y(_01096_));
 sky130_fd_sc_hd__a21oi_1 _12219_ (.A1(\genblk2.pcpi_div.quotient_msk[23] ),
    .A2(net273),
    .B1(net2766),
    .Y(_06602_));
 sky130_fd_sc_hd__nor2_1 _12220_ (.A(net749),
    .B(net2767),
    .Y(_01097_));
 sky130_fd_sc_hd__a21oi_1 _12221_ (.A1(\genblk2.pcpi_div.quotient_msk[24] ),
    .A2(net273),
    .B1(net2725),
    .Y(_06603_));
 sky130_fd_sc_hd__nor2_1 _12222_ (.A(net749),
    .B(net2726),
    .Y(_01098_));
 sky130_fd_sc_hd__a21oi_1 _12223_ (.A1(net2791),
    .A2(net273),
    .B1(net2820),
    .Y(_06604_));
 sky130_fd_sc_hd__nor2_1 _12224_ (.A(net750),
    .B(_06604_),
    .Y(_01099_));
 sky130_fd_sc_hd__a21oi_1 _12225_ (.A1(\genblk2.pcpi_div.quotient_msk[26] ),
    .A2(net275),
    .B1(net2595),
    .Y(_06605_));
 sky130_fd_sc_hd__nor2_1 _12226_ (.A(net750),
    .B(net2596),
    .Y(_01100_));
 sky130_fd_sc_hd__a21oi_1 _12227_ (.A1(net3072),
    .A2(net275),
    .B1(net2854),
    .Y(_06606_));
 sky130_fd_sc_hd__nor2_1 _12228_ (.A(net750),
    .B(_06606_),
    .Y(_01101_));
 sky130_fd_sc_hd__a21oi_1 _12229_ (.A1(\genblk2.pcpi_div.quotient_msk[28] ),
    .A2(net274),
    .B1(net2806),
    .Y(_06607_));
 sky130_fd_sc_hd__nor2_1 _12230_ (.A(net750),
    .B(net2807),
    .Y(_01102_));
 sky130_fd_sc_hd__a21oi_1 _12231_ (.A1(net2732),
    .A2(net274),
    .B1(net2985),
    .Y(_06608_));
 sky130_fd_sc_hd__nor2_1 _12232_ (.A(net750),
    .B(_06608_),
    .Y(_01103_));
 sky130_fd_sc_hd__a21oi_1 _12233_ (.A1(\genblk2.pcpi_div.quotient_msk[30] ),
    .A2(net275),
    .B1(net2753),
    .Y(_06609_));
 sky130_fd_sc_hd__nor2_1 _12234_ (.A(net750),
    .B(net2754),
    .Y(_01104_));
 sky130_fd_sc_hd__a21oi_1 _12235_ (.A1(\genblk2.pcpi_div.quotient_msk[31] ),
    .A2(net275),
    .B1(net2618),
    .Y(_06610_));
 sky130_fd_sc_hd__nor2_1 _12236_ (.A(net750),
    .B(net2619),
    .Y(_01105_));
 sky130_fd_sc_hd__a22o_1 _12237_ (.A1(net2579),
    .A2(net385),
    .B1(net371),
    .B2(\genblk2.pcpi_div.divisor[1] ),
    .X(_01106_));
 sky130_fd_sc_hd__a22o_1 _12238_ (.A1(\genblk2.pcpi_div.divisor[1] ),
    .A2(net385),
    .B1(net371),
    .B2(net2964),
    .X(_01107_));
 sky130_fd_sc_hd__a22o_1 _12239_ (.A1(\genblk2.pcpi_div.divisor[2] ),
    .A2(net385),
    .B1(net371),
    .B2(net2898),
    .X(_01108_));
 sky130_fd_sc_hd__a22o_1 _12240_ (.A1(\genblk2.pcpi_div.divisor[3] ),
    .A2(net383),
    .B1(net371),
    .B2(net2717),
    .X(_01109_));
 sky130_fd_sc_hd__a22o_1 _12241_ (.A1(net2717),
    .A2(net383),
    .B1(net372),
    .B2(net2734),
    .X(_01110_));
 sky130_fd_sc_hd__a22o_1 _12242_ (.A1(net2734),
    .A2(net382),
    .B1(net371),
    .B2(net2887),
    .X(_01111_));
 sky130_fd_sc_hd__a22o_1 _12243_ (.A1(\genblk2.pcpi_div.divisor[6] ),
    .A2(net382),
    .B1(net371),
    .B2(net2715),
    .X(_01112_));
 sky130_fd_sc_hd__a22o_1 _12244_ (.A1(net2715),
    .A2(net382),
    .B1(net366),
    .B2(\genblk2.pcpi_div.divisor[8] ),
    .X(_01113_));
 sky130_fd_sc_hd__a22o_1 _12245_ (.A1(\genblk2.pcpi_div.divisor[8] ),
    .A2(net379),
    .B1(net366),
    .B2(net2661),
    .X(_01114_));
 sky130_fd_sc_hd__a22o_1 _12246_ (.A1(net2661),
    .A2(net379),
    .B1(net366),
    .B2(net2742),
    .X(_01115_));
 sky130_fd_sc_hd__a22o_1 _12247_ (.A1(net2742),
    .A2(net379),
    .B1(net366),
    .B2(net2853),
    .X(_01116_));
 sky130_fd_sc_hd__a22o_1 _12248_ (.A1(\genblk2.pcpi_div.divisor[11] ),
    .A2(net379),
    .B1(net366),
    .B2(net2704),
    .X(_01117_));
 sky130_fd_sc_hd__a22o_1 _12249_ (.A1(\genblk2.pcpi_div.divisor[12] ),
    .A2(net379),
    .B1(net366),
    .B2(net2677),
    .X(_01118_));
 sky130_fd_sc_hd__a22o_1 _12250_ (.A1(net2677),
    .A2(net379),
    .B1(net364),
    .B2(net2728),
    .X(_01119_));
 sky130_fd_sc_hd__a22o_1 _12251_ (.A1(\genblk2.pcpi_div.divisor[14] ),
    .A2(net377),
    .B1(net364),
    .B2(net2657),
    .X(_01120_));
 sky130_fd_sc_hd__a22o_1 _12252_ (.A1(net2657),
    .A2(net377),
    .B1(net364),
    .B2(net2719),
    .X(_01121_));
 sky130_fd_sc_hd__a22o_1 _12253_ (.A1(net3069),
    .A2(net377),
    .B1(net364),
    .B2(net2702),
    .X(_01122_));
 sky130_fd_sc_hd__a22o_1 _12254_ (.A1(net2702),
    .A2(net377),
    .B1(net364),
    .B2(\genblk2.pcpi_div.divisor[18] ),
    .X(_01123_));
 sky130_fd_sc_hd__a22o_1 _12255_ (.A1(net2769),
    .A2(net377),
    .B1(net364),
    .B2(net2818),
    .X(_01124_));
 sky130_fd_sc_hd__a22o_1 _12256_ (.A1(net2818),
    .A2(net377),
    .B1(net364),
    .B2(\genblk2.pcpi_div.divisor[20] ),
    .X(_01125_));
 sky130_fd_sc_hd__a22o_1 _12257_ (.A1(\genblk2.pcpi_div.divisor[20] ),
    .A2(net377),
    .B1(net364),
    .B2(net2731),
    .X(_01126_));
 sky130_fd_sc_hd__a22o_1 _12258_ (.A1(net2731),
    .A2(net377),
    .B1(net364),
    .B2(net2816),
    .X(_01127_));
 sky130_fd_sc_hd__a22o_1 _12259_ (.A1(net2816),
    .A2(net381),
    .B1(net369),
    .B2(net2876),
    .X(_01128_));
 sky130_fd_sc_hd__a22o_1 _12260_ (.A1(\genblk2.pcpi_div.divisor[23] ),
    .A2(net381),
    .B1(net369),
    .B2(net2692),
    .X(_01129_));
 sky130_fd_sc_hd__a22o_1 _12261_ (.A1(net2692),
    .A2(net381),
    .B1(net369),
    .B2(net2775),
    .X(_01130_));
 sky130_fd_sc_hd__a22o_1 _12262_ (.A1(net2775),
    .A2(net381),
    .B1(net369),
    .B2(net2782),
    .X(_01131_));
 sky130_fd_sc_hd__a22o_1 _12263_ (.A1(\genblk2.pcpi_div.divisor[26] ),
    .A2(net381),
    .B1(net369),
    .B2(net2743),
    .X(_01132_));
 sky130_fd_sc_hd__a22o_1 _12264_ (.A1(net2743),
    .A2(net381),
    .B1(net369),
    .B2(net2903),
    .X(_01133_));
 sky130_fd_sc_hd__a22o_1 _12265_ (.A1(\genblk2.pcpi_div.divisor[28] ),
    .A2(net381),
    .B1(net369),
    .B2(net2873),
    .X(_01134_));
 sky130_fd_sc_hd__a22o_1 _12266_ (.A1(net2873),
    .A2(net380),
    .B1(net368),
    .B2(net2891),
    .X(_01135_));
 sky130_fd_sc_hd__a22o_1 _12267_ (.A1(\genblk2.pcpi_div.divisor[30] ),
    .A2(net380),
    .B1(net368),
    .B2(net2173),
    .X(_01136_));
 sky130_fd_sc_hd__nor2_1 _12268_ (.A(net1192),
    .B(_05096_),
    .Y(_01137_));
 sky130_fd_sc_hd__nor2_1 _12269_ (.A(net176),
    .B(_04298_),
    .Y(_06611_));
 sky130_fd_sc_hd__and3_1 _12270_ (.A(net175),
    .B(net174),
    .C(_06611_),
    .X(_01138_));
 sky130_fd_sc_hd__a31o_1 _12271_ (.A1(_02369_),
    .A2(_02448_),
    .A3(_06238_),
    .B1(_06252_),
    .X(_06612_));
 sky130_fd_sc_hd__a21o_1 _12272_ (.A1(net1234),
    .A2(net268),
    .B1(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__or4b_1 _12273_ (.A(mem_do_rdata),
    .B(mem_do_rinst),
    .C(\mem_state[1] ),
    .D_N(\mem_state[0] ),
    .X(_06614_));
 sky130_fd_sc_hd__a211o_1 _12274_ (.A1(_06250_),
    .A2(_06614_),
    .B1(_06612_),
    .C1(_06239_),
    .X(_06615_));
 sky130_fd_sc_hd__a21bo_1 _12275_ (.A1(net2760),
    .A2(_06613_),
    .B1_N(_06615_),
    .X(_01139_));
 sky130_fd_sc_hd__o21bai_1 _12276_ (.A1(_06239_),
    .A2(_06614_),
    .B1_N(net730),
    .Y(_06616_));
 sky130_fd_sc_hd__mux2_1 _12277_ (.A0(_06616_),
    .A1(net2960),
    .S(_06613_),
    .X(_01140_));
 sky130_fd_sc_hd__and3b_1 _12278_ (.A_N(net175),
    .B(net174),
    .C(_04299_),
    .X(_01141_));
 sky130_fd_sc_hd__and3b_1 _12279_ (.A_N(net174),
    .B(_04299_),
    .C(net175),
    .X(_01142_));
 sky130_fd_sc_hd__or2_1 _12280_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(is_sb_sh_sw),
    .X(_06617_));
 sky130_fd_sc_hd__or2_1 _12281_ (.A(_06223_),
    .B(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__a22o_1 _12282_ (.A1(net1150),
    .A2(net1128),
    .B1(_06618_),
    .B2(\mem_rdata_q[31] ),
    .X(_06619_));
 sky130_fd_sc_hd__and2_1 _12283_ (.A(net745),
    .B(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__and2_1 _12284_ (.A(\decoded_imm[31] ),
    .B(net739),
    .X(_06621_));
 sky130_fd_sc_hd__and2_1 _12285_ (.A(_02428_),
    .B(net745),
    .X(_06622_));
 sky130_fd_sc_hd__a211o_1 _12286_ (.A1(\mem_rdata_q[31] ),
    .A2(net559),
    .B1(_06621_),
    .C1(net532),
    .X(_01143_));
 sky130_fd_sc_hd__a221o_1 _12287_ (.A1(\decoded_imm[30] ),
    .A2(net739),
    .B1(net559),
    .B2(\mem_rdata_q[30] ),
    .C1(net532),
    .X(_01144_));
 sky130_fd_sc_hd__and2_1 _12288_ (.A(\decoded_imm[29] ),
    .B(net739),
    .X(_06623_));
 sky130_fd_sc_hd__a211o_1 _12289_ (.A1(\mem_rdata_q[29] ),
    .A2(_06622_),
    .B1(_06623_),
    .C1(_06620_),
    .X(_01145_));
 sky130_fd_sc_hd__and2_1 _12290_ (.A(\decoded_imm[28] ),
    .B(net739),
    .X(_06624_));
 sky130_fd_sc_hd__a211o_1 _12291_ (.A1(\mem_rdata_q[28] ),
    .A2(_06622_),
    .B1(_06624_),
    .C1(_06620_),
    .X(_01146_));
 sky130_fd_sc_hd__and2_1 _12292_ (.A(\decoded_imm[27] ),
    .B(net733),
    .X(_06625_));
 sky130_fd_sc_hd__a211o_1 _12293_ (.A1(\mem_rdata_q[27] ),
    .A2(net559),
    .B1(_06625_),
    .C1(net532),
    .X(_01147_));
 sky130_fd_sc_hd__and2_1 _12294_ (.A(\decoded_imm[26] ),
    .B(net733),
    .X(_06626_));
 sky130_fd_sc_hd__a211o_1 _12295_ (.A1(\mem_rdata_q[26] ),
    .A2(net559),
    .B1(_06626_),
    .C1(net532),
    .X(_01148_));
 sky130_fd_sc_hd__and2_1 _12296_ (.A(\decoded_imm[25] ),
    .B(net733),
    .X(_06627_));
 sky130_fd_sc_hd__a211o_1 _12297_ (.A1(\mem_rdata_q[25] ),
    .A2(net559),
    .B1(_06627_),
    .C1(net532),
    .X(_01149_));
 sky130_fd_sc_hd__and2_1 _12298_ (.A(\decoded_imm[24] ),
    .B(net733),
    .X(_06628_));
 sky130_fd_sc_hd__a211o_1 _12299_ (.A1(\mem_rdata_q[24] ),
    .A2(net559),
    .B1(_06628_),
    .C1(net532),
    .X(_01150_));
 sky130_fd_sc_hd__and2_1 _12300_ (.A(\decoded_imm[23] ),
    .B(net733),
    .X(_06629_));
 sky130_fd_sc_hd__a211o_1 _12301_ (.A1(\mem_rdata_q[23] ),
    .A2(net559),
    .B1(_06629_),
    .C1(net532),
    .X(_01151_));
 sky130_fd_sc_hd__and2_1 _12302_ (.A(\decoded_imm[22] ),
    .B(net733),
    .X(_06630_));
 sky130_fd_sc_hd__a211o_1 _12303_ (.A1(\mem_rdata_q[22] ),
    .A2(net559),
    .B1(_06630_),
    .C1(net532),
    .X(_01152_));
 sky130_fd_sc_hd__and2_1 _12304_ (.A(\decoded_imm[21] ),
    .B(net733),
    .X(_06631_));
 sky130_fd_sc_hd__a211o_1 _12305_ (.A1(\mem_rdata_q[21] ),
    .A2(net559),
    .B1(_06631_),
    .C1(net532),
    .X(_01153_));
 sky130_fd_sc_hd__a221o_1 _12306_ (.A1(\decoded_imm[20] ),
    .A2(net733),
    .B1(net559),
    .B2(\mem_rdata_q[20] ),
    .C1(net532),
    .X(_01154_));
 sky130_fd_sc_hd__a21o_2 _12307_ (.A1(\mem_rdata_q[31] ),
    .A2(_06618_),
    .B1(net733),
    .X(_06632_));
 sky130_fd_sc_hd__a22o_1 _12308_ (.A1(net1146),
    .A2(\decoded_imm_j[19] ),
    .B1(net970),
    .B2(\mem_rdata_q[19] ),
    .X(_06633_));
 sky130_fd_sc_hd__o22a_1 _12309_ (.A1(net3056),
    .A2(net743),
    .B1(_06632_),
    .B2(_06633_),
    .X(_01155_));
 sky130_fd_sc_hd__a22o_1 _12310_ (.A1(net1146),
    .A2(\decoded_imm_j[18] ),
    .B1(net970),
    .B2(\mem_rdata_q[18] ),
    .X(_06634_));
 sky130_fd_sc_hd__o22a_1 _12311_ (.A1(\decoded_imm[18] ),
    .A2(net743),
    .B1(_06632_),
    .B2(_06634_),
    .X(_01156_));
 sky130_fd_sc_hd__a22o_1 _12312_ (.A1(net1147),
    .A2(\decoded_imm_j[17] ),
    .B1(net970),
    .B2(\mem_rdata_q[17] ),
    .X(_06635_));
 sky130_fd_sc_hd__o22a_1 _12313_ (.A1(\decoded_imm[17] ),
    .A2(net743),
    .B1(_06632_),
    .B2(_06635_),
    .X(_01157_));
 sky130_fd_sc_hd__a22o_1 _12314_ (.A1(net1146),
    .A2(\decoded_imm_j[16] ),
    .B1(net970),
    .B2(\mem_rdata_q[16] ),
    .X(_06636_));
 sky130_fd_sc_hd__o22a_1 _12315_ (.A1(net3055),
    .A2(net743),
    .B1(_06632_),
    .B2(_06636_),
    .X(_01158_));
 sky130_fd_sc_hd__a22o_1 _12316_ (.A1(net1146),
    .A2(\decoded_imm_j[15] ),
    .B1(net970),
    .B2(\mem_rdata_q[15] ),
    .X(_06637_));
 sky130_fd_sc_hd__o22a_1 _12317_ (.A1(net3063),
    .A2(net743),
    .B1(_06632_),
    .B2(_06637_),
    .X(_01159_));
 sky130_fd_sc_hd__a22o_1 _12318_ (.A1(net1146),
    .A2(\decoded_imm_j[14] ),
    .B1(net970),
    .B2(\mem_rdata_q[14] ),
    .X(_06638_));
 sky130_fd_sc_hd__o22a_1 _12319_ (.A1(\decoded_imm[14] ),
    .A2(net743),
    .B1(_06632_),
    .B2(_06638_),
    .X(_01160_));
 sky130_fd_sc_hd__a22o_1 _12320_ (.A1(net1147),
    .A2(\decoded_imm_j[13] ),
    .B1(net970),
    .B2(\mem_rdata_q[13] ),
    .X(_06639_));
 sky130_fd_sc_hd__o22a_1 _12321_ (.A1(\decoded_imm[13] ),
    .A2(net743),
    .B1(_06632_),
    .B2(_06639_),
    .X(_01161_));
 sky130_fd_sc_hd__a22o_1 _12322_ (.A1(net1147),
    .A2(\decoded_imm_j[12] ),
    .B1(net970),
    .B2(\mem_rdata_q[12] ),
    .X(_06640_));
 sky130_fd_sc_hd__o22a_1 _12323_ (.A1(\decoded_imm[12] ),
    .A2(net743),
    .B1(_06632_),
    .B2(_06640_),
    .X(_01162_));
 sky130_fd_sc_hd__o21a_1 _12324_ (.A1(is_sb_sh_sw),
    .A2(_06223_),
    .B1(\mem_rdata_q[31] ),
    .X(_06641_));
 sky130_fd_sc_hd__a221o_1 _12325_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(\mem_rdata_q[7] ),
    .B1(\decoded_imm_j[11] ),
    .B2(net1151),
    .C1(net734),
    .X(_06642_));
 sky130_fd_sc_hd__o22a_1 _12326_ (.A1(\decoded_imm[11] ),
    .A2(net745),
    .B1(_06641_),
    .B2(_06642_),
    .X(_01163_));
 sky130_fd_sc_hd__and2_1 _12327_ (.A(net744),
    .B(_06618_),
    .X(_06643_));
 sky130_fd_sc_hd__and3_1 _12328_ (.A(net1148),
    .B(\decoded_imm_j[10] ),
    .C(net743),
    .X(_06644_));
 sky130_fd_sc_hd__a221o_1 _12329_ (.A1(\decoded_imm[10] ),
    .A2(net735),
    .B1(_06643_),
    .B2(\mem_rdata_q[30] ),
    .C1(_06644_),
    .X(_01164_));
 sky130_fd_sc_hd__and3_1 _12330_ (.A(net1148),
    .B(\decoded_imm_j[9] ),
    .C(net744),
    .X(_06645_));
 sky130_fd_sc_hd__a221o_1 _12331_ (.A1(\decoded_imm[9] ),
    .A2(net735),
    .B1(_06643_),
    .B2(\mem_rdata_q[29] ),
    .C1(_06645_),
    .X(_01165_));
 sky130_fd_sc_hd__and3_1 _12332_ (.A(net1148),
    .B(\decoded_imm_j[8] ),
    .C(net744),
    .X(_06646_));
 sky130_fd_sc_hd__a221o_1 _12333_ (.A1(\decoded_imm[8] ),
    .A2(net735),
    .B1(_06643_),
    .B2(\mem_rdata_q[28] ),
    .C1(_06646_),
    .X(_01166_));
 sky130_fd_sc_hd__and3_1 _12334_ (.A(net1148),
    .B(\decoded_imm_j[7] ),
    .C(net744),
    .X(_06647_));
 sky130_fd_sc_hd__a221o_1 _12335_ (.A1(\decoded_imm[7] ),
    .A2(net735),
    .B1(_06643_),
    .B2(\mem_rdata_q[27] ),
    .C1(_06647_),
    .X(_01167_));
 sky130_fd_sc_hd__and3_1 _12336_ (.A(net1148),
    .B(\decoded_imm_j[6] ),
    .C(net744),
    .X(_06648_));
 sky130_fd_sc_hd__a221o_1 _12337_ (.A1(\decoded_imm[6] ),
    .A2(net735),
    .B1(_06643_),
    .B2(\mem_rdata_q[26] ),
    .C1(_06648_),
    .X(_01168_));
 sky130_fd_sc_hd__and3_1 _12338_ (.A(net1148),
    .B(\decoded_imm_j[5] ),
    .C(net743),
    .X(_06649_));
 sky130_fd_sc_hd__a221o_1 _12339_ (.A1(\decoded_imm[5] ),
    .A2(net735),
    .B1(_06643_),
    .B2(\mem_rdata_q[25] ),
    .C1(_06649_),
    .X(_01169_));
 sky130_fd_sc_hd__and2_1 _12340_ (.A(\mem_rdata_q[24] ),
    .B(_06223_),
    .X(_06650_));
 sky130_fd_sc_hd__a221o_1 _12341_ (.A1(net1151),
    .A2(\decoded_imm_j[4] ),
    .B1(_06617_),
    .B2(\mem_rdata_q[11] ),
    .C1(net734),
    .X(_06651_));
 sky130_fd_sc_hd__o22a_1 _12342_ (.A1(\decoded_imm[4] ),
    .A2(net745),
    .B1(_06650_),
    .B2(_06651_),
    .X(_01170_));
 sky130_fd_sc_hd__and2_1 _12343_ (.A(\mem_rdata_q[23] ),
    .B(_06223_),
    .X(_06652_));
 sky130_fd_sc_hd__a221o_1 _12344_ (.A1(net1151),
    .A2(\decoded_imm_j[3] ),
    .B1(_06617_),
    .B2(\mem_rdata_q[10] ),
    .C1(net734),
    .X(_06653_));
 sky130_fd_sc_hd__o22a_1 _12345_ (.A1(\decoded_imm[3] ),
    .A2(net745),
    .B1(_06652_),
    .B2(_06653_),
    .X(_01171_));
 sky130_fd_sc_hd__and2_1 _12346_ (.A(\mem_rdata_q[22] ),
    .B(_06223_),
    .X(_06654_));
 sky130_fd_sc_hd__a221o_1 _12347_ (.A1(net1151),
    .A2(\decoded_imm_j[2] ),
    .B1(_06617_),
    .B2(\mem_rdata_q[9] ),
    .C1(net733),
    .X(_06655_));
 sky130_fd_sc_hd__o22a_1 _12348_ (.A1(net3019),
    .A2(net745),
    .B1(_06654_),
    .B2(_06655_),
    .X(_01172_));
 sky130_fd_sc_hd__and2_1 _12349_ (.A(\mem_rdata_q[8] ),
    .B(_06617_),
    .X(_06656_));
 sky130_fd_sc_hd__a221o_1 _12350_ (.A1(net1151),
    .A2(\decoded_imm_j[1] ),
    .B1(_06223_),
    .B2(\mem_rdata_q[21] ),
    .C1(net734),
    .X(_06657_));
 sky130_fd_sc_hd__o22a_1 _12351_ (.A1(\decoded_imm[1] ),
    .A2(net745),
    .B1(_06656_),
    .B2(_06657_),
    .X(_01173_));
 sky130_fd_sc_hd__or4_1 _12352_ (.A(\genblk1.genblk1.pcpi_mul.mul_counter[0] ),
    .B(\genblk1.genblk1.pcpi_mul.mul_counter[3] ),
    .C(\genblk1.genblk1.pcpi_mul.mul_counter[2] ),
    .D(\genblk1.genblk1.pcpi_mul.mul_counter[1] ),
    .X(_06658_));
 sky130_fd_sc_hd__or3_1 _12353_ (.A(\genblk1.genblk1.pcpi_mul.mul_counter[4] ),
    .B(_02415_),
    .C(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__o21ai_1 _12354_ (.A1(\genblk1.genblk1.pcpi_mul.mul_counter[4] ),
    .A2(_06658_),
    .B1(_02415_),
    .Y(_06660_));
 sky130_fd_sc_hd__a22o_1 _12355_ (.A1(net1218),
    .A2(\genblk1.genblk1.pcpi_mul.mul_counter[5] ),
    .B1(net956),
    .B2(net917),
    .X(_06661_));
 sky130_fd_sc_hd__a31o_1 _12356_ (.A1(net910),
    .A2(_06659_),
    .A3(_06660_),
    .B1(_06661_),
    .X(_01174_));
 sky130_fd_sc_hd__and3b_1 _12357_ (.A_N(\latched_rd[0] ),
    .B(_04290_),
    .C(\latched_rd[1] ),
    .X(_06662_));
 sky130_fd_sc_hd__mux2_1 _12358_ (.A0(net1873),
    .A1(net586),
    .S(net362),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _12359_ (.A0(net1636),
    .A1(net584),
    .S(net362),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _12360_ (.A0(net1387),
    .A1(net582),
    .S(net362),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _12361_ (.A0(net1376),
    .A1(net578),
    .S(net361),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _12362_ (.A0(net1377),
    .A1(net573),
    .S(net361),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(net1372),
    .A1(net543),
    .S(net361),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(net1411),
    .A1(net540),
    .S(net361),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _12365_ (.A0(net1522),
    .A1(net525),
    .S(net360),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _12366_ (.A0(net1547),
    .A1(net522),
    .S(net360),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _12367_ (.A0(net1362),
    .A1(net409),
    .S(net360),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(net1627),
    .A1(net405),
    .S(net360),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _12369_ (.A0(net1849),
    .A1(net355),
    .S(net360),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _12370_ (.A0(net1340),
    .A1(net351),
    .S(net360),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _12371_ (.A0(net1446),
    .A1(net348),
    .S(net360),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(net1441),
    .A1(net345),
    .S(net361),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _12373_ (.A0(net1383),
    .A1(net340),
    .S(net360),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(net1452),
    .A1(_03810_),
    .S(net361),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _12375_ (.A0(net1388),
    .A1(net332),
    .S(net360),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(net1391),
    .A1(net328),
    .S(net360),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _12377_ (.A0(net1809),
    .A1(net325),
    .S(net362),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(net1342),
    .A1(net322),
    .S(net361),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _12379_ (.A0(net1645),
    .A1(net316),
    .S(net361),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(net2122),
    .A1(net313),
    .S(net362),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _12381_ (.A0(net1432),
    .A1(net310),
    .S(net362),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(net1423),
    .A1(net307),
    .S(net362),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _12383_ (.A0(net1341),
    .A1(net303),
    .S(net362),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(net1571),
    .A1(net300),
    .S(net362),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _12385_ (.A0(net1457),
    .A1(net295),
    .S(net363),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(net1487),
    .A1(net291),
    .S(net363),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _12387_ (.A0(net1403),
    .A1(net288),
    .S(net362),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(net1597),
    .A1(net282),
    .S(net363),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _12389_ (.A0(net1418),
    .A1(net280),
    .S(net363),
    .X(_01206_));
 sky130_fd_sc_hd__or3b_1 _12390_ (.A(\latched_rd[4] ),
    .B(\latched_rd[3] ),
    .C_N(\latched_rd[2] ),
    .X(_06663_));
 sky130_fd_sc_hd__or2_2 _12391_ (.A(_04273_),
    .B(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__mux2_1 _12392_ (.A0(net588),
    .A1(net1990),
    .S(net474),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(_03751_),
    .A1(net2063),
    .S(net473),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(net579),
    .A1(net1828),
    .S(net473),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(net575),
    .A1(net2046),
    .S(net472),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _12396_ (.A0(net571),
    .A1(net2032),
    .S(net472),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _12397_ (.A0(net541),
    .A1(net1942),
    .S(net472),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(net538),
    .A1(net1717),
    .S(net472),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(net527),
    .A1(net1866),
    .S(net471),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _12400_ (.A0(net522),
    .A1(net2135),
    .S(net471),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _12401_ (.A0(net408),
    .A1(net2015),
    .S(net472),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(net403),
    .A1(net2043),
    .S(net471),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(net356),
    .A1(net2123),
    .S(net471),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _12404_ (.A0(net352),
    .A1(net1879),
    .S(net471),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _12405_ (.A0(_03799_),
    .A1(net1727),
    .S(net471),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _12406_ (.A0(_03802_),
    .A1(net2000),
    .S(net471),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(net342),
    .A1(net1954),
    .S(net471),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _12408_ (.A0(net338),
    .A1(net1756),
    .S(net472),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(net335),
    .A1(net1977),
    .S(net471),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(net330),
    .A1(net2218),
    .S(net471),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _12411_ (.A0(net326),
    .A1(net1891),
    .S(net474),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(net323),
    .A1(net1738),
    .S(net472),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _12413_ (.A0(net317),
    .A1(net1919),
    .S(net474),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(net314),
    .A1(net2166),
    .S(net473),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _12415_ (.A0(net309),
    .A1(net1986),
    .S(net472),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _12416_ (.A0(net306),
    .A1(net2363),
    .S(net473),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(net301),
    .A1(net1939),
    .S(net474),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(net297),
    .A1(net1516),
    .S(net473),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(net293),
    .A1(net2039),
    .S(net473),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _12420_ (.A0(net291),
    .A1(net1966),
    .S(net473),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _12421_ (.A0(net285),
    .A1(net1590),
    .S(net473),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _12422_ (.A0(net284),
    .A1(net1999),
    .S(net473),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _12423_ (.A0(net279),
    .A1(net2010),
    .S(net473),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(net910),
    .A1(net1217),
    .S(net2990),
    .X(_01239_));
 sky130_fd_sc_hd__o21a_1 _12425_ (.A1(net1218),
    .A2(\genblk1.genblk1.pcpi_mul.mul_counter[0] ),
    .B1(net3012),
    .X(_06665_));
 sky130_fd_sc_hd__or3_1 _12426_ (.A(net1218),
    .B(\genblk1.genblk1.pcpi_mul.mul_counter[0] ),
    .C(\genblk1.genblk1.pcpi_mul.mul_counter[1] ),
    .X(_06666_));
 sky130_fd_sc_hd__or3b_1 _12427_ (.A(net917),
    .B(_06665_),
    .C_N(_06666_),
    .X(_01240_));
 sky130_fd_sc_hd__a21oi_1 _12428_ (.A1(net2709),
    .A2(_06666_),
    .B1(net917),
    .Y(_06667_));
 sky130_fd_sc_hd__o21ai_1 _12429_ (.A1(net2709),
    .A2(_06666_),
    .B1(_06667_),
    .Y(_01241_));
 sky130_fd_sc_hd__o21a_1 _12430_ (.A1(\genblk1.genblk1.pcpi_mul.mul_counter[2] ),
    .A2(_06666_),
    .B1(\genblk1.genblk1.pcpi_mul.mul_counter[3] ),
    .X(_06668_));
 sky130_fd_sc_hd__or3_1 _12431_ (.A(\genblk1.genblk1.pcpi_mul.mul_counter[3] ),
    .B(\genblk1.genblk1.pcpi_mul.mul_counter[2] ),
    .C(_06666_),
    .X(_06669_));
 sky130_fd_sc_hd__or3b_1 _12432_ (.A(net917),
    .B(_06668_),
    .C_N(_06669_),
    .X(_01242_));
 sky130_fd_sc_hd__or2_1 _12433_ (.A(\genblk1.genblk1.pcpi_mul.mul_counter[4] ),
    .B(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__a21oi_1 _12434_ (.A1(net2811),
    .A2(_06669_),
    .B1(net917),
    .Y(_06671_));
 sky130_fd_sc_hd__nand2_1 _12435_ (.A(_06670_),
    .B(_06671_),
    .Y(_01243_));
 sky130_fd_sc_hd__mux2_1 _12436_ (.A0(net1180),
    .A1(\genblk2.pcpi_div.divisor[32] ),
    .S(net865),
    .X(_06672_));
 sky130_fd_sc_hd__mux2_1 _12437_ (.A0(_06672_),
    .A1(net2173),
    .S(net384),
    .X(_01244_));
 sky130_fd_sc_hd__and2_1 _12438_ (.A(net1157),
    .B(_02507_),
    .X(_06673_));
 sky130_fd_sc_hd__nand2_1 _12439_ (.A(net1157),
    .B(_02507_),
    .Y(_06674_));
 sky130_fd_sc_hd__nand2_1 _12440_ (.A(net1180),
    .B(net717),
    .Y(_06675_));
 sky130_fd_sc_hd__xnor2_1 _12441_ (.A(net1178),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__mux2_1 _12442_ (.A0(\genblk2.pcpi_div.divisor[33] ),
    .A1(_06676_),
    .S(net868),
    .X(_06677_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(_06677_),
    .A1(net2771),
    .S(net383),
    .X(_01245_));
 sky130_fd_sc_hd__o21ai_1 _12444_ (.A1(net1180),
    .A2(net1178),
    .B1(net717),
    .Y(_06678_));
 sky130_fd_sc_hd__xnor2_1 _12445_ (.A(net1177),
    .B(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__mux2_1 _12446_ (.A0(\genblk2.pcpi_div.divisor[34] ),
    .A1(_06679_),
    .S(net868),
    .X(_06680_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(_06680_),
    .A1(net2552),
    .S(net383),
    .X(_01246_));
 sky130_fd_sc_hd__o31a_1 _12448_ (.A1(net1180),
    .A2(net1179),
    .A3(net1177),
    .B1(net717),
    .X(_06681_));
 sky130_fd_sc_hd__xnor2_1 _12449_ (.A(_02392_),
    .B(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__mux2_1 _12450_ (.A0(\genblk2.pcpi_div.divisor[35] ),
    .A1(_06682_),
    .S(net868),
    .X(_06683_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(_06683_),
    .A1(net2570),
    .S(net383),
    .X(_01247_));
 sky130_fd_sc_hd__a21oi_1 _12452_ (.A1(_05098_),
    .A2(net717),
    .B1(net1174),
    .Y(_06684_));
 sky130_fd_sc_hd__a31o_1 _12453_ (.A1(net1174),
    .A2(_05098_),
    .A3(net717),
    .B1(net865),
    .X(_06685_));
 sky130_fd_sc_hd__a2bb2o_1 _12454_ (.A1_N(_06684_),
    .A2_N(_06685_),
    .B1(\genblk2.pcpi_div.divisor[36] ),
    .B2(net865),
    .X(_06686_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(_06686_),
    .A1(net2545),
    .S(net383),
    .X(_01248_));
 sky130_fd_sc_hd__a21oi_1 _12456_ (.A1(_05099_),
    .A2(net717),
    .B1(net1172),
    .Y(_06687_));
 sky130_fd_sc_hd__a31o_1 _12457_ (.A1(net1172),
    .A2(_05099_),
    .A3(net717),
    .B1(net865),
    .X(_06688_));
 sky130_fd_sc_hd__a2bb2o_1 _12458_ (.A1_N(_06687_),
    .A2_N(_06688_),
    .B1(\genblk2.pcpi_div.divisor[37] ),
    .B2(net865),
    .X(_06689_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(_06689_),
    .A1(net2551),
    .S(net383),
    .X(_01249_));
 sky130_fd_sc_hd__o31a_1 _12460_ (.A1(net1172),
    .A2(net1175),
    .A3(_05098_),
    .B1(net717),
    .X(_06690_));
 sky130_fd_sc_hd__xor2_1 _12461_ (.A(net1171),
    .B(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(\genblk2.pcpi_div.divisor[38] ),
    .A1(_06691_),
    .S(net869),
    .X(_06692_));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(_06692_),
    .A1(net2546),
    .S(net383),
    .X(_01250_));
 sky130_fd_sc_hd__nand2_1 _12464_ (.A(_05100_),
    .B(net717),
    .Y(_06693_));
 sky130_fd_sc_hd__xnor2_1 _12465_ (.A(net1169),
    .B(_06693_),
    .Y(_06694_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(\genblk2.pcpi_div.divisor[39] ),
    .A1(_06694_),
    .S(net868),
    .X(_06695_));
 sky130_fd_sc_hd__mux2_1 _12467_ (.A0(_06695_),
    .A1(net2571),
    .S(net384),
    .X(_01251_));
 sky130_fd_sc_hd__o21ai_1 _12468_ (.A1(net1169),
    .A2(_05100_),
    .B1(net718),
    .Y(_06696_));
 sky130_fd_sc_hd__xnor2_1 _12469_ (.A(net1168),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(\genblk2.pcpi_div.divisor[40] ),
    .A1(_06697_),
    .S(net868),
    .X(_06698_));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(_06698_),
    .A1(net2566),
    .S(net386),
    .X(_01252_));
 sky130_fd_sc_hd__or3b_1 _12472_ (.A(net1167),
    .B(net715),
    .C_N(_05101_),
    .X(_06699_));
 sky130_fd_sc_hd__a21bo_1 _12473_ (.A1(_05101_),
    .A2(net717),
    .B1_N(net1167),
    .X(_06700_));
 sky130_fd_sc_hd__or2_1 _12474_ (.A(net2533),
    .B(net868),
    .X(_06701_));
 sky130_fd_sc_hd__a31oi_1 _12475_ (.A1(net868),
    .A2(_06699_),
    .A3(_06700_),
    .B1(net386),
    .Y(_06702_));
 sky130_fd_sc_hd__a22o_1 _12476_ (.A1(net2599),
    .A2(net386),
    .B1(_06701_),
    .B2(_06702_),
    .X(_01253_));
 sky130_fd_sc_hd__or3b_1 _12477_ (.A(net1166),
    .B(net715),
    .C_N(_05102_),
    .X(_06703_));
 sky130_fd_sc_hd__a21bo_1 _12478_ (.A1(_05102_),
    .A2(net718),
    .B1_N(net1166),
    .X(_06704_));
 sky130_fd_sc_hd__nor2_1 _12479_ (.A(\genblk2.pcpi_div.divisor[42] ),
    .B(net870),
    .Y(_06705_));
 sky130_fd_sc_hd__a31o_1 _12480_ (.A1(net870),
    .A2(_06703_),
    .A3(_06704_),
    .B1(net386),
    .X(_06706_));
 sky130_fd_sc_hd__a2bb2o_1 _12481_ (.A1_N(_06705_),
    .A2_N(_06706_),
    .B1(net2533),
    .B2(net386),
    .X(_01254_));
 sky130_fd_sc_hd__or3_1 _12482_ (.A(net1165),
    .B(_05103_),
    .C(net715),
    .X(_06707_));
 sky130_fd_sc_hd__o21ai_1 _12483_ (.A1(_05103_),
    .A2(net715),
    .B1(net1165),
    .Y(_06708_));
 sky130_fd_sc_hd__nor2_1 _12484_ (.A(\genblk2.pcpi_div.divisor[43] ),
    .B(net870),
    .Y(_06709_));
 sky130_fd_sc_hd__a31o_1 _12485_ (.A1(net870),
    .A2(_06707_),
    .A3(_06708_),
    .B1(net386),
    .X(_06710_));
 sky130_fd_sc_hd__a2bb2o_1 _12486_ (.A1_N(_06709_),
    .A2_N(_06710_),
    .B1(net2687),
    .B2(net386),
    .X(_01255_));
 sky130_fd_sc_hd__or3b_1 _12487_ (.A(net1164),
    .B(net715),
    .C_N(_05104_),
    .X(_06711_));
 sky130_fd_sc_hd__a21bo_1 _12488_ (.A1(_05104_),
    .A2(net718),
    .B1_N(net1164),
    .X(_06712_));
 sky130_fd_sc_hd__or2_1 _12489_ (.A(net2536),
    .B(net871),
    .X(_06713_));
 sky130_fd_sc_hd__a31oi_1 _12490_ (.A1(net871),
    .A2(_06711_),
    .A3(_06712_),
    .B1(net386),
    .Y(_06714_));
 sky130_fd_sc_hd__a22o_1 _12491_ (.A1(net2669),
    .A2(net386),
    .B1(_06713_),
    .B2(_06714_),
    .X(_01256_));
 sky130_fd_sc_hd__or3b_1 _12492_ (.A(net1163),
    .B(net715),
    .C_N(_05105_),
    .X(_06715_));
 sky130_fd_sc_hd__a21bo_1 _12493_ (.A1(_05105_),
    .A2(net718),
    .B1_N(net1163),
    .X(_01990_));
 sky130_fd_sc_hd__nor2_1 _12494_ (.A(\genblk2.pcpi_div.divisor[45] ),
    .B(net871),
    .Y(_01991_));
 sky130_fd_sc_hd__a31o_1 _12495_ (.A1(net871),
    .A2(_06715_),
    .A3(_01990_),
    .B1(net387),
    .X(_01992_));
 sky130_fd_sc_hd__a2bb2o_1 _12496_ (.A1_N(_01991_),
    .A2_N(_01992_),
    .B1(net2536),
    .B2(net387),
    .X(_01257_));
 sky130_fd_sc_hd__or3_1 _12497_ (.A(net240),
    .B(_05106_),
    .C(net715),
    .X(_01993_));
 sky130_fd_sc_hd__o21ai_1 _12498_ (.A1(_05106_),
    .A2(net716),
    .B1(net240),
    .Y(_01994_));
 sky130_fd_sc_hd__nor2_1 _12499_ (.A(\genblk2.pcpi_div.divisor[46] ),
    .B(net870),
    .Y(_01995_));
 sky130_fd_sc_hd__a31o_1 _12500_ (.A1(net871),
    .A2(_01993_),
    .A3(_01994_),
    .B1(net387),
    .X(_01996_));
 sky130_fd_sc_hd__a2bb2o_1 _12501_ (.A1_N(_01995_),
    .A2_N(_01996_),
    .B1(net2623),
    .B2(net386),
    .X(_01258_));
 sky130_fd_sc_hd__or3b_1 _12502_ (.A(net1162),
    .B(net715),
    .C_N(_05107_),
    .X(_01997_));
 sky130_fd_sc_hd__a21bo_1 _12503_ (.A1(_05107_),
    .A2(net718),
    .B1_N(net241),
    .X(_01998_));
 sky130_fd_sc_hd__or2_1 _12504_ (.A(\genblk2.pcpi_div.divisor[47] ),
    .B(net870),
    .X(_01999_));
 sky130_fd_sc_hd__a31oi_1 _12505_ (.A1(net870),
    .A2(_01997_),
    .A3(_01998_),
    .B1(net387),
    .Y(_02000_));
 sky130_fd_sc_hd__a22o_1 _12506_ (.A1(net2666),
    .A2(net387),
    .B1(_01999_),
    .B2(_02000_),
    .X(_01259_));
 sky130_fd_sc_hd__a21oi_1 _12507_ (.A1(_05108_),
    .A2(net718),
    .B1(_02395_),
    .Y(_02001_));
 sky130_fd_sc_hd__a31o_1 _12508_ (.A1(_02395_),
    .A2(_05108_),
    .A3(net720),
    .B1(net866),
    .X(_02002_));
 sky130_fd_sc_hd__or2_1 _12509_ (.A(\genblk2.pcpi_div.divisor[48] ),
    .B(net870),
    .X(_02003_));
 sky130_fd_sc_hd__o21ba_1 _12510_ (.A1(_02001_),
    .A2(_02002_),
    .B1_N(net385),
    .X(_02004_));
 sky130_fd_sc_hd__a22o_1 _12511_ (.A1(net2543),
    .A2(net387),
    .B1(_02003_),
    .B2(_02004_),
    .X(_01260_));
 sky130_fd_sc_hd__o21ai_1 _12512_ (.A1(_05109_),
    .A2(net715),
    .B1(net1160),
    .Y(_02005_));
 sky130_fd_sc_hd__or3_1 _12513_ (.A(net1160),
    .B(_05109_),
    .C(net715),
    .X(_02006_));
 sky130_fd_sc_hd__nor2_1 _12514_ (.A(\genblk2.pcpi_div.divisor[49] ),
    .B(net870),
    .Y(_02007_));
 sky130_fd_sc_hd__a31o_1 _12515_ (.A1(net870),
    .A2(_02005_),
    .A3(_02006_),
    .B1(net385),
    .X(_02008_));
 sky130_fd_sc_hd__a2bb2o_1 _12516_ (.A1_N(_02007_),
    .A2_N(_02008_),
    .B1(net2563),
    .B2(net385),
    .X(_01261_));
 sky130_fd_sc_hd__or3b_1 _12517_ (.A(net244),
    .B(net716),
    .C_N(_05110_),
    .X(_02009_));
 sky130_fd_sc_hd__a21bo_1 _12518_ (.A1(_05110_),
    .A2(net718),
    .B1_N(net244),
    .X(_02010_));
 sky130_fd_sc_hd__or2_1 _12519_ (.A(\genblk2.pcpi_div.divisor[50] ),
    .B(net872),
    .X(_02011_));
 sky130_fd_sc_hd__a31oi_1 _12520_ (.A1(net871),
    .A2(_02009_),
    .A3(_02010_),
    .B1(net388),
    .Y(_02012_));
 sky130_fd_sc_hd__a22o_1 _12521_ (.A1(net2664),
    .A2(net385),
    .B1(_02011_),
    .B2(_02012_),
    .X(_01262_));
 sky130_fd_sc_hd__or3b_1 _12522_ (.A(net1159),
    .B(net716),
    .C_N(_05111_),
    .X(_02013_));
 sky130_fd_sc_hd__a21bo_1 _12523_ (.A1(_05111_),
    .A2(net718),
    .B1_N(net245),
    .X(_02014_));
 sky130_fd_sc_hd__nor2_1 _12524_ (.A(\genblk2.pcpi_div.divisor[51] ),
    .B(net872),
    .Y(_02015_));
 sky130_fd_sc_hd__a31o_1 _12525_ (.A1(net872),
    .A2(_02013_),
    .A3(_02014_),
    .B1(net388),
    .X(_02016_));
 sky130_fd_sc_hd__a2bb2o_1 _12526_ (.A1_N(_02015_),
    .A2_N(_02016_),
    .B1(net2600),
    .B2(net385),
    .X(_01263_));
 sky130_fd_sc_hd__o21a_1 _12527_ (.A1(net245),
    .A2(_05111_),
    .B1(net718),
    .X(_02017_));
 sky130_fd_sc_hd__xor2_1 _12528_ (.A(net247),
    .B(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _12529_ (.A0(\genblk2.pcpi_div.divisor[52] ),
    .A1(_02018_),
    .S(net872),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _12530_ (.A0(_02019_),
    .A1(net2653),
    .S(net385),
    .X(_01264_));
 sky130_fd_sc_hd__nand2_1 _12531_ (.A(_05112_),
    .B(net719),
    .Y(_02020_));
 sky130_fd_sc_hd__xnor2_1 _12532_ (.A(net248),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__mux2_1 _12533_ (.A0(\genblk2.pcpi_div.divisor[53] ),
    .A1(_02021_),
    .S(net872),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_1 _12534_ (.A0(_02022_),
    .A1(net2690),
    .S(net389),
    .X(_01265_));
 sky130_fd_sc_hd__nand2_1 _12535_ (.A(_05113_),
    .B(net719),
    .Y(_02023_));
 sky130_fd_sc_hd__xnor2_1 _12536_ (.A(net1158),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(\genblk2.pcpi_div.divisor[54] ),
    .A1(_02024_),
    .S(_05082_),
    .X(_02025_));
 sky130_fd_sc_hd__mux2_1 _12538_ (.A0(_02025_),
    .A1(net2534),
    .S(net389),
    .X(_01266_));
 sky130_fd_sc_hd__o21ai_1 _12539_ (.A1(net1158),
    .A2(_05113_),
    .B1(net719),
    .Y(_02026_));
 sky130_fd_sc_hd__xnor2_1 _12540_ (.A(net250),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\genblk2.pcpi_div.divisor[55] ),
    .A1(_02027_),
    .S(net874),
    .X(_02028_));
 sky130_fd_sc_hd__mux2_1 _12542_ (.A0(_02028_),
    .A1(net2581),
    .S(net389),
    .X(_01267_));
 sky130_fd_sc_hd__a21oi_1 _12543_ (.A1(_05114_),
    .A2(net719),
    .B1(_02396_),
    .Y(_02029_));
 sky130_fd_sc_hd__a31o_1 _12544_ (.A1(_02396_),
    .A2(_05114_),
    .A3(net719),
    .B1(net866),
    .X(_02030_));
 sky130_fd_sc_hd__o22a_1 _12545_ (.A1(\genblk2.pcpi_div.divisor[56] ),
    .A2(net874),
    .B1(_02029_),
    .B2(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(_02031_),
    .A1(net2722),
    .S(net390),
    .X(_01268_));
 sky130_fd_sc_hd__o21ai_1 _12547_ (.A1(net251),
    .A2(_05114_),
    .B1(net719),
    .Y(_02032_));
 sky130_fd_sc_hd__xnor2_1 _12548_ (.A(net252),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__mux2_1 _12549_ (.A0(\genblk2.pcpi_div.divisor[57] ),
    .A1(_02033_),
    .S(net874),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(_02034_),
    .A1(net2631),
    .S(net389),
    .X(_01269_));
 sky130_fd_sc_hd__nand2_1 _12551_ (.A(_05115_),
    .B(net719),
    .Y(_02035_));
 sky130_fd_sc_hd__xnor2_1 _12552_ (.A(net253),
    .B(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(\genblk2.pcpi_div.divisor[58] ),
    .A1(_02036_),
    .S(net874),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(_02037_),
    .A1(net2535),
    .S(net389),
    .X(_01270_));
 sky130_fd_sc_hd__or3b_1 _12555_ (.A(net254),
    .B(net716),
    .C_N(_05116_),
    .X(_02038_));
 sky130_fd_sc_hd__a21o_1 _12556_ (.A1(_05116_),
    .A2(net719),
    .B1(_02397_),
    .X(_02039_));
 sky130_fd_sc_hd__or2_1 _12557_ (.A(\genblk2.pcpi_div.divisor[59] ),
    .B(net874),
    .X(_02040_));
 sky130_fd_sc_hd__a31oi_1 _12558_ (.A1(net874),
    .A2(_02038_),
    .A3(_02039_),
    .B1(net389),
    .Y(_02041_));
 sky130_fd_sc_hd__a22o_1 _12559_ (.A1(net2553),
    .A2(net389),
    .B1(_02040_),
    .B2(_02041_),
    .X(_01271_));
 sky130_fd_sc_hd__a21oi_1 _12560_ (.A1(_05117_),
    .A2(net720),
    .B1(_02399_),
    .Y(_02042_));
 sky130_fd_sc_hd__a31o_1 _12561_ (.A1(_02399_),
    .A2(_05117_),
    .A3(net720),
    .B1(_05083_),
    .X(_02043_));
 sky130_fd_sc_hd__o22a_1 _12562_ (.A1(\genblk2.pcpi_div.divisor[60] ),
    .A2(net874),
    .B1(_02042_),
    .B2(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _12563_ (.A0(_02044_),
    .A1(net2627),
    .S(net390),
    .X(_01272_));
 sky130_fd_sc_hd__o21a_1 _12564_ (.A1(net255),
    .A2(_05117_),
    .B1(net719),
    .X(_02045_));
 sky130_fd_sc_hd__xnor2_1 _12565_ (.A(_02398_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(\genblk2.pcpi_div.divisor[61] ),
    .A1(_02046_),
    .S(net874),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _12567_ (.A0(_02047_),
    .A1(net2634),
    .S(net389),
    .X(_01273_));
 sky130_fd_sc_hd__nand2_1 _12568_ (.A(_05118_),
    .B(net719),
    .Y(_02048_));
 sky130_fd_sc_hd__xnor2_1 _12569_ (.A(net258),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__mux2_1 _12570_ (.A0(\genblk2.pcpi_div.divisor[62] ),
    .A1(_02049_),
    .S(net874),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _12571_ (.A0(_02050_),
    .A1(net2589),
    .S(net389),
    .X(_01274_));
 sky130_fd_sc_hd__or2_2 _12572_ (.A(_04275_),
    .B(_06663_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _12573_ (.A0(net588),
    .A1(net1910),
    .S(net470),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _12574_ (.A0(net585),
    .A1(net2350),
    .S(net469),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(net580),
    .A1(net2319),
    .S(net469),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _12576_ (.A0(net576),
    .A1(net2283),
    .S(net468),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(net571),
    .A1(net2268),
    .S(net468),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _12578_ (.A0(net541),
    .A1(net2211),
    .S(net468),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(net538),
    .A1(net2304),
    .S(net468),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _12580_ (.A0(net527),
    .A1(net1922),
    .S(net467),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(net521),
    .A1(net1911),
    .S(net467),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _12582_ (.A0(net408),
    .A1(net2402),
    .S(net468),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _12583_ (.A0(net403),
    .A1(net2023),
    .S(net467),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(net357),
    .A1(net2181),
    .S(net467),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(net352),
    .A1(net2030),
    .S(net467),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _12586_ (.A0(net349),
    .A1(net2159),
    .S(net467),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(net346),
    .A1(net2401),
    .S(net467),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(net341),
    .A1(net2223),
    .S(net467),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _12589_ (.A0(net338),
    .A1(net2141),
    .S(net468),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(net335),
    .A1(net2031),
    .S(net467),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(net331),
    .A1(net1913),
    .S(net467),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _12592_ (.A0(net327),
    .A1(net2425),
    .S(net470),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _12593_ (.A0(net322),
    .A1(net2215),
    .S(net468),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(net317),
    .A1(net2356),
    .S(net470),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _12595_ (.A0(net314),
    .A1(net2382),
    .S(net469),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(net309),
    .A1(net2027),
    .S(net468),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _12597_ (.A0(net306),
    .A1(net2381),
    .S(net469),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(net301),
    .A1(net2179),
    .S(net470),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _12599_ (.A0(net297),
    .A1(net2397),
    .S(net469),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(net293),
    .A1(net2353),
    .S(net469),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _12601_ (.A0(net291),
    .A1(net2503),
    .S(net469),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(net285),
    .A1(net2169),
    .S(net469),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _12603_ (.A0(net284),
    .A1(net2468),
    .S(net469),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(net279),
    .A1(net2352),
    .S(net469),
    .X(_01306_));
 sky130_fd_sc_hd__a22o_1 _12605_ (.A1(net1199),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[2] ),
    .B1(net916),
    .B2(net1179),
    .X(_02052_));
 sky130_fd_sc_hd__a21o_1 _12606_ (.A1(net2759),
    .A2(net894),
    .B1(_02052_),
    .X(_01307_));
 sky130_fd_sc_hd__a22o_1 _12607_ (.A1(net1199),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[3] ),
    .B1(net916),
    .B2(net119),
    .X(_02053_));
 sky130_fd_sc_hd__a21o_1 _12608_ (.A1(net2700),
    .A2(net894),
    .B1(_02053_),
    .X(_01308_));
 sky130_fd_sc_hd__nor2_1 _12609_ (.A(_02392_),
    .B(net912),
    .Y(_02054_));
 sky130_fd_sc_hd__a221o_1 _12610_ (.A1(net1199),
    .A2(net2950),
    .B1(net893),
    .B2(net3022),
    .C1(_02054_),
    .X(_01309_));
 sky130_fd_sc_hd__nor2_1 _12611_ (.A(_02393_),
    .B(net911),
    .Y(_02055_));
 sky130_fd_sc_hd__a221o_1 _12612_ (.A1(net1200),
    .A2(net2914),
    .B1(net893),
    .B2(\genblk1.genblk1.pcpi_mul.next_rs2[4] ),
    .C1(_02055_),
    .X(_01310_));
 sky130_fd_sc_hd__and3_1 _12613_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1224),
    .C(net1172),
    .X(_02056_));
 sky130_fd_sc_hd__a221o_1 _12614_ (.A1(net1200),
    .A2(net2902),
    .B1(net893),
    .B2(net2914),
    .C1(_02056_),
    .X(_01311_));
 sky130_fd_sc_hd__a22o_1 _12615_ (.A1(net1201),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[7] ),
    .B1(net916),
    .B2(net125),
    .X(_02057_));
 sky130_fd_sc_hd__a21o_1 _12616_ (.A1(net2902),
    .A2(net892),
    .B1(_02057_),
    .X(_01312_));
 sky130_fd_sc_hd__a22o_1 _12617_ (.A1(net1195),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[8] ),
    .B1(net915),
    .B2(net1169),
    .X(_02058_));
 sky130_fd_sc_hd__a21o_1 _12618_ (.A1(net2983),
    .A2(net888),
    .B1(_02058_),
    .X(_01313_));
 sky130_fd_sc_hd__a22o_1 _12619_ (.A1(net1195),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[9] ),
    .B1(net915),
    .B2(net1168),
    .X(_02059_));
 sky130_fd_sc_hd__a21o_1 _12620_ (.A1(net2668),
    .A2(net888),
    .B1(_02059_),
    .X(_01314_));
 sky130_fd_sc_hd__a22o_1 _12621_ (.A1(net1193),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[10] ),
    .B1(net915),
    .B2(net1167),
    .X(_02060_));
 sky130_fd_sc_hd__a21o_1 _12622_ (.A1(net2723),
    .A2(net888),
    .B1(_02060_),
    .X(_01315_));
 sky130_fd_sc_hd__and3_1 _12623_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1223),
    .C(net1166),
    .X(_02061_));
 sky130_fd_sc_hd__a221o_1 _12624_ (.A1(net1194),
    .A2(net2629),
    .B1(net887),
    .B2(net3004),
    .C1(_02061_),
    .X(_01316_));
 sky130_fd_sc_hd__a22o_1 _12625_ (.A1(net1194),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[12] ),
    .B1(net915),
    .B2(net1165),
    .X(_02062_));
 sky130_fd_sc_hd__a21o_1 _12626_ (.A1(net2629),
    .A2(net887),
    .B1(_02062_),
    .X(_01317_));
 sky130_fd_sc_hd__a22o_1 _12627_ (.A1(net1194),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[13] ),
    .B1(net915),
    .B2(net238),
    .X(_02063_));
 sky130_fd_sc_hd__a21o_1 _12628_ (.A1(net2830),
    .A2(net886),
    .B1(_02063_),
    .X(_01318_));
 sky130_fd_sc_hd__a22o_1 _12629_ (.A1(net1192),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[14] ),
    .B1(net915),
    .B2(net1163),
    .X(_02064_));
 sky130_fd_sc_hd__a21o_1 _12630_ (.A1(net2993),
    .A2(net885),
    .B1(_02064_),
    .X(_01319_));
 sky130_fd_sc_hd__nor2_1 _12631_ (.A(_02394_),
    .B(net911),
    .Y(_02065_));
 sky130_fd_sc_hd__a221o_1 _12632_ (.A1(net1192),
    .A2(net2814),
    .B1(net885),
    .B2(\genblk1.genblk1.pcpi_mul.next_rs2[14] ),
    .C1(_02065_),
    .X(_01320_));
 sky130_fd_sc_hd__a22o_1 _12633_ (.A1(net1198),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[16] ),
    .B1(net915),
    .B2(net1162),
    .X(_02066_));
 sky130_fd_sc_hd__a21o_1 _12634_ (.A1(net2814),
    .A2(net890),
    .B1(_02066_),
    .X(_01321_));
 sky130_fd_sc_hd__a22o_1 _12635_ (.A1(net1196),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[17] ),
    .B1(net914),
    .B2(net1161),
    .X(_02067_));
 sky130_fd_sc_hd__a21o_1 _12636_ (.A1(net2890),
    .A2(net890),
    .B1(_02067_),
    .X(_01322_));
 sky130_fd_sc_hd__a22o_1 _12637_ (.A1(net1196),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[18] ),
    .B1(net915),
    .B2(net1160),
    .X(_02068_));
 sky130_fd_sc_hd__a21o_1 _12638_ (.A1(net2633),
    .A2(net890),
    .B1(_02068_),
    .X(_01323_));
 sky130_fd_sc_hd__a22o_1 _12639_ (.A1(net1200),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[19] ),
    .B1(net919),
    .B2(net244),
    .X(_02069_));
 sky130_fd_sc_hd__a21o_1 _12640_ (.A1(net2970),
    .A2(net893),
    .B1(_02069_),
    .X(_01324_));
 sky130_fd_sc_hd__a22o_1 _12641_ (.A1(net1202),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[20] ),
    .B1(net916),
    .B2(net245),
    .X(_02070_));
 sky130_fd_sc_hd__a21o_1 _12642_ (.A1(net2752),
    .A2(net895),
    .B1(_02070_),
    .X(_01325_));
 sky130_fd_sc_hd__a22o_1 _12643_ (.A1(net1202),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[21] ),
    .B1(net916),
    .B2(net247),
    .X(_02071_));
 sky130_fd_sc_hd__a21o_1 _12644_ (.A1(net2763),
    .A2(net895),
    .B1(_02071_),
    .X(_01326_));
 sky130_fd_sc_hd__a22o_1 _12645_ (.A1(net1202),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[22] ),
    .B1(net916),
    .B2(net248),
    .X(_02072_));
 sky130_fd_sc_hd__a21o_1 _12646_ (.A1(net2823),
    .A2(net895),
    .B1(_02072_),
    .X(_01327_));
 sky130_fd_sc_hd__a22o_1 _12647_ (.A1(net1210),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[23] ),
    .B1(net918),
    .B2(net249),
    .X(_02073_));
 sky130_fd_sc_hd__a21o_1 _12648_ (.A1(net2923),
    .A2(net899),
    .B1(_02073_),
    .X(_01328_));
 sky130_fd_sc_hd__and3_1 _12649_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1227),
    .C(net250),
    .X(_02074_));
 sky130_fd_sc_hd__a221o_1 _12650_ (.A1(net1210),
    .A2(net2971),
    .B1(net899),
    .B2(net3002),
    .C1(_02074_),
    .X(_01329_));
 sky130_fd_sc_hd__nor2_1 _12651_ (.A(_02396_),
    .B(net913),
    .Y(_02075_));
 sky130_fd_sc_hd__a221o_1 _12652_ (.A1(net1210),
    .A2(net2724),
    .B1(net900),
    .B2(net2971),
    .C1(_02075_),
    .X(_01330_));
 sky130_fd_sc_hd__a22o_1 _12653_ (.A1(net1212),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[26] ),
    .B1(net918),
    .B2(net252),
    .X(_02076_));
 sky130_fd_sc_hd__a21o_1 _12654_ (.A1(net2724),
    .A2(net902),
    .B1(_02076_),
    .X(_01331_));
 sky130_fd_sc_hd__a22o_1 _12655_ (.A1(net1212),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[27] ),
    .B1(net917),
    .B2(net253),
    .X(_02077_));
 sky130_fd_sc_hd__a21o_1 _12656_ (.A1(net3014),
    .A2(net902),
    .B1(_02077_),
    .X(_01332_));
 sky130_fd_sc_hd__nor2_1 _12657_ (.A(_02397_),
    .B(net913),
    .Y(_02078_));
 sky130_fd_sc_hd__a221o_1 _12658_ (.A1(net1212),
    .A2(net2730),
    .B1(net902),
    .B2(net3009),
    .C1(_02078_),
    .X(_01333_));
 sky130_fd_sc_hd__a22o_1 _12659_ (.A1(net1212),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[29] ),
    .B1(net917),
    .B2(net255),
    .X(_02079_));
 sky130_fd_sc_hd__a21o_1 _12660_ (.A1(net2730),
    .A2(net902),
    .B1(_02079_),
    .X(_01334_));
 sky130_fd_sc_hd__nor2_1 _12661_ (.A(_02398_),
    .B(net913),
    .Y(_02080_));
 sky130_fd_sc_hd__a221o_1 _12662_ (.A1(net1212),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[30] ),
    .B1(net905),
    .B2(net3003),
    .C1(_02080_),
    .X(_01335_));
 sky130_fd_sc_hd__a22o_1 _12663_ (.A1(net1218),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[31] ),
    .B1(net917),
    .B2(net258),
    .X(_02081_));
 sky130_fd_sc_hd__a21o_1 _12664_ (.A1(net3027),
    .A2(net905),
    .B1(_02081_),
    .X(_01336_));
 sky130_fd_sc_hd__and3_1 _12665_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1237),
    .C(net1157),
    .X(_02082_));
 sky130_fd_sc_hd__a221o_1 _12666_ (.A1(net1218),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[32] ),
    .B1(net905),
    .B2(net3023),
    .C1(_02082_),
    .X(_01337_));
 sky130_fd_sc_hd__and2_2 _12667_ (.A(\genblk1.genblk1.pcpi_mul.instr_mulh ),
    .B(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__a221o_1 _12668_ (.A1(net1210),
    .A2(net2939),
    .B1(net899),
    .B2(\genblk1.genblk1.pcpi_mul.next_rs2[32] ),
    .C1(net713),
    .X(_01338_));
 sky130_fd_sc_hd__a221o_1 _12669_ (.A1(net1203),
    .A2(net3071),
    .B1(net899),
    .B2(net2939),
    .C1(net713),
    .X(_01339_));
 sky130_fd_sc_hd__a221o_1 _12670_ (.A1(net1202),
    .A2(net2979),
    .B1(net894),
    .B2(net3007),
    .C1(net713),
    .X(_01340_));
 sky130_fd_sc_hd__a221o_1 _12671_ (.A1(net1202),
    .A2(net2953),
    .B1(net894),
    .B2(net2979),
    .C1(net712),
    .X(_01341_));
 sky130_fd_sc_hd__a221o_1 _12672_ (.A1(net1200),
    .A2(net2894),
    .B1(net892),
    .B2(net2953),
    .C1(net712),
    .X(_01342_));
 sky130_fd_sc_hd__a221o_1 _12673_ (.A1(net1201),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[38] ),
    .B1(net892),
    .B2(net2894),
    .C1(net712),
    .X(_01343_));
 sky130_fd_sc_hd__a221o_1 _12674_ (.A1(net1201),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[39] ),
    .B1(net892),
    .B2(net3035),
    .C1(net712),
    .X(_01344_));
 sky130_fd_sc_hd__a221o_1 _12675_ (.A1(net1195),
    .A2(net3006),
    .B1(net889),
    .B2(\genblk1.genblk1.pcpi_mul.next_rs2[39] ),
    .C1(net712),
    .X(_01345_));
 sky130_fd_sc_hd__a221o_1 _12676_ (.A1(net1195),
    .A2(net2942),
    .B1(net888),
    .B2(net3006),
    .C1(net711),
    .X(_01346_));
 sky130_fd_sc_hd__a221o_1 _12677_ (.A1(net1197),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[42] ),
    .B1(net887),
    .B2(net2942),
    .C1(net711),
    .X(_01347_));
 sky130_fd_sc_hd__a221o_1 _12678_ (.A1(net1193),
    .A2(net2938),
    .B1(net886),
    .B2(net2975),
    .C1(net711),
    .X(_01348_));
 sky130_fd_sc_hd__a221o_1 _12679_ (.A1(net1193),
    .A2(net2826),
    .B1(net886),
    .B2(net2938),
    .C1(net711),
    .X(_01349_));
 sky130_fd_sc_hd__a221o_1 _12680_ (.A1(net1193),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[45] ),
    .B1(net886),
    .B2(net2826),
    .C1(net711),
    .X(_01350_));
 sky130_fd_sc_hd__a221o_1 _12681_ (.A1(net1194),
    .A2(net3070),
    .B1(net885),
    .B2(\genblk1.genblk1.pcpi_mul.next_rs2[45] ),
    .C1(net711),
    .X(_01351_));
 sky130_fd_sc_hd__a221o_1 _12682_ (.A1(net1194),
    .A2(net2915),
    .B1(net885),
    .B2(net2978),
    .C1(net711),
    .X(_01352_));
 sky130_fd_sc_hd__a221o_1 _12683_ (.A1(net1194),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[48] ),
    .B1(net886),
    .B2(net2915),
    .C1(net711),
    .X(_01353_));
 sky130_fd_sc_hd__a221o_1 _12684_ (.A1(net1196),
    .A2(net2928),
    .B1(net888),
    .B2(net2948),
    .C1(net711),
    .X(_01354_));
 sky130_fd_sc_hd__a221o_1 _12685_ (.A1(net1197),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[50] ),
    .B1(net889),
    .B2(net2928),
    .C1(net711),
    .X(_01355_));
 sky130_fd_sc_hd__a221o_1 _12686_ (.A1(net1195),
    .A2(net2845),
    .B1(net889),
    .B2(net3046),
    .C1(net712),
    .X(_01356_));
 sky130_fd_sc_hd__a221o_1 _12687_ (.A1(net1200),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[52] ),
    .B1(net895),
    .B2(net2845),
    .C1(net712),
    .X(_01357_));
 sky130_fd_sc_hd__a221o_1 _12688_ (.A1(net1203),
    .A2(net2905),
    .B1(net895),
    .B2(net2977),
    .C1(net713),
    .X(_01358_));
 sky130_fd_sc_hd__a221o_1 _12689_ (.A1(net1203),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[54] ),
    .B1(net895),
    .B2(net2905),
    .C1(net713),
    .X(_01359_));
 sky130_fd_sc_hd__a221o_1 _12690_ (.A1(net1210),
    .A2(net2955),
    .B1(net900),
    .B2(\genblk1.genblk1.pcpi_mul.next_rs2[54] ),
    .C1(net713),
    .X(_01360_));
 sky130_fd_sc_hd__a221o_1 _12691_ (.A1(net1211),
    .A2(net2952),
    .B1(net900),
    .B2(net2955),
    .C1(net713),
    .X(_01361_));
 sky130_fd_sc_hd__a221o_1 _12692_ (.A1(net1211),
    .A2(net2900),
    .B1(net903),
    .B2(net2952),
    .C1(net713),
    .X(_01362_));
 sky130_fd_sc_hd__a221o_1 _12693_ (.A1(net1211),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[58] ),
    .B1(net901),
    .B2(net2900),
    .C1(net713),
    .X(_01363_));
 sky130_fd_sc_hd__a221o_1 _12694_ (.A1(net1212),
    .A2(net2958),
    .B1(net901),
    .B2(net2969),
    .C1(net714),
    .X(_01364_));
 sky130_fd_sc_hd__a221o_1 _12695_ (.A1(net1213),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[60] ),
    .B1(net901),
    .B2(net2958),
    .C1(net714),
    .X(_01365_));
 sky130_fd_sc_hd__a221o_1 _12696_ (.A1(net1213),
    .A2(net2945),
    .B1(net901),
    .B2(net2963),
    .C1(net714),
    .X(_01366_));
 sky130_fd_sc_hd__a221o_1 _12697_ (.A1(net1217),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[62] ),
    .B1(net904),
    .B2(net2945),
    .C1(net714),
    .X(_01367_));
 sky130_fd_sc_hd__a221o_1 _12698_ (.A1(net1217),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs2[63] ),
    .B1(net904),
    .B2(net2956),
    .C1(net713),
    .X(_01368_));
 sky130_fd_sc_hd__a221o_1 _12699_ (.A1(net1217),
    .A2(net2527),
    .B1(net904),
    .B2(\genblk1.genblk1.pcpi_mul.next_rs2[63] ),
    .C1(net714),
    .X(_01369_));
 sky130_fd_sc_hd__nor2_1 _12700_ (.A(_02384_),
    .B(net912),
    .Y(_02084_));
 sky130_fd_sc_hd__a221o_1 _12701_ (.A1(net1199),
    .A2(net1098),
    .B1(net897),
    .B2(net2772),
    .C1(_02084_),
    .X(_01370_));
 sky130_fd_sc_hd__nor2_1 _12702_ (.A(_02383_),
    .B(net912),
    .Y(_02085_));
 sky130_fd_sc_hd__a221o_1 _12703_ (.A1(net1191),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[0] ),
    .B1(net2409),
    .B2(net897),
    .C1(_02085_),
    .X(_01371_));
 sky130_fd_sc_hd__a22o_1 _12704_ (.A1(net1191),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[1] ),
    .B1(net916),
    .B2(net1046),
    .X(_02086_));
 sky130_fd_sc_hd__a21o_1 _12705_ (.A1(net1491),
    .A2(net897),
    .B1(_02086_),
    .X(_01372_));
 sky130_fd_sc_hd__nor2_1 _12706_ (.A(_02402_),
    .B(net911),
    .Y(_02087_));
 sky130_fd_sc_hd__a221o_1 _12707_ (.A1(net1191),
    .A2(net1491),
    .B1(net2544),
    .B2(net897),
    .C1(_02087_),
    .X(_01373_));
 sky130_fd_sc_hd__a22o_1 _12708_ (.A1(net1198),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[3] ),
    .B1(net914),
    .B2(net1043),
    .X(_02088_));
 sky130_fd_sc_hd__a21o_1 _12709_ (.A1(net1339),
    .A2(net884),
    .B1(_02088_),
    .X(_01374_));
 sky130_fd_sc_hd__a22o_1 _12710_ (.A1(net1198),
    .A2(net1339),
    .B1(net914),
    .B2(net1041),
    .X(_02089_));
 sky130_fd_sc_hd__a21o_1 _12711_ (.A1(net1688),
    .A2(net884),
    .B1(_02089_),
    .X(_01375_));
 sky130_fd_sc_hd__a22o_1 _12712_ (.A1(net1192),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[5] ),
    .B1(net914),
    .B2(net231),
    .X(_02090_));
 sky130_fd_sc_hd__a21o_1 _12713_ (.A1(net1364),
    .A2(net883),
    .B1(_02090_),
    .X(_01376_));
 sky130_fd_sc_hd__a22o_1 _12714_ (.A1(net1192),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[6] ),
    .B1(net914),
    .B2(net1037),
    .X(_02091_));
 sky130_fd_sc_hd__a21o_1 _12715_ (.A1(net1354),
    .A2(net883),
    .B1(_02091_),
    .X(_01377_));
 sky130_fd_sc_hd__and3_1 _12716_ (.A(\genblk1.genblk1.pcpi_mul.mul_waiting ),
    .B(net1223),
    .C(net1034),
    .X(_02092_));
 sky130_fd_sc_hd__a221o_1 _12717_ (.A1(net1192),
    .A2(net1354),
    .B1(net2520),
    .B2(net883),
    .C1(_02092_),
    .X(_01378_));
 sky130_fd_sc_hd__nor2_1 _12718_ (.A(_02403_),
    .B(net911),
    .Y(_02093_));
 sky130_fd_sc_hd__a221o_1 _12719_ (.A1(net1190),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[8] ),
    .B1(net1542),
    .B2(net883),
    .C1(_02093_),
    .X(_01379_));
 sky130_fd_sc_hd__a22o_1 _12720_ (.A1(net1190),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[9] ),
    .B1(net914),
    .B2(net1030),
    .X(_02094_));
 sky130_fd_sc_hd__a21o_1 _12721_ (.A1(net1335),
    .A2(net883),
    .B1(_02094_),
    .X(_01380_));
 sky130_fd_sc_hd__nor2_1 _12722_ (.A(_02404_),
    .B(net911),
    .Y(_02095_));
 sky130_fd_sc_hd__a221o_1 _12723_ (.A1(net1190),
    .A2(net1335),
    .B1(net1732),
    .B2(net883),
    .C1(_02095_),
    .X(_01381_));
 sky130_fd_sc_hd__nor2_1 _12724_ (.A(_02405_),
    .B(net911),
    .Y(_02096_));
 sky130_fd_sc_hd__a221o_1 _12725_ (.A1(net1190),
    .A2(net1732),
    .B1(net2133),
    .B2(net883),
    .C1(_02096_),
    .X(_01382_));
 sky130_fd_sc_hd__nor2_1 _12726_ (.A(_02406_),
    .B(net911),
    .Y(_02097_));
 sky130_fd_sc_hd__a221o_1 _12727_ (.A1(net1190),
    .A2(net2133),
    .B1(net2421),
    .B2(net883),
    .C1(_02097_),
    .X(_01383_));
 sky130_fd_sc_hd__a22o_1 _12728_ (.A1(net1190),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[13] ),
    .B1(net914),
    .B2(net1023),
    .X(_02098_));
 sky130_fd_sc_hd__a21o_1 _12729_ (.A1(net1331),
    .A2(net883),
    .B1(_02098_),
    .X(_01384_));
 sky130_fd_sc_hd__a22o_1 _12730_ (.A1(net1190),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[14] ),
    .B1(net914),
    .B2(net1021),
    .X(_02099_));
 sky130_fd_sc_hd__a21o_1 _12731_ (.A1(net1326),
    .A2(net884),
    .B1(_02099_),
    .X(_01385_));
 sky130_fd_sc_hd__nor2_1 _12732_ (.A(_02407_),
    .B(net911),
    .Y(_02100_));
 sky130_fd_sc_hd__a221o_1 _12733_ (.A1(net1191),
    .A2(net1326),
    .B1(net2197),
    .B2(net884),
    .C1(_02100_),
    .X(_01386_));
 sky130_fd_sc_hd__nor2_1 _12734_ (.A(_02408_),
    .B(net911),
    .Y(_02101_));
 sky130_fd_sc_hd__a221o_1 _12735_ (.A1(net1191),
    .A2(net2197),
    .B1(net2364),
    .B2(net884),
    .C1(_02101_),
    .X(_01387_));
 sky130_fd_sc_hd__a22o_1 _12736_ (.A1(net1190),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[17] ),
    .B1(net914),
    .B2(net1015),
    .X(_02102_));
 sky130_fd_sc_hd__a21o_1 _12737_ (.A1(net1337),
    .A2(net884),
    .B1(_02102_),
    .X(_01388_));
 sky130_fd_sc_hd__nor2_1 _12738_ (.A(_02409_),
    .B(net912),
    .Y(_02103_));
 sky130_fd_sc_hd__a221o_1 _12739_ (.A1(net1190),
    .A2(net1337),
    .B1(net2089),
    .B2(net883),
    .C1(_02103_),
    .X(_01389_));
 sky130_fd_sc_hd__a22o_1 _12740_ (.A1(net1190),
    .A2(net2089),
    .B1(net914),
    .B2(net1011),
    .X(_02104_));
 sky130_fd_sc_hd__a21o_1 _12741_ (.A1(net2511),
    .A2(net897),
    .B1(_02104_),
    .X(_01390_));
 sky130_fd_sc_hd__nor2_1 _12742_ (.A(_02410_),
    .B(net912),
    .Y(_02105_));
 sky130_fd_sc_hd__a221o_1 _12743_ (.A1(net1191),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[20] ),
    .B1(net2105),
    .B2(net897),
    .C1(_02105_),
    .X(_01391_));
 sky130_fd_sc_hd__a22o_1 _12744_ (.A1(net1191),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[21] ),
    .B1(net916),
    .B2(net1008),
    .X(_02106_));
 sky130_fd_sc_hd__a21o_1 _12745_ (.A1(net1328),
    .A2(net897),
    .B1(_02106_),
    .X(_01392_));
 sky130_fd_sc_hd__nor2_1 _12746_ (.A(_02411_),
    .B(net911),
    .Y(_02107_));
 sky130_fd_sc_hd__a221o_1 _12747_ (.A1(net1191),
    .A2(net1328),
    .B1(net2392),
    .B2(net897),
    .C1(_02107_),
    .X(_01393_));
 sky130_fd_sc_hd__a22o_1 _12748_ (.A1(net1199),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[23] ),
    .B1(net916),
    .B2(net1005),
    .X(_02108_));
 sky130_fd_sc_hd__a21o_1 _12749_ (.A1(net2293),
    .A2(net897),
    .B1(_02108_),
    .X(_01394_));
 sky130_fd_sc_hd__a22o_1 _12750_ (.A1(net1214),
    .A2(net3068),
    .B1(net918),
    .B2(net1003),
    .X(_02109_));
 sky130_fd_sc_hd__a21o_1 _12751_ (.A1(net1550),
    .A2(net903),
    .B1(_02109_),
    .X(_01395_));
 sky130_fd_sc_hd__a22o_1 _12752_ (.A1(net1214),
    .A2(net1550),
    .B1(net918),
    .B2(net1001),
    .X(_02110_));
 sky130_fd_sc_hd__a21o_1 _12753_ (.A1(net1641),
    .A2(net899),
    .B1(_02110_),
    .X(_01396_));
 sky130_fd_sc_hd__a22o_1 _12754_ (.A1(net1214),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[26] ),
    .B1(net918),
    .B2(net999),
    .X(_02111_));
 sky130_fd_sc_hd__a21o_1 _12755_ (.A1(net1578),
    .A2(net899),
    .B1(_02111_),
    .X(_01397_));
 sky130_fd_sc_hd__nor2_1 _12756_ (.A(_02412_),
    .B(net913),
    .Y(_02112_));
 sky130_fd_sc_hd__a221o_1 _12757_ (.A1(net1214),
    .A2(net1578),
    .B1(net2575),
    .B2(net900),
    .C1(_02112_),
    .X(_01398_));
 sky130_fd_sc_hd__a22o_1 _12758_ (.A1(net1216),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[28] ),
    .B1(net917),
    .B2(net995),
    .X(_02113_));
 sky130_fd_sc_hd__a21o_1 _12759_ (.A1(net1450),
    .A2(net905),
    .B1(_02113_),
    .X(_01399_));
 sky130_fd_sc_hd__a22o_1 _12760_ (.A1(net1216),
    .A2(net1450),
    .B1(net918),
    .B2(net993),
    .X(_02114_));
 sky130_fd_sc_hd__a21o_1 _12761_ (.A1(net1836),
    .A2(net905),
    .B1(_02114_),
    .X(_01400_));
 sky130_fd_sc_hd__a221o_1 _12762_ (.A1(net1216),
    .A2(net1836),
    .B1(net2477),
    .B2(net907),
    .C1(_03876_),
    .X(_01401_));
 sky130_fd_sc_hd__a221o_1 _12763_ (.A1(net1216),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[31] ),
    .B1(net2337),
    .B2(net907),
    .C1(net762),
    .X(_01402_));
 sky130_fd_sc_hd__a221o_1 _12764_ (.A1(net1215),
    .A2(net2337),
    .B1(net2521),
    .B2(net906),
    .C1(net762),
    .X(_01403_));
 sky130_fd_sc_hd__a221o_1 _12765_ (.A1(net1215),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[33] ),
    .B1(net2501),
    .B2(net906),
    .C1(net762),
    .X(_01404_));
 sky130_fd_sc_hd__a221o_1 _12766_ (.A1(net1219),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[34] ),
    .B1(net2478),
    .B2(net907),
    .C1(net763),
    .X(_01405_));
 sky130_fd_sc_hd__a221o_1 _12767_ (.A1(net1219),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[35] ),
    .B1(net2472),
    .B2(net907),
    .C1(net763),
    .X(_01406_));
 sky130_fd_sc_hd__a221o_1 _12768_ (.A1(net1219),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[36] ),
    .B1(net2432),
    .B2(net906),
    .C1(net763),
    .X(_01407_));
 sky130_fd_sc_hd__a221o_1 _12769_ (.A1(net1219),
    .A2(net2432),
    .B1(net2594),
    .B2(net906),
    .C1(net763),
    .X(_01408_));
 sky130_fd_sc_hd__a221o_1 _12770_ (.A1(net1219),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[38] ),
    .B1(net2480),
    .B2(net908),
    .C1(net764),
    .X(_01409_));
 sky130_fd_sc_hd__a221o_1 _12771_ (.A1(net1219),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[39] ),
    .B1(net2289),
    .B2(net908),
    .C1(net764),
    .X(_01410_));
 sky130_fd_sc_hd__a221o_1 _12772_ (.A1(net1220),
    .A2(net2289),
    .B1(net2540),
    .B2(net908),
    .C1(net764),
    .X(_01411_));
 sky130_fd_sc_hd__a221o_1 _12773_ (.A1(net1220),
    .A2(net2540),
    .B1(net2573),
    .B2(net908),
    .C1(net764),
    .X(_01412_));
 sky130_fd_sc_hd__a221o_1 _12774_ (.A1(net1220),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[42] ),
    .B1(net2504),
    .B2(net908),
    .C1(net764),
    .X(_01413_));
 sky130_fd_sc_hd__a221o_1 _12775_ (.A1(net1220),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[43] ),
    .B1(net2107),
    .B2(net909),
    .C1(net764),
    .X(_01414_));
 sky130_fd_sc_hd__a221o_1 _12776_ (.A1(net1220),
    .A2(net2107),
    .B1(net2541),
    .B2(net909),
    .C1(net765),
    .X(_01415_));
 sky130_fd_sc_hd__a221o_1 _12777_ (.A1(net1220),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[45] ),
    .B1(net2517),
    .B2(net909),
    .C1(net765),
    .X(_01416_));
 sky130_fd_sc_hd__a221o_1 _12778_ (.A1(net1221),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[46] ),
    .B1(net2233),
    .B2(net909),
    .C1(net765),
    .X(_01417_));
 sky130_fd_sc_hd__a221o_1 _12779_ (.A1(net1221),
    .A2(net2233),
    .B1(net2489),
    .B2(net909),
    .C1(net765),
    .X(_01418_));
 sky130_fd_sc_hd__a221o_1 _12780_ (.A1(net1220),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[48] ),
    .B1(net2469),
    .B2(net908),
    .C1(net765),
    .X(_01419_));
 sky130_fd_sc_hd__a221o_1 _12781_ (.A1(net1220),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[49] ),
    .B1(net2264),
    .B2(net909),
    .C1(net765),
    .X(_01420_));
 sky130_fd_sc_hd__a221o_1 _12782_ (.A1(net1220),
    .A2(net2264),
    .B1(net2393),
    .B2(net908),
    .C1(net765),
    .X(_01421_));
 sky130_fd_sc_hd__a221o_1 _12783_ (.A1(net1220),
    .A2(net2393),
    .B1(net2519),
    .B2(net908),
    .C1(net764),
    .X(_01422_));
 sky130_fd_sc_hd__a221o_1 _12784_ (.A1(net1219),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[52] ),
    .B1(net2375),
    .B2(net908),
    .C1(net764),
    .X(_01423_));
 sky130_fd_sc_hd__a221o_1 _12785_ (.A1(net1219),
    .A2(net2375),
    .B1(net2443),
    .B2(net908),
    .C1(net764),
    .X(_01424_));
 sky130_fd_sc_hd__a221o_1 _12786_ (.A1(net1219),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[54] ),
    .B1(net2236),
    .B2(net907),
    .C1(net764),
    .X(_01425_));
 sky130_fd_sc_hd__a221o_1 _12787_ (.A1(net1219),
    .A2(net2236),
    .B1(net2286),
    .B2(net907),
    .C1(net763),
    .X(_01426_));
 sky130_fd_sc_hd__a221o_1 _12788_ (.A1(net1221),
    .A2(net2286),
    .B1(net2491),
    .B2(net906),
    .C1(net762),
    .X(_01427_));
 sky130_fd_sc_hd__a221o_1 _12789_ (.A1(net1221),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[57] ),
    .B1(net2367),
    .B2(net906),
    .C1(net762),
    .X(_01428_));
 sky130_fd_sc_hd__a221o_1 _12790_ (.A1(net1215),
    .A2(net2367),
    .B1(net2476),
    .B2(net906),
    .C1(net762),
    .X(_01429_));
 sky130_fd_sc_hd__a221o_1 _12791_ (.A1(net1215),
    .A2(net2476),
    .B1(net2508),
    .B2(net906),
    .C1(net762),
    .X(_01430_));
 sky130_fd_sc_hd__a221o_1 _12792_ (.A1(net1215),
    .A2(\genblk1.genblk1.pcpi_mul.next_rs1[60] ),
    .B1(net1961),
    .B2(net906),
    .C1(net762),
    .X(_01431_));
 sky130_fd_sc_hd__a221o_1 _12793_ (.A1(net1215),
    .A2(net1961),
    .B1(net1582),
    .B2(net906),
    .C1(net762),
    .X(_01432_));
 sky130_fd_sc_hd__or2_1 _12794_ (.A(\genblk1.genblk1.pcpi_mul.mul_counter[5] ),
    .B(_06670_),
    .X(_02115_));
 sky130_fd_sc_hd__a21oi_1 _12795_ (.A1(_02414_),
    .A2(_02115_),
    .B1(net918),
    .Y(_02116_));
 sky130_fd_sc_hd__o21a_1 _12796_ (.A1(_02414_),
    .A2(_02115_),
    .B1(_02116_),
    .X(_01433_));
 sky130_fd_sc_hd__or2_2 _12797_ (.A(_03745_),
    .B(_06663_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _12798_ (.A0(net588),
    .A1(net1938),
    .S(net465),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _12799_ (.A0(net585),
    .A1(net2074),
    .S(net465),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _12800_ (.A0(net579),
    .A1(net1884),
    .S(net465),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _12801_ (.A0(net575),
    .A1(net2311),
    .S(net464),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _12802_ (.A0(net571),
    .A1(net1881),
    .S(net465),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _12803_ (.A0(net543),
    .A1(net2064),
    .S(net464),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _12804_ (.A0(net538),
    .A1(net1846),
    .S(net463),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _12805_ (.A0(net527),
    .A1(net2242),
    .S(net463),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(net521),
    .A1(net2083),
    .S(net464),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _12807_ (.A0(net409),
    .A1(net2026),
    .S(net464),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _12808_ (.A0(net403),
    .A1(net2148),
    .S(net464),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(net357),
    .A1(net1914),
    .S(net463),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _12810_ (.A0(net352),
    .A1(net1781),
    .S(net463),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _12811_ (.A0(net349),
    .A1(net1996),
    .S(net463),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _12812_ (.A0(net346),
    .A1(net2200),
    .S(net463),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _12813_ (.A0(net341),
    .A1(net1972),
    .S(net463),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _12814_ (.A0(net338),
    .A1(net2189),
    .S(net463),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _12815_ (.A0(net335),
    .A1(net1971),
    .S(net463),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _12816_ (.A0(net331),
    .A1(net1872),
    .S(net463),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _12817_ (.A0(net327),
    .A1(net2307),
    .S(net465),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _12818_ (.A0(net323),
    .A1(net2068),
    .S(net464),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _12819_ (.A0(net317),
    .A1(net2069),
    .S(net465),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _12820_ (.A0(net315),
    .A1(net2016),
    .S(net465),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _12821_ (.A0(net309),
    .A1(net2257),
    .S(net464),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _12822_ (.A0(net306),
    .A1(net2058),
    .S(net466),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _12823_ (.A0(net301),
    .A1(net2086),
    .S(net465),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _12824_ (.A0(net297),
    .A1(net1842),
    .S(net465),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(net293),
    .A1(net1979),
    .S(net466),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _12826_ (.A0(net291),
    .A1(net1923),
    .S(net466),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _12827_ (.A0(net285),
    .A1(net1724),
    .S(net465),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _12828_ (.A0(net284),
    .A1(net2128),
    .S(net466),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _12829_ (.A0(net279),
    .A1(net2119),
    .S(net466),
    .X(_01465_));
 sky130_fd_sc_hd__or2_4 _12830_ (.A(_03742_),
    .B(_04283_),
    .X(_02118_));
 sky130_fd_sc_hd__mux2_1 _12831_ (.A0(net587),
    .A1(net2308),
    .S(net461),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _12832_ (.A0(net584),
    .A1(net2460),
    .S(net461),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _12833_ (.A0(net581),
    .A1(net2203),
    .S(net462),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _12834_ (.A0(net577),
    .A1(net2274),
    .S(net459),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _12835_ (.A0(net574),
    .A1(net2292),
    .S(net462),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _12836_ (.A0(net542),
    .A1(net2448),
    .S(net459),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _12837_ (.A0(net539),
    .A1(net2390),
    .S(net459),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _12838_ (.A0(_03774_),
    .A1(net2345),
    .S(net460),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _12839_ (.A0(net520),
    .A1(net2110),
    .S(net460),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _12840_ (.A0(net409),
    .A1(net2240),
    .S(net460),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(net405),
    .A1(net2049),
    .S(net460),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _12842_ (.A0(net355),
    .A1(net2157),
    .S(net460),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(net351),
    .A1(net2339),
    .S(net459),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _12844_ (.A0(net347),
    .A1(net2245),
    .S(net459),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _12845_ (.A0(net344),
    .A1(net2380),
    .S(net460),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(net339),
    .A1(net2176),
    .S(net459),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _12847_ (.A0(net337),
    .A1(net2306),
    .S(net459),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _12848_ (.A0(net333),
    .A1(net2522),
    .S(net459),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _12849_ (.A0(net328),
    .A1(net2147),
    .S(net459),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _12850_ (.A0(net325),
    .A1(net2357),
    .S(net461),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(net321),
    .A1(net2260),
    .S(net459),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _12852_ (.A0(net316),
    .A1(net2057),
    .S(net461),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(net313),
    .A1(net2429),
    .S(net461),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _12854_ (.A0(net311),
    .A1(net2454),
    .S(net461),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(net306),
    .A1(net2395),
    .S(net462),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _12856_ (.A0(net302),
    .A1(net2287),
    .S(net462),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _12857_ (.A0(net298),
    .A1(net2252),
    .S(net462),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _12858_ (.A0(net293),
    .A1(net2492),
    .S(net461),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(net289),
    .A1(net2383),
    .S(net461),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(net285),
    .A1(net2104),
    .S(net462),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(net283),
    .A1(net2295),
    .S(net461),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _12862_ (.A0(net278),
    .A1(net2466),
    .S(net461),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _12863_ (.A0(net1),
    .A1(net2699),
    .S(_02450_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _12864_ (.A0(net12),
    .A1(net2645),
    .S(_02450_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(net23),
    .A1(\mem_rdata_q[2] ),
    .S(_02450_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _12866_ (.A0(net26),
    .A1(net2793),
    .S(_02450_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _12867_ (.A0(net27),
    .A1(net2936),
    .S(_02450_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _12868_ (.A0(net28),
    .A1(net3015),
    .S(_02450_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _12869_ (.A0(net29),
    .A1(net2947),
    .S(_02450_),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _12870_ (.A0(\mem_rdata_q[7] ),
    .A1(net30),
    .S(net962),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _12871_ (.A0(\mem_rdata_q[8] ),
    .A1(net31),
    .S(net963),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _12872_ (.A0(\mem_rdata_q[9] ),
    .A1(net32),
    .S(net963),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _12873_ (.A0(\mem_rdata_q[10] ),
    .A1(net2),
    .S(net964),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(\mem_rdata_q[11] ),
    .A1(net3),
    .S(net963),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _12875_ (.A0(\mem_rdata_q[12] ),
    .A1(net4),
    .S(net963),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(\mem_rdata_q[13] ),
    .A1(net5),
    .S(net963),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _12877_ (.A0(\mem_rdata_q[14] ),
    .A1(net6),
    .S(net962),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(\mem_rdata_q[15] ),
    .A1(net7),
    .S(net962),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _12879_ (.A0(\mem_rdata_q[16] ),
    .A1(net8),
    .S(net962),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _12880_ (.A0(\mem_rdata_q[17] ),
    .A1(net9),
    .S(net962),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _12881_ (.A0(\mem_rdata_q[18] ),
    .A1(net10),
    .S(net962),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _12882_ (.A0(\mem_rdata_q[19] ),
    .A1(net11),
    .S(net962),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _12883_ (.A0(\mem_rdata_q[20] ),
    .A1(net13),
    .S(net964),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _12884_ (.A0(\mem_rdata_q[21] ),
    .A1(net14),
    .S(net962),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _12885_ (.A0(\mem_rdata_q[22] ),
    .A1(net15),
    .S(net962),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _12886_ (.A0(\mem_rdata_q[23] ),
    .A1(net16),
    .S(net964),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _12887_ (.A0(\mem_rdata_q[24] ),
    .A1(net17),
    .S(net964),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(\mem_rdata_q[25] ),
    .A1(net18),
    .S(net964),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _12889_ (.A0(\mem_rdata_q[26] ),
    .A1(net19),
    .S(net964),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _12890_ (.A0(\mem_rdata_q[27] ),
    .A1(net20),
    .S(net964),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _12891_ (.A0(\mem_rdata_q[28] ),
    .A1(net21),
    .S(net964),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _12892_ (.A0(\mem_rdata_q[29] ),
    .A1(net22),
    .S(net964),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _12893_ (.A0(\mem_rdata_q[30] ),
    .A1(net24),
    .S(net965),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(\mem_rdata_q[31] ),
    .A1(net25),
    .S(net962),
    .X(_01529_));
 sky130_fd_sc_hd__or2_2 _12895_ (.A(_04283_),
    .B(_06663_),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _12896_ (.A0(net588),
    .A1(net2340),
    .S(net457),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _12897_ (.A0(net585),
    .A1(net2444),
    .S(net457),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _12898_ (.A0(net579),
    .A1(net2099),
    .S(net457),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _12899_ (.A0(net576),
    .A1(net1907),
    .S(net456),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _12900_ (.A0(net571),
    .A1(net1967),
    .S(net457),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _12901_ (.A0(net543),
    .A1(net2323),
    .S(net456),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _12902_ (.A0(net538),
    .A1(net2038),
    .S(net455),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _12903_ (.A0(net527),
    .A1(net2249),
    .S(net455),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _12904_ (.A0(net521),
    .A1(net2102),
    .S(net456),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _12905_ (.A0(net409),
    .A1(net2117),
    .S(net456),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _12906_ (.A0(net404),
    .A1(net2005),
    .S(net456),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _12907_ (.A0(net357),
    .A1(net1926),
    .S(net455),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _12908_ (.A0(net352),
    .A1(net2006),
    .S(net455),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _12909_ (.A0(net349),
    .A1(net1960),
    .S(net455),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _12910_ (.A0(net346),
    .A1(net2347),
    .S(net455),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _12911_ (.A0(net341),
    .A1(net2139),
    .S(net455),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _12912_ (.A0(net338),
    .A1(net2365),
    .S(net455),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _12913_ (.A0(net335),
    .A1(net2449),
    .S(net455),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _12914_ (.A0(net331),
    .A1(net2153),
    .S(net455),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _12915_ (.A0(net326),
    .A1(net2278),
    .S(net457),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _12916_ (.A0(net323),
    .A1(net2034),
    .S(net456),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _12917_ (.A0(net317),
    .A1(net2336),
    .S(net457),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _12918_ (.A0(net314),
    .A1(net2437),
    .S(net457),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _12919_ (.A0(net309),
    .A1(net2471),
    .S(net456),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _12920_ (.A0(net306),
    .A1(net2384),
    .S(net458),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _12921_ (.A0(net301),
    .A1(net1956),
    .S(net457),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _12922_ (.A0(net297),
    .A1(net1793),
    .S(net457),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _12923_ (.A0(net294),
    .A1(net2438),
    .S(net458),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _12924_ (.A0(net291),
    .A1(net2463),
    .S(net458),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(net285),
    .A1(net2314),
    .S(net457),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _12926_ (.A0(net284),
    .A1(net2253),
    .S(net458),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _12927_ (.A0(net279),
    .A1(net2404),
    .S(net458),
    .X(_01561_));
 sky130_fd_sc_hd__and3b_1 _12928_ (.A_N(net174),
    .B(_06611_),
    .C(net175),
    .X(_01562_));
 sky130_fd_sc_hd__and3b_1 _12929_ (.A_N(net175),
    .B(net174),
    .C(_06611_),
    .X(_01563_));
 sky130_fd_sc_hd__a221o_1 _12930_ (.A1(net1066),
    .A2(_02385_),
    .B1(\decoded_imm_j[11] ),
    .B2(_02701_),
    .C1(net710),
    .X(_02120_));
 sky130_fd_sc_hd__o22a_1 _12931_ (.A1(net3016),
    .A2(_02502_),
    .B1(_05169_),
    .B2(_02120_),
    .X(_01564_));
 sky130_fd_sc_hd__a32o_1 _12932_ (.A1(net1066),
    .A2(\reg_sh[1] ),
    .A3(\reg_sh[0] ),
    .B1(\decoded_imm_j[1] ),
    .B2(_02701_),
    .X(_02121_));
 sky130_fd_sc_hd__o32a_1 _12933_ (.A1(_03192_),
    .A2(_05204_),
    .A3(_02121_),
    .B1(_02502_),
    .B2(net2170),
    .X(_01565_));
 sky130_fd_sc_hd__or2_1 _12934_ (.A(_03744_),
    .B(_04283_),
    .X(_02122_));
 sky130_fd_sc_hd__mux2_1 _12935_ (.A0(net588),
    .A1(net2532),
    .S(net453),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _12936_ (.A0(net585),
    .A1(net2415),
    .S(net453),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _12937_ (.A0(net580),
    .A1(net2184),
    .S(net453),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _12938_ (.A0(net576),
    .A1(net2114),
    .S(net451),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _12939_ (.A0(net571),
    .A1(net2036),
    .S(net451),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(net541),
    .A1(net2316),
    .S(net454),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _12941_ (.A0(net537),
    .A1(net1848),
    .S(net451),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _12942_ (.A0(net526),
    .A1(net2261),
    .S(net451),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _12943_ (.A0(net521),
    .A1(net2202),
    .S(net451),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(net408),
    .A1(net2185),
    .S(net451),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _12945_ (.A0(net403),
    .A1(net2142),
    .S(net451),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _12946_ (.A0(net356),
    .A1(net2434),
    .S(net451),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _12947_ (.A0(net353),
    .A1(net2231),
    .S(net452),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _12948_ (.A0(net349),
    .A1(net2024),
    .S(net452),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _12949_ (.A0(net346),
    .A1(net2196),
    .S(net451),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _12950_ (.A0(net342),
    .A1(net1944),
    .S(net452),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _12951_ (.A0(net338),
    .A1(net2155),
    .S(net452),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _12952_ (.A0(net334),
    .A1(net2178),
    .S(net452),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _12953_ (.A0(net331),
    .A1(net1951),
    .S(net452),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _12954_ (.A0(net326),
    .A1(net2427),
    .S(net452),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _12955_ (.A0(net323),
    .A1(net2028),
    .S(net452),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _12956_ (.A0(net317),
    .A1(net2065),
    .S(net452),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _12957_ (.A0(net315),
    .A1(net2414),
    .S(net453),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _12958_ (.A0(net309),
    .A1(net2164),
    .S(net451),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _12959_ (.A0(net306),
    .A1(net2209),
    .S(net453),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _12960_ (.A0(net301),
    .A1(net2172),
    .S(net454),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _12961_ (.A0(net297),
    .A1(net2035),
    .S(net454),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _12962_ (.A0(net293),
    .A1(net2227),
    .S(net453),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _12963_ (.A0(net291),
    .A1(net2495),
    .S(net453),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _12964_ (.A0(net286),
    .A1(net2453),
    .S(net453),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _12965_ (.A0(net284),
    .A1(net2456),
    .S(net453),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _12966_ (.A0(net279),
    .A1(net2525),
    .S(net453),
    .X(_01597_));
 sky130_fd_sc_hd__nor2_1 _12967_ (.A(_03745_),
    .B(_04281_),
    .Y(_02123_));
 sky130_fd_sc_hd__mux2_1 _12968_ (.A0(net1397),
    .A1(net586),
    .S(net449),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _12969_ (.A0(net1785),
    .A1(net585),
    .S(net449),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _12970_ (.A0(net1874),
    .A1(net582),
    .S(net449),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _12971_ (.A0(net1532),
    .A1(net578),
    .S(net448),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _12972_ (.A0(net1821),
    .A1(net573),
    .S(net448),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _12973_ (.A0(net1871),
    .A1(net542),
    .S(net448),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _12974_ (.A0(net1497),
    .A1(net539),
    .S(net447),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _12975_ (.A0(net1739),
    .A1(net525),
    .S(net447),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _12976_ (.A0(net1712),
    .A1(net523),
    .S(net447),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _12977_ (.A0(net1695),
    .A1(_03782_),
    .S(net447),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _12978_ (.A0(net1622),
    .A1(net406),
    .S(net448),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _12979_ (.A0(net1563),
    .A1(net354),
    .S(net448),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _12980_ (.A0(net1344),
    .A1(net350),
    .S(net447),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _12981_ (.A0(net1480),
    .A1(net347),
    .S(net447),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _12982_ (.A0(net1632),
    .A1(net343),
    .S(net447),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _12983_ (.A0(net1518),
    .A1(net340),
    .S(net447),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _12984_ (.A0(net2127),
    .A1(net338),
    .S(net448),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _12985_ (.A0(net1812),
    .A1(net333),
    .S(net447),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _12986_ (.A0(net1346),
    .A1(net330),
    .S(net447),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _12987_ (.A0(net1567),
    .A1(net327),
    .S(net449),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _12988_ (.A0(net1425),
    .A1(net323),
    .S(net448),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _12989_ (.A0(net1541),
    .A1(net318),
    .S(net448),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _12990_ (.A0(net1826),
    .A1(net314),
    .S(net449),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _12991_ (.A0(net1442),
    .A1(net310),
    .S(net449),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _12992_ (.A0(net1381),
    .A1(net307),
    .S(net449),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _12993_ (.A0(net1510),
    .A1(net303),
    .S(net450),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _12994_ (.A0(net2547),
    .A1(net300),
    .S(net450),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _12995_ (.A0(net1672),
    .A1(net296),
    .S(net450),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _12996_ (.A0(net1408),
    .A1(net292),
    .S(net449),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _12997_ (.A0(net1638),
    .A1(net287),
    .S(net449),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _12998_ (.A0(net1428),
    .A1(net284),
    .S(net449),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _12999_ (.A0(net1527),
    .A1(net280),
    .S(net450),
    .X(_01638_));
 sky130_fd_sc_hd__and2_1 _13000_ (.A(_06255_),
    .B(_06611_),
    .X(_01639_));
 sky130_fd_sc_hd__and2_1 _13001_ (.A(net2515),
    .B(net907),
    .X(_01640_));
 sky130_fd_sc_hd__or2_1 _13002_ (.A(_04272_),
    .B(_04275_),
    .X(_02124_));
 sky130_fd_sc_hd__mux2_1 _13003_ (.A0(_03749_),
    .A1(net2328),
    .S(net445),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _13004_ (.A0(net584),
    .A1(net2280),
    .S(net445),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _13005_ (.A0(net580),
    .A1(net2344),
    .S(net445),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _13006_ (.A0(net575),
    .A1(net2333),
    .S(net444),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _13007_ (.A0(net572),
    .A1(net2220),
    .S(net445),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _13008_ (.A0(net541),
    .A1(net2243),
    .S(net444),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _13009_ (.A0(net538),
    .A1(net2394),
    .S(net443),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _13010_ (.A0(net526),
    .A1(net2299),
    .S(net443),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _13011_ (.A0(net521),
    .A1(net2447),
    .S(net443),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _13012_ (.A0(net408),
    .A1(net2317),
    .S(net443),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _13013_ (.A0(net403),
    .A1(net2134),
    .S(net444),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _13014_ (.A0(net356),
    .A1(net1984),
    .S(net443),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _13015_ (.A0(net352),
    .A1(net2269),
    .S(net443),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _13016_ (.A0(net349),
    .A1(net2198),
    .S(net443),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _13017_ (.A0(net346),
    .A1(net2162),
    .S(net444),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _13018_ (.A0(net341),
    .A1(net2152),
    .S(net443),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _13019_ (.A0(net337),
    .A1(net2488),
    .S(net444),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _13020_ (.A0(net334),
    .A1(net2235),
    .S(net443),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _13021_ (.A0(net331),
    .A1(net2462),
    .S(net443),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _13022_ (.A0(net326),
    .A1(net2284),
    .S(net445),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _13023_ (.A0(net322),
    .A1(net2194),
    .S(net444),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _13024_ (.A0(net317),
    .A1(net2391),
    .S(net444),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _13025_ (.A0(net313),
    .A1(net2371),
    .S(net445),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _13026_ (.A0(net308),
    .A1(net2465),
    .S(net444),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _13027_ (.A0(net305),
    .A1(net2377),
    .S(net445),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _13028_ (.A0(net304),
    .A1(net2330),
    .S(net446),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _13029_ (.A0(net299),
    .A1(net2510),
    .S(net445),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _13030_ (.A0(net296),
    .A1(net2334),
    .S(net445),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(net289),
    .A1(net2273),
    .S(net446),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _13032_ (.A0(net287),
    .A1(net2313),
    .S(net446),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _13033_ (.A0(net282),
    .A1(net2342),
    .S(net445),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _13034_ (.A0(net281),
    .A1(net2490),
    .S(net446),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _13035_ (.A0(net1459),
    .A1(net86),
    .S(net535),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _13036_ (.A0(net1593),
    .A1(net89),
    .S(net535),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _13037_ (.A0(net1366),
    .A1(net90),
    .S(net535),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _13038_ (.A0(net1464),
    .A1(net91),
    .S(net535),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _13039_ (.A0(net1348),
    .A1(net92),
    .S(net535),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _13040_ (.A0(net1333),
    .A1(net93),
    .S(net535),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(net1345),
    .A1(net94),
    .S(net535),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _13042_ (.A0(net1334),
    .A1(net95),
    .S(net535),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _13043_ (.A0(net1419),
    .A1(net66),
    .S(net535),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _13044_ (.A0(net1347),
    .A1(net67),
    .S(net534),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _13045_ (.A0(net1477),
    .A1(net68),
    .S(net534),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _13046_ (.A0(net1352),
    .A1(net69),
    .S(net534),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _13047_ (.A0(net1363),
    .A1(net70),
    .S(net535),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _13048_ (.A0(net1681),
    .A1(net71),
    .S(net534),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _13049_ (.A0(net1623),
    .A1(net72),
    .S(net534),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _13050_ (.A0(net1494),
    .A1(net73),
    .S(net534),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _13051_ (.A0(net1585),
    .A1(net74),
    .S(net533),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _13052_ (.A0(net1827),
    .A1(net75),
    .S(net533),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _13053_ (.A0(net1723),
    .A1(net76),
    .S(net533),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _13054_ (.A0(net1461),
    .A1(net77),
    .S(net533),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _13055_ (.A0(net2001),
    .A1(net78),
    .S(net533),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _13056_ (.A0(net1596),
    .A1(net79),
    .S(net533),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _13057_ (.A0(net2467),
    .A1(net80),
    .S(net536),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _13058_ (.A0(net1373),
    .A1(net81),
    .S(net536),
    .X(_01696_));
 sky130_fd_sc_hd__mux2_1 _13059_ (.A0(net1646),
    .A1(net82),
    .S(net533),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(net1614),
    .A1(net83),
    .S(net533),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _13061_ (.A0(net1556),
    .A1(net84),
    .S(net533),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _13062_ (.A0(net2498),
    .A1(net85),
    .S(net534),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _13063_ (.A0(net1439),
    .A1(net87),
    .S(net533),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _13064_ (.A0(net2258),
    .A1(net88),
    .S(net534),
    .X(_01702_));
 sky130_fd_sc_hd__or2_1 _13065_ (.A(_03745_),
    .B(_04272_),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _13066_ (.A0(net586),
    .A1(net2161),
    .S(net441),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _13067_ (.A0(net584),
    .A1(net2277),
    .S(net442),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _13068_ (.A0(net579),
    .A1(net1953),
    .S(net441),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _13069_ (.A0(net575),
    .A1(net2008),
    .S(net440),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _13070_ (.A0(net572),
    .A1(net2160),
    .S(net441),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _13071_ (.A0(net544),
    .A1(net2205),
    .S(net440),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _13072_ (.A0(net537),
    .A1(net1770),
    .S(net439),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _13073_ (.A0(net526),
    .A1(net1716),
    .S(net439),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _13074_ (.A0(net521),
    .A1(net1895),
    .S(net439),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _13075_ (.A0(net407),
    .A1(net1631),
    .S(net439),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _13076_ (.A0(net403),
    .A1(net1639),
    .S(net440),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _13077_ (.A0(net356),
    .A1(net1893),
    .S(net439),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _13078_ (.A0(net352),
    .A1(net1833),
    .S(net439),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _13079_ (.A0(net349),
    .A1(net1733),
    .S(net439),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _13080_ (.A0(net346),
    .A1(net1682),
    .S(net440),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _13081_ (.A0(net341),
    .A1(net1628),
    .S(net439),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _13082_ (.A0(net337),
    .A1(net2060),
    .S(net440),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _13083_ (.A0(net334),
    .A1(net1815),
    .S(net439),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _13084_ (.A0(net329),
    .A1(net1561),
    .S(net439),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _13085_ (.A0(net325),
    .A1(net2025),
    .S(net441),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _13086_ (.A0(net321),
    .A1(net2003),
    .S(net440),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _13087_ (.A0(net318),
    .A1(net1698),
    .S(net440),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _13088_ (.A0(net313),
    .A1(net2062),
    .S(net441),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _13089_ (.A0(net308),
    .A1(net1814),
    .S(net440),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _13090_ (.A0(net305),
    .A1(net2318),
    .S(net441),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _13091_ (.A0(net304),
    .A1(net1902),
    .S(net442),
    .X(_01728_));
 sky130_fd_sc_hd__mux2_1 _13092_ (.A0(net299),
    .A1(net1985),
    .S(net441),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _13093_ (.A0(net296),
    .A1(net2335),
    .S(net441),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(net290),
    .A1(net2130),
    .S(net441),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _13095_ (.A0(net286),
    .A1(net2386),
    .S(net441),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _13096_ (.A0(net283),
    .A1(net1917),
    .S(net442),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _13097_ (.A0(net279),
    .A1(net2175),
    .S(net442),
    .X(_01734_));
 sky130_fd_sc_hd__or2_1 _13098_ (.A(_04272_),
    .B(_04283_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _13099_ (.A0(net588),
    .A1(net2497),
    .S(net437),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_1 _13100_ (.A0(net584),
    .A1(net2507),
    .S(net438),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _13101_ (.A0(net579),
    .A1(net2461),
    .S(net437),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _13102_ (.A0(net575),
    .A1(net2405),
    .S(net436),
    .X(_01738_));
 sky130_fd_sc_hd__mux2_1 _13103_ (.A0(net572),
    .A1(net2183),
    .S(net437),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _13104_ (.A0(net544),
    .A1(net2310),
    .S(net436),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _13105_ (.A0(net537),
    .A1(net2451),
    .S(net435),
    .X(_01741_));
 sky130_fd_sc_hd__mux2_1 _13106_ (.A0(net526),
    .A1(net2248),
    .S(net435),
    .X(_01742_));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(net521),
    .A1(net2408),
    .S(net435),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _13108_ (.A0(net407),
    .A1(net2207),
    .S(net435),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _13109_ (.A0(net403),
    .A1(net2121),
    .S(net436),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _13110_ (.A0(net356),
    .A1(net2097),
    .S(net435),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(net352),
    .A1(net2239),
    .S(net435),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_1 _13112_ (.A0(net349),
    .A1(net2138),
    .S(net435),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _13113_ (.A0(net346),
    .A1(net2126),
    .S(net436),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _13114_ (.A0(net341),
    .A1(net2270),
    .S(net435),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _13115_ (.A0(net337),
    .A1(net2213),
    .S(net436),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _13116_ (.A0(net334),
    .A1(net2354),
    .S(net435),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(net329),
    .A1(net2464),
    .S(net435),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _13118_ (.A0(net325),
    .A1(net2424),
    .S(net437),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _13119_ (.A0(net321),
    .A1(net2276),
    .S(net436),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _13120_ (.A0(net318),
    .A1(net2259),
    .S(net436),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(net313),
    .A1(net2343),
    .S(net437),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _13122_ (.A0(net308),
    .A1(net2360),
    .S(net436),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _13123_ (.A0(net305),
    .A1(net2302),
    .S(net437),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _13124_ (.A0(net304),
    .A1(net2496),
    .S(net438),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _13125_ (.A0(net299),
    .A1(net2500),
    .S(net437),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _13126_ (.A0(net296),
    .A1(net2294),
    .S(net437),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _13127_ (.A0(net290),
    .A1(net2509),
    .S(net437),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _13128_ (.A0(net286),
    .A1(net2399),
    .S(net437),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _13129_ (.A0(net282),
    .A1(net2486),
    .S(net438),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _13130_ (.A0(net281),
    .A1(net2378),
    .S(net438),
    .X(_01766_));
 sky130_fd_sc_hd__nand3b_1 _13131_ (.A_N(\latched_rd[4] ),
    .B(\latched_rd[3] ),
    .C(\latched_rd[2] ),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _13132_ (.A(_04273_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__mux2_1 _13133_ (.A0(net1535),
    .A1(net588),
    .S(net433),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(net1484),
    .A1(net583),
    .S(net433),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _13135_ (.A0(net1444),
    .A1(net579),
    .S(net433),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(net1489),
    .A1(net575),
    .S(net432),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _13137_ (.A0(net1601),
    .A1(net571),
    .S(net433),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _13138_ (.A0(net1524),
    .A1(net541),
    .S(net432),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _13139_ (.A0(net1670),
    .A1(net537),
    .S(net431),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _13140_ (.A0(net1463),
    .A1(net526),
    .S(net431),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _13141_ (.A0(net1472),
    .A1(net520),
    .S(net431),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _13142_ (.A0(net1588),
    .A1(net407),
    .S(net431),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _13143_ (.A0(net1367),
    .A1(net404),
    .S(net432),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _13144_ (.A0(net1409),
    .A1(net357),
    .S(net431),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _13145_ (.A0(net1946),
    .A1(net351),
    .S(net431),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _13146_ (.A0(net1499),
    .A1(net348),
    .S(net431),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _13147_ (.A0(net1476),
    .A1(net345),
    .S(net432),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _13148_ (.A0(net1615),
    .A1(net341),
    .S(net431),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _13149_ (.A0(net1448),
    .A1(net336),
    .S(net432),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _13150_ (.A0(net1664),
    .A1(net334),
    .S(net431),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(net1493),
    .A1(net328),
    .S(net431),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _13152_ (.A0(net1625),
    .A1(net325),
    .S(net433),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(net1647),
    .A1(net320),
    .S(net432),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _13154_ (.A0(net1759),
    .A1(net318),
    .S(net432),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _13155_ (.A0(net1680),
    .A1(net312),
    .S(net433),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _13156_ (.A0(net1506),
    .A1(net308),
    .S(net432),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _13157_ (.A0(net2324),
    .A1(net305),
    .S(net433),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _13158_ (.A0(net1412),
    .A1(net303),
    .S(net434),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(net1832),
    .A1(net300),
    .S(net433),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _13160_ (.A0(net1375),
    .A1(net295),
    .S(net433),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _13161_ (.A0(net2389),
    .A1(net290),
    .S(net434),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _13162_ (.A0(net1396),
    .A1(net287),
    .S(net433),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _13163_ (.A0(net1458),
    .A1(_03870_),
    .S(net434),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _13164_ (.A0(net1594),
    .A1(net281),
    .S(net434),
    .X(_01798_));
 sky130_fd_sc_hd__nor2_1 _13165_ (.A(_04275_),
    .B(_02127_),
    .Y(_02129_));
 sky130_fd_sc_hd__mux2_1 _13166_ (.A0(net2059),
    .A1(net588),
    .S(net429),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _13167_ (.A0(net1915),
    .A1(net583),
    .S(net429),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _13168_ (.A0(net1526),
    .A1(net579),
    .S(net429),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _13169_ (.A0(net1470),
    .A1(net575),
    .S(net428),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _13170_ (.A0(net1640),
    .A1(net571),
    .S(net429),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _13171_ (.A0(net1753),
    .A1(net541),
    .S(net428),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _13172_ (.A0(net1549),
    .A1(net537),
    .S(net427),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _13173_ (.A0(net2116),
    .A1(net526),
    .S(net427),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _13174_ (.A0(net1540),
    .A1(net520),
    .S(net427),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _13175_ (.A0(net1824),
    .A1(net407),
    .S(net427),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(net1755),
    .A1(net404),
    .S(net428),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _13177_ (.A0(net1566),
    .A1(net357),
    .S(net427),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _13178_ (.A0(net1806),
    .A1(net351),
    .S(net427),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _13179_ (.A0(net1883),
    .A1(_03799_),
    .S(net427),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(net1857),
    .A1(net345),
    .S(net428),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _13181_ (.A0(net1574),
    .A1(net341),
    .S(net427),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _13182_ (.A0(net1777),
    .A1(net337),
    .S(net428),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _13183_ (.A0(net1671),
    .A1(net334),
    .S(net427),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _13184_ (.A0(net1515),
    .A1(net329),
    .S(net427),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(net2428),
    .A1(net324),
    .S(net429),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _13186_ (.A0(net1720),
    .A1(net320),
    .S(net428),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _13187_ (.A0(net1711),
    .A1(net318),
    .S(net428),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _13188_ (.A0(net1860),
    .A1(net312),
    .S(net429),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _13189_ (.A0(net1604),
    .A1(net308),
    .S(net428),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(net2369),
    .A1(net305),
    .S(net429),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _13191_ (.A0(net2154),
    .A1(net303),
    .S(net430),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _13192_ (.A0(net2303),
    .A1(net300),
    .S(net429),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _13193_ (.A0(net2158),
    .A1(net295),
    .S(net429),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(net2246),
    .A1(net290),
    .S(net430),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _13195_ (.A0(net1936),
    .A1(net287),
    .S(net429),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _13196_ (.A0(net1981),
    .A1(net282),
    .S(net430),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _13197_ (.A0(net2048),
    .A1(net281),
    .S(net430),
    .X(_01830_));
 sky130_fd_sc_hd__nor2_1 _13198_ (.A(net569),
    .B(_05168_),
    .Y(_02130_));
 sky130_fd_sc_hd__a21oi_1 _13199_ (.A1(net1051),
    .A2(\decoded_imm[0] ),
    .B1(net961),
    .Y(_02131_));
 sky130_fd_sc_hd__o21a_1 _13200_ (.A1(net1051),
    .A2(\decoded_imm[0] ),
    .B1(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__and2_2 _13201_ (.A(net1063),
    .B(_02474_),
    .X(_02133_));
 sky130_fd_sc_hd__a22o_1 _13202_ (.A1(net1042),
    .A2(net709),
    .B1(net557),
    .B2(net1047),
    .X(_02134_));
 sky130_fd_sc_hd__a211o_1 _13203_ (.A1(net755),
    .A2(_02134_),
    .B1(_02132_),
    .C1(net393),
    .X(_02135_));
 sky130_fd_sc_hd__o22a_1 _13204_ (.A1(net1051),
    .A2(net397),
    .B1(_02130_),
    .B2(_02135_),
    .X(_01831_));
 sky130_fd_sc_hd__nor2_1 _13205_ (.A(net569),
    .B(_05203_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _13206_ (.A(_02384_),
    .B(net759),
    .Y(_02137_));
 sky130_fd_sc_hd__or2_1 _13207_ (.A(net1045),
    .B(net759),
    .X(_02138_));
 sky130_fd_sc_hd__a21o_1 _13208_ (.A1(_02137_),
    .A2(_02138_),
    .B1(_02475_),
    .X(_02139_));
 sky130_fd_sc_hd__a31o_1 _13209_ (.A1(net1065),
    .A2(net1040),
    .A3(net755),
    .B1(net557),
    .X(_02140_));
 sky130_fd_sc_hd__a22o_1 _13210_ (.A1(net1051),
    .A2(\decoded_imm[0] ),
    .B1(_04951_),
    .B2(_04952_),
    .X(_02141_));
 sky130_fd_sc_hd__and3_1 _13211_ (.A(net958),
    .B(_04953_),
    .C(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__a221o_1 _13212_ (.A1(\reg_pc[1] ),
    .A2(net565),
    .B1(_02139_),
    .B2(_02140_),
    .C1(net392),
    .X(_02143_));
 sky130_fd_sc_hd__o32a_1 _13213_ (.A1(_02136_),
    .A2(_02142_),
    .A3(_02143_),
    .B1(net397),
    .B2(net1047),
    .X(_01832_));
 sky130_fd_sc_hd__and2b_1 _13214_ (.A_N(net569),
    .B(_03189_),
    .X(_02144_));
 sky130_fd_sc_hd__a21o_1 _13215_ (.A1(_04949_),
    .A2(_04955_),
    .B1(_04954_),
    .X(_02145_));
 sky130_fd_sc_hd__and3_1 _13216_ (.A(net959),
    .B(_04956_),
    .C(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(_02383_),
    .A1(_02402_),
    .S(net755),
    .X(_02147_));
 sky130_fd_sc_hd__nand2_1 _13218_ (.A(_02474_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__a31o_1 _13219_ (.A1(net1063),
    .A2(net1038),
    .A3(net754),
    .B1(net557),
    .X(_02149_));
 sky130_fd_sc_hd__a221o_1 _13220_ (.A1(\reg_pc[2] ),
    .A2(net565),
    .B1(_02148_),
    .B2(_02149_),
    .C1(net392),
    .X(_02150_));
 sky130_fd_sc_hd__o32a_1 _13221_ (.A1(_02144_),
    .A2(_02146_),
    .A3(_02150_),
    .B1(net397),
    .B2(net1045),
    .X(_01833_));
 sky130_fd_sc_hd__nor2_1 _13222_ (.A(_03227_),
    .B(net568),
    .Y(_02151_));
 sky130_fd_sc_hd__o211a_1 _13223_ (.A1(_04948_),
    .A2(_04957_),
    .B1(_04956_),
    .C1(_04949_),
    .X(_02152_));
 sky130_fd_sc_hd__nor3_1 _13224_ (.A(net960),
    .B(_04958_),
    .C(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(net1045),
    .A1(net1042),
    .S(net757),
    .X(_02154_));
 sky130_fd_sc_hd__or2_1 _13226_ (.A(_02475_),
    .B(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__a31o_1 _13227_ (.A1(net1063),
    .A2(net1035),
    .A3(net754),
    .B1(net557),
    .X(_02156_));
 sky130_fd_sc_hd__a221o_1 _13228_ (.A1(\reg_pc[3] ),
    .A2(net565),
    .B1(_02155_),
    .B2(_02156_),
    .C1(net392),
    .X(_02157_));
 sky130_fd_sc_hd__o32a_1 _13229_ (.A1(_02151_),
    .A2(_02153_),
    .A3(_02157_),
    .B1(net396),
    .B2(net1044),
    .X(_01834_));
 sky130_fd_sc_hd__nor2_1 _13230_ (.A(_03263_),
    .B(net568),
    .Y(_02158_));
 sky130_fd_sc_hd__a211o_1 _13231_ (.A1(_04947_),
    .A2(_04959_),
    .B1(_04958_),
    .C1(_04948_),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _13232_ (.A0(net1044),
    .A1(net1040),
    .S(net755),
    .X(_02160_));
 sky130_fd_sc_hd__or2_1 _13233_ (.A(net1033),
    .B(net758),
    .X(_02161_));
 sky130_fd_sc_hd__a221o_1 _13234_ (.A1(\reg_pc[4] ),
    .A2(net565),
    .B1(net557),
    .B2(_02160_),
    .C1(net392),
    .X(_02162_));
 sky130_fd_sc_hd__a31o_1 _13235_ (.A1(net709),
    .A2(_02137_),
    .A3(_02161_),
    .B1(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__a31o_1 _13236_ (.A1(net959),
    .A2(_04960_),
    .A3(_02159_),
    .B1(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__o22a_1 _13237_ (.A1(net1042),
    .A2(net396),
    .B1(_02158_),
    .B2(_02164_),
    .X(_01835_));
 sky130_fd_sc_hd__xnor2_1 _13238_ (.A(_04961_),
    .B(_04968_),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_1 _13239_ (.A(_02403_),
    .B(net753),
    .Y(_02166_));
 sky130_fd_sc_hd__o211a_1 _13240_ (.A1(net1047),
    .A2(net754),
    .B1(_02166_),
    .C1(net709),
    .X(_02167_));
 sky130_fd_sc_hd__or2_1 _13241_ (.A(net1042),
    .B(net753),
    .X(_02168_));
 sky130_fd_sc_hd__o2111a_1 _13242_ (.A1(net1038),
    .A2(net758),
    .B1(_02168_),
    .C1(_02474_),
    .D1(net1063),
    .X(_02169_));
 sky130_fd_sc_hd__a2111oi_1 _13243_ (.A1(\reg_pc[5] ),
    .A2(net565),
    .B1(_02167_),
    .C1(_02169_),
    .D1(net391),
    .Y(_02170_));
 sky130_fd_sc_hd__o221a_1 _13244_ (.A1(net568),
    .A2(_05242_),
    .B1(_02165_),
    .B2(net960),
    .C1(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__o21ba_1 _13245_ (.A1(net1040),
    .A2(net396),
    .B1_N(_02171_),
    .X(_01836_));
 sky130_fd_sc_hd__xnor2_1 _13246_ (.A(_04943_),
    .B(_04962_),
    .Y(_02172_));
 sky130_fd_sc_hd__or2_1 _13247_ (.A(net1040),
    .B(net752),
    .X(_02173_));
 sky130_fd_sc_hd__o2111a_1 _13248_ (.A1(net1035),
    .A2(net758),
    .B1(_02173_),
    .C1(_02474_),
    .D1(net1064),
    .X(_02174_));
 sky130_fd_sc_hd__or2_1 _13249_ (.A(net1029),
    .B(net758),
    .X(_02175_));
 sky130_fd_sc_hd__o211a_1 _13250_ (.A1(net1045),
    .A2(net754),
    .B1(_02175_),
    .C1(net709),
    .X(_02176_));
 sky130_fd_sc_hd__a2111oi_1 _13251_ (.A1(\reg_pc[6] ),
    .A2(net565),
    .B1(_02174_),
    .C1(_02176_),
    .D1(net392),
    .Y(_02177_));
 sky130_fd_sc_hd__o221a_1 _13252_ (.A1(net568),
    .A2(_05278_),
    .B1(_02172_),
    .B2(net960),
    .C1(_02177_),
    .X(_02178_));
 sky130_fd_sc_hd__o21ba_1 _13253_ (.A1(net1038),
    .A2(net396),
    .B1_N(_02178_),
    .X(_01837_));
 sky130_fd_sc_hd__xnor2_1 _13254_ (.A(_04963_),
    .B(_04965_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_1 _13255_ (.A(net960),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _13256_ (.A(net567),
    .B(_05316_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _13257_ (.A(_02404_),
    .B(net753),
    .Y(_02182_));
 sky130_fd_sc_hd__o211a_1 _13258_ (.A1(net1044),
    .A2(net753),
    .B1(_02182_),
    .C1(net708),
    .X(_02183_));
 sky130_fd_sc_hd__o211a_1 _13259_ (.A1(net1038),
    .A2(net753),
    .B1(net556),
    .C1(_02161_),
    .X(_02184_));
 sky130_fd_sc_hd__a2111o_1 _13260_ (.A1(\reg_pc[7] ),
    .A2(net564),
    .B1(_02183_),
    .C1(_02184_),
    .D1(net391),
    .X(_02185_));
 sky130_fd_sc_hd__o32a_1 _13261_ (.A1(_02180_),
    .A2(_02181_),
    .A3(_02185_),
    .B1(net395),
    .B2(net1035),
    .X(_01838_));
 sky130_fd_sc_hd__a221o_1 _13262_ (.A1(_04940_),
    .A2(_04963_),
    .B1(_04971_),
    .B2(_04936_),
    .C1(_04937_),
    .X(_02186_));
 sky130_fd_sc_hd__and3_1 _13263_ (.A(net959),
    .B(_04973_),
    .C(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__nor2_1 _13264_ (.A(net567),
    .B(_05351_),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _13265_ (.A(_02405_),
    .B(net752),
    .Y(_02189_));
 sky130_fd_sc_hd__or2_1 _13266_ (.A(net1035),
    .B(net752),
    .X(_02190_));
 sky130_fd_sc_hd__a32o_1 _13267_ (.A1(net556),
    .A2(_02166_),
    .A3(_02190_),
    .B1(net564),
    .B2(\reg_pc[8] ),
    .X(_02191_));
 sky130_fd_sc_hd__a311o_1 _13268_ (.A1(net708),
    .A2(_02168_),
    .A3(_02189_),
    .B1(_02191_),
    .C1(net391),
    .X(_02192_));
 sky130_fd_sc_hd__o32a_1 _13269_ (.A1(_02187_),
    .A2(_02188_),
    .A3(_02192_),
    .B1(net395),
    .B2(net1033),
    .X(_01839_));
 sky130_fd_sc_hd__o21ai_1 _13270_ (.A1(_04974_),
    .A2(_04981_),
    .B1(net959),
    .Y(_02193_));
 sky130_fd_sc_hd__a21oi_1 _13271_ (.A1(_04974_),
    .A2(_04981_),
    .B1(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__nor2_1 _13272_ (.A(net567),
    .B(_05386_),
    .Y(_02195_));
 sky130_fd_sc_hd__or2_1 _13273_ (.A(net1033),
    .B(net752),
    .X(_02196_));
 sky130_fd_sc_hd__nand2_1 _13274_ (.A(_02406_),
    .B(net752),
    .Y(_02197_));
 sky130_fd_sc_hd__a32o_1 _13275_ (.A1(net708),
    .A2(_02173_),
    .A3(_02197_),
    .B1(net564),
    .B2(\reg_pc[9] ),
    .X(_02198_));
 sky130_fd_sc_hd__a311o_1 _13276_ (.A1(net556),
    .A2(_02175_),
    .A3(_02196_),
    .B1(_02198_),
    .C1(net391),
    .X(_02199_));
 sky130_fd_sc_hd__o32a_1 _13277_ (.A1(_02194_),
    .A2(_02195_),
    .A3(_02199_),
    .B1(net395),
    .B2(net1032),
    .X(_01840_));
 sky130_fd_sc_hd__nand2_1 _13278_ (.A(_04933_),
    .B(_04975_),
    .Y(_02200_));
 sky130_fd_sc_hd__and3_1 _13279_ (.A(net959),
    .B(_04976_),
    .C(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__nor2_1 _13280_ (.A(net567),
    .B(_05421_),
    .Y(_02202_));
 sky130_fd_sc_hd__o211a_1 _13281_ (.A1(net1031),
    .A2(net753),
    .B1(net556),
    .C1(_02182_),
    .X(_02203_));
 sky130_fd_sc_hd__or2_1 _13282_ (.A(net1022),
    .B(net758),
    .X(_02204_));
 sky130_fd_sc_hd__o211a_1 _13283_ (.A1(net1038),
    .A2(net752),
    .B1(_02204_),
    .C1(net708),
    .X(_02205_));
 sky130_fd_sc_hd__a2111o_1 _13284_ (.A1(\reg_pc[10] ),
    .A2(net564),
    .B1(_02203_),
    .C1(_02205_),
    .D1(net391),
    .X(_02206_));
 sky130_fd_sc_hd__o32a_1 _13285_ (.A1(_02201_),
    .A2(_02202_),
    .A3(_02206_),
    .B1(net395),
    .B2(net1029),
    .X(_01841_));
 sky130_fd_sc_hd__xor2_1 _13286_ (.A(_04977_),
    .B(_04979_),
    .X(_02207_));
 sky130_fd_sc_hd__nor2_1 _13287_ (.A(net960),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__nor2_1 _13288_ (.A(net567),
    .B(_05456_),
    .Y(_02209_));
 sky130_fd_sc_hd__or2_1 _13289_ (.A(net1029),
    .B(net752),
    .X(_02210_));
 sky130_fd_sc_hd__or2_1 _13290_ (.A(net1020),
    .B(net758),
    .X(_02211_));
 sky130_fd_sc_hd__a32o_1 _13291_ (.A1(net708),
    .A2(_02190_),
    .A3(_02211_),
    .B1(net564),
    .B2(\reg_pc[11] ),
    .X(_02212_));
 sky130_fd_sc_hd__a311o_1 _13292_ (.A1(net556),
    .A2(_02189_),
    .A3(_02210_),
    .B1(_02212_),
    .C1(net391),
    .X(_02213_));
 sky130_fd_sc_hd__o32a_1 _13293_ (.A1(_02208_),
    .A2(_02209_),
    .A3(_02213_),
    .B1(net395),
    .B2(net205),
    .X(_01842_));
 sky130_fd_sc_hd__and3_1 _13294_ (.A(_04928_),
    .B(_04978_),
    .C(_04982_),
    .X(_02214_));
 sky130_fd_sc_hd__nor3_1 _13295_ (.A(net960),
    .B(_04983_),
    .C(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _13296_ (.A(net567),
    .B(_05491_),
    .Y(_02216_));
 sky130_fd_sc_hd__nand2_1 _13297_ (.A(_02404_),
    .B(net758),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _13298_ (.A(_02407_),
    .B(net753),
    .Y(_02218_));
 sky130_fd_sc_hd__a32o_1 _13299_ (.A1(net708),
    .A2(_02196_),
    .A3(_02218_),
    .B1(net564),
    .B2(\reg_pc[12] ),
    .X(_02219_));
 sky130_fd_sc_hd__a311o_1 _13300_ (.A1(net556),
    .A2(_02197_),
    .A3(_02217_),
    .B1(_02219_),
    .C1(net391),
    .X(_02220_));
 sky130_fd_sc_hd__o32a_1 _13301_ (.A1(_02215_),
    .A2(_02216_),
    .A3(_02220_),
    .B1(net395),
    .B2(net1027),
    .X(_01843_));
 sky130_fd_sc_hd__a21o_1 _13302_ (.A1(\decoded_imm[12] ),
    .A2(net1026),
    .B1(_04983_),
    .X(_02221_));
 sky130_fd_sc_hd__xnor2_1 _13303_ (.A(_04927_),
    .B(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__nand2_1 _13304_ (.A(_02408_),
    .B(net754),
    .Y(_02223_));
 sky130_fd_sc_hd__o211a_1 _13305_ (.A1(net1031),
    .A2(net752),
    .B1(_02223_),
    .C1(net708),
    .X(_02224_));
 sky130_fd_sc_hd__nand2_1 _13306_ (.A(_02405_),
    .B(net758),
    .Y(_02225_));
 sky130_fd_sc_hd__and3_1 _13307_ (.A(net556),
    .B(_02204_),
    .C(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__a211o_1 _13308_ (.A1(\reg_pc[13] ),
    .A2(net564),
    .B1(_02224_),
    .C1(net391),
    .X(_02227_));
 sky130_fd_sc_hd__a2bb2o_1 _13309_ (.A1_N(net567),
    .A2_N(_05527_),
    .B1(_02222_),
    .B2(net959),
    .X(_02228_));
 sky130_fd_sc_hd__o32a_1 _13310_ (.A1(_02226_),
    .A2(_02227_),
    .A3(_02228_),
    .B1(net395),
    .B2(net1024),
    .X(_01844_));
 sky130_fd_sc_hd__a21oi_1 _13311_ (.A1(_04922_),
    .A2(_04984_),
    .B1(net960),
    .Y(_02229_));
 sky130_fd_sc_hd__o21a_1 _13312_ (.A1(_04922_),
    .A2(_04984_),
    .B1(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__nor2_1 _13313_ (.A(net567),
    .B(_05563_),
    .Y(_02231_));
 sky130_fd_sc_hd__nand2_1 _13314_ (.A(_02406_),
    .B(net758),
    .Y(_02232_));
 sky130_fd_sc_hd__or2_1 _13315_ (.A(net1014),
    .B(net758),
    .X(_02233_));
 sky130_fd_sc_hd__a32o_1 _13316_ (.A1(net708),
    .A2(_02210_),
    .A3(_02233_),
    .B1(net564),
    .B2(\reg_pc[14] ),
    .X(_02234_));
 sky130_fd_sc_hd__a311o_1 _13317_ (.A1(net556),
    .A2(_02211_),
    .A3(_02232_),
    .B1(_02234_),
    .C1(net391),
    .X(_02235_));
 sky130_fd_sc_hd__o32a_1 _13318_ (.A1(_02230_),
    .A2(_02231_),
    .A3(_02235_),
    .B1(net395),
    .B2(net1022),
    .X(_01845_));
 sky130_fd_sc_hd__o21ai_1 _13319_ (.A1(_04922_),
    .A2(_04984_),
    .B1(_04917_),
    .Y(_02236_));
 sky130_fd_sc_hd__xnor2_1 _13320_ (.A(_04920_),
    .B(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__nor2_1 _13321_ (.A(net960),
    .B(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__nand2_1 _13322_ (.A(_02409_),
    .B(net754),
    .Y(_02239_));
 sky130_fd_sc_hd__or2_1 _13323_ (.A(net1022),
    .B(net752),
    .X(_02240_));
 sky130_fd_sc_hd__a32o_1 _13324_ (.A1(net556),
    .A2(_02218_),
    .A3(_02240_),
    .B1(net564),
    .B2(\reg_pc[15] ),
    .X(_02241_));
 sky130_fd_sc_hd__a31o_1 _13325_ (.A1(net708),
    .A2(_02217_),
    .A3(_02239_),
    .B1(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__o21ai_1 _13326_ (.A1(net567),
    .A2(_05599_),
    .B1(net395),
    .Y(_02243_));
 sky130_fd_sc_hd__o32a_1 _13327_ (.A1(_02238_),
    .A2(_02242_),
    .A3(_02243_),
    .B1(net395),
    .B2(net1020),
    .X(_01846_));
 sky130_fd_sc_hd__and3_1 _13328_ (.A(_04987_),
    .B(_04989_),
    .C(_04990_),
    .X(_02244_));
 sky130_fd_sc_hd__nor3_1 _13329_ (.A(net960),
    .B(_04991_),
    .C(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _13330_ (.A(net567),
    .B(_05637_),
    .Y(_02246_));
 sky130_fd_sc_hd__or2_1 _13331_ (.A(net1010),
    .B(net759),
    .X(_02247_));
 sky130_fd_sc_hd__or2_1 _13332_ (.A(net1020),
    .B(net754),
    .X(_02248_));
 sky130_fd_sc_hd__a32o_1 _13333_ (.A1(net557),
    .A2(_02223_),
    .A3(_02248_),
    .B1(net564),
    .B2(\reg_pc[16] ),
    .X(_02249_));
 sky130_fd_sc_hd__a311o_1 _13334_ (.A1(net708),
    .A2(_02225_),
    .A3(_02247_),
    .B1(_02249_),
    .C1(net391),
    .X(_02250_));
 sky130_fd_sc_hd__o32a_1 _13335_ (.A1(_02245_),
    .A2(_02246_),
    .A3(_02250_),
    .B1(net396),
    .B2(net1018),
    .X(_01847_));
 sky130_fd_sc_hd__a21oi_1 _13336_ (.A1(_04992_),
    .A2(_04994_),
    .B1(net960),
    .Y(_02251_));
 sky130_fd_sc_hd__o21a_1 _13337_ (.A1(_04992_),
    .A2(_04994_),
    .B1(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__nor2_1 _13338_ (.A(net568),
    .B(_05675_),
    .Y(_02253_));
 sky130_fd_sc_hd__o211a_1 _13339_ (.A1(net1018),
    .A2(net752),
    .B1(net556),
    .C1(_02233_),
    .X(_02254_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_02410_),
    .B(net755),
    .Y(_02255_));
 sky130_fd_sc_hd__a32o_1 _13341_ (.A1(net709),
    .A2(_02232_),
    .A3(_02255_),
    .B1(net565),
    .B2(\reg_pc[17] ),
    .X(_02256_));
 sky130_fd_sc_hd__or4_1 _13342_ (.A(net392),
    .B(_02253_),
    .C(_02254_),
    .D(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__o22a_1 _13343_ (.A1(net1017),
    .A2(net396),
    .B1(_02252_),
    .B2(_02257_),
    .X(_01848_));
 sky130_fd_sc_hd__or3_1 _13344_ (.A(_04996_),
    .B(_05000_),
    .C(_05004_),
    .X(_02258_));
 sky130_fd_sc_hd__o21ai_1 _13345_ (.A1(_05000_),
    .A2(_05004_),
    .B1(_04996_),
    .Y(_02259_));
 sky130_fd_sc_hd__and3_1 _13346_ (.A(net959),
    .B(_02258_),
    .C(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__nor2_1 _13347_ (.A(net568),
    .B(_05710_),
    .Y(_02261_));
 sky130_fd_sc_hd__or2_1 _13348_ (.A(net1007),
    .B(net759),
    .X(_02262_));
 sky130_fd_sc_hd__nand2_1 _13349_ (.A(_02408_),
    .B(net759),
    .Y(_02263_));
 sky130_fd_sc_hd__a32o_1 _13350_ (.A1(net557),
    .A2(_02239_),
    .A3(_02263_),
    .B1(net565),
    .B2(\reg_pc[18] ),
    .X(_02264_));
 sky130_fd_sc_hd__a311o_1 _13351_ (.A1(net709),
    .A2(_02240_),
    .A3(_02262_),
    .B1(_02264_),
    .C1(net392),
    .X(_02265_));
 sky130_fd_sc_hd__o32a_1 _13352_ (.A1(_02260_),
    .A2(_02261_),
    .A3(_02265_),
    .B1(net396),
    .B2(net1014),
    .X(_01849_));
 sky130_fd_sc_hd__a211o_1 _13353_ (.A1(_05001_),
    .A2(_02258_),
    .B1(_04998_),
    .C1(_04999_),
    .X(_02266_));
 sky130_fd_sc_hd__o211ai_1 _13354_ (.A1(_04998_),
    .A2(_04999_),
    .B1(_05001_),
    .C1(_02258_),
    .Y(_02267_));
 sky130_fd_sc_hd__and3_1 _13355_ (.A(net959),
    .B(_02266_),
    .C(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__nor2_1 _13356_ (.A(net569),
    .B(_05748_),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _13357_ (.A(_02411_),
    .B(net755),
    .Y(_02270_));
 sky130_fd_sc_hd__or2_1 _13358_ (.A(net1014),
    .B(net755),
    .X(_02271_));
 sky130_fd_sc_hd__a32o_1 _13359_ (.A1(net557),
    .A2(_02247_),
    .A3(_02271_),
    .B1(net565),
    .B2(\reg_pc[19] ),
    .X(_02272_));
 sky130_fd_sc_hd__a311o_1 _13360_ (.A1(net709),
    .A2(_02248_),
    .A3(_02270_),
    .B1(_02272_),
    .C1(net392),
    .X(_02273_));
 sky130_fd_sc_hd__o32a_1 _13361_ (.A1(_02268_),
    .A2(_02269_),
    .A3(_02273_),
    .B1(net397),
    .B2(net1012),
    .X(_01850_));
 sky130_fd_sc_hd__o21ai_1 _13362_ (.A1(_05003_),
    .A2(_05005_),
    .B1(_05007_),
    .Y(_02274_));
 sky130_fd_sc_hd__and3_1 _13363_ (.A(net958),
    .B(_05008_),
    .C(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__nor2_1 _13364_ (.A(net569),
    .B(_05784_),
    .Y(_02276_));
 sky130_fd_sc_hd__or2_1 _13365_ (.A(net1004),
    .B(net760),
    .X(_02277_));
 sky130_fd_sc_hd__o211a_1 _13366_ (.A1(net1019),
    .A2(net755),
    .B1(_02277_),
    .C1(net710),
    .X(_02278_));
 sky130_fd_sc_hd__o211a_1 _13367_ (.A1(net1012),
    .A2(net755),
    .B1(net558),
    .C1(_02255_),
    .X(_02279_));
 sky130_fd_sc_hd__a2111o_1 _13368_ (.A1(\reg_pc[20] ),
    .A2(net566),
    .B1(_02278_),
    .C1(_02279_),
    .D1(net393),
    .X(_02280_));
 sky130_fd_sc_hd__o32a_1 _13369_ (.A1(_02275_),
    .A2(_02276_),
    .A3(_02280_),
    .B1(net397),
    .B2(net1010),
    .X(_01851_));
 sky130_fd_sc_hd__a21oi_1 _13370_ (.A1(_05009_),
    .A2(_05018_),
    .B1(net961),
    .Y(_02281_));
 sky130_fd_sc_hd__o21a_1 _13371_ (.A1(_05009_),
    .A2(_05018_),
    .B1(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__nor2_1 _13372_ (.A(net569),
    .B(_05820_),
    .Y(_02283_));
 sky130_fd_sc_hd__or2_1 _13373_ (.A(net1010),
    .B(net756),
    .X(_02284_));
 sky130_fd_sc_hd__or2_1 _13374_ (.A(net1002),
    .B(net760),
    .X(_02285_));
 sky130_fd_sc_hd__a32o_1 _13375_ (.A1(net710),
    .A2(_02263_),
    .A3(_02285_),
    .B1(net566),
    .B2(\reg_pc[21] ),
    .X(_02286_));
 sky130_fd_sc_hd__a311o_1 _13376_ (.A1(net558),
    .A2(_02262_),
    .A3(_02284_),
    .B1(_02286_),
    .C1(net393),
    .X(_02287_));
 sky130_fd_sc_hd__o32a_1 _13377_ (.A1(_02282_),
    .A2(_02283_),
    .A3(_02287_),
    .B1(net397),
    .B2(net2556),
    .X(_01852_));
 sky130_fd_sc_hd__nand2_1 _13378_ (.A(_04910_),
    .B(_05011_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2_1 _13379_ (.A(_02410_),
    .B(net760),
    .Y(_02289_));
 sky130_fd_sc_hd__or2_1 _13380_ (.A(net1000),
    .B(net760),
    .X(_02290_));
 sky130_fd_sc_hd__a31o_1 _13381_ (.A1(net710),
    .A2(_02271_),
    .A3(_02290_),
    .B1(_04879_),
    .X(_02291_));
 sky130_fd_sc_hd__a31o_1 _13382_ (.A1(net558),
    .A2(_02270_),
    .A3(_02289_),
    .B1(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__a31o_1 _13383_ (.A1(net958),
    .A2(_05012_),
    .A3(_02288_),
    .B1(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__o2bb2a_1 _13384_ (.A1_N(\reg_pc[22] ),
    .A2_N(_05079_),
    .B1(_05855_),
    .B2(is_lui_auipc_jal),
    .X(_02294_));
 sky130_fd_sc_hd__a21oi_1 _13385_ (.A1(_04879_),
    .A2(_02294_),
    .B1(net393),
    .Y(_02295_));
 sky130_fd_sc_hd__a22o_1 _13386_ (.A1(net1007),
    .A2(net393),
    .B1(_02293_),
    .B2(_02295_),
    .X(_01853_));
 sky130_fd_sc_hd__xor2_1 _13387_ (.A(_05013_),
    .B(_05015_),
    .X(_02296_));
 sky130_fd_sc_hd__nor2_1 _13388_ (.A(net961),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _13389_ (.A(net569),
    .B(_05890_),
    .Y(_02298_));
 sky130_fd_sc_hd__or2_1 _13390_ (.A(net998),
    .B(_04884_),
    .X(_02299_));
 sky130_fd_sc_hd__o211a_1 _13391_ (.A1(net1012),
    .A2(net756),
    .B1(_02299_),
    .C1(net710),
    .X(_02300_));
 sky130_fd_sc_hd__or2_1 _13392_ (.A(net1007),
    .B(net756),
    .X(_02301_));
 sky130_fd_sc_hd__a32o_1 _13393_ (.A1(net558),
    .A2(_02277_),
    .A3(_02301_),
    .B1(net566),
    .B2(\reg_pc[23] ),
    .X(_02302_));
 sky130_fd_sc_hd__or4_1 _13394_ (.A(net393),
    .B(_02298_),
    .C(_02300_),
    .D(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__o22a_1 _13395_ (.A1(net2764),
    .A2(net397),
    .B1(_02297_),
    .B2(_02303_),
    .X(_01854_));
 sky130_fd_sc_hd__o21ai_1 _13396_ (.A1(_05021_),
    .A2(_05023_),
    .B1(net959),
    .Y(_02304_));
 sky130_fd_sc_hd__a21oi_1 _13397_ (.A1(_05021_),
    .A2(_05023_),
    .B1(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _13398_ (.A(net569),
    .B(_05926_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand2_1 _13399_ (.A(_02412_),
    .B(net756),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_1 _13400_ (.A(_02411_),
    .B(net760),
    .Y(_02308_));
 sky130_fd_sc_hd__a32o_1 _13401_ (.A1(net558),
    .A2(_02285_),
    .A3(_02308_),
    .B1(net566),
    .B2(\reg_pc[24] ),
    .X(_02309_));
 sky130_fd_sc_hd__a311o_1 _13402_ (.A1(_02501_),
    .A2(_02284_),
    .A3(_02307_),
    .B1(_02309_),
    .C1(net394),
    .X(_02310_));
 sky130_fd_sc_hd__o32a_1 _13403_ (.A1(_02305_),
    .A2(_02306_),
    .A3(_02310_),
    .B1(net397),
    .B2(net1004),
    .X(_01855_));
 sky130_fd_sc_hd__o21ai_1 _13404_ (.A1(_05024_),
    .A2(_05029_),
    .B1(net958),
    .Y(_02311_));
 sky130_fd_sc_hd__a21oi_1 _13405_ (.A1(_05024_),
    .A2(_05029_),
    .B1(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _13406_ (.A(net570),
    .B(_05964_),
    .Y(_02313_));
 sky130_fd_sc_hd__o211a_1 _13407_ (.A1(net1004),
    .A2(net756),
    .B1(net558),
    .C1(_02290_),
    .X(_02314_));
 sky130_fd_sc_hd__or2_1 _13408_ (.A(net994),
    .B(net760),
    .X(_02315_));
 sky130_fd_sc_hd__a32o_1 _13409_ (.A1(net710),
    .A2(_02289_),
    .A3(_02315_),
    .B1(net566),
    .B2(\reg_pc[25] ),
    .X(_02316_));
 sky130_fd_sc_hd__or4_1 _13410_ (.A(net394),
    .B(_02313_),
    .C(_02314_),
    .D(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__o22a_1 _13411_ (.A1(net1002),
    .A2(net397),
    .B1(_02312_),
    .B2(_02317_),
    .X(_01856_));
 sky130_fd_sc_hd__o21a_1 _13412_ (.A1(_04902_),
    .A2(_05025_),
    .B1(_04900_),
    .X(_02318_));
 sky130_fd_sc_hd__nor3_1 _13413_ (.A(net961),
    .B(_05026_),
    .C(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _13414_ (.A(net569),
    .B(_05999_),
    .Y(_02320_));
 sky130_fd_sc_hd__or2_1 _13415_ (.A(net992),
    .B(net760),
    .X(_02321_));
 sky130_fd_sc_hd__or2_1 _13416_ (.A(net1002),
    .B(net757),
    .X(_02322_));
 sky130_fd_sc_hd__a32o_1 _13417_ (.A1(net558),
    .A2(_02299_),
    .A3(_02322_),
    .B1(net566),
    .B2(\reg_pc[26] ),
    .X(_02323_));
 sky130_fd_sc_hd__a311o_1 _13418_ (.A1(net710),
    .A2(_02301_),
    .A3(_02321_),
    .B1(_02323_),
    .C1(net394),
    .X(_02324_));
 sky130_fd_sc_hd__o32a_1 _13419_ (.A1(_02319_),
    .A2(_02320_),
    .A3(_02324_),
    .B1(net398),
    .B2(net1000),
    .X(_01857_));
 sky130_fd_sc_hd__a211o_1 _13420_ (.A1(_04897_),
    .A2(_05028_),
    .B1(_05026_),
    .C1(_04898_),
    .X(_02325_));
 sky130_fd_sc_hd__o211ai_1 _13421_ (.A1(_04898_),
    .A2(_05026_),
    .B1(_05028_),
    .C1(_04897_),
    .Y(_02326_));
 sky130_fd_sc_hd__or2_1 _13422_ (.A(net1000),
    .B(net756),
    .X(_02327_));
 sky130_fd_sc_hd__or2_1 _13423_ (.A(net1188),
    .B(net760),
    .X(_02328_));
 sky130_fd_sc_hd__a31o_1 _13424_ (.A1(net558),
    .A2(_02307_),
    .A3(_02327_),
    .B1(_04879_),
    .X(_02329_));
 sky130_fd_sc_hd__a31o_1 _13425_ (.A1(net710),
    .A2(_02308_),
    .A3(_02328_),
    .B1(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__a31o_1 _13426_ (.A1(_02463_),
    .A2(_02325_),
    .A3(_02326_),
    .B1(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__o2bb2a_1 _13427_ (.A1_N(\reg_pc[27] ),
    .A2_N(_05079_),
    .B1(_06034_),
    .B2(is_lui_auipc_jal),
    .X(_02332_));
 sky130_fd_sc_hd__a21oi_1 _13428_ (.A1(_04879_),
    .A2(_02332_),
    .B1(net393),
    .Y(_02333_));
 sky130_fd_sc_hd__a22o_1 _13429_ (.A1(net998),
    .A2(net393),
    .B1(_02331_),
    .B2(_02333_),
    .X(_01858_));
 sky130_fd_sc_hd__o21ai_1 _13430_ (.A1(_04896_),
    .A2(_05030_),
    .B1(net958),
    .Y(_02334_));
 sky130_fd_sc_hd__a21oi_1 _13431_ (.A1(_04896_),
    .A2(_05030_),
    .B1(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__a21o_1 _13432_ (.A1(net1188),
    .A2(_04883_),
    .B1(net760),
    .X(_02336_));
 sky130_fd_sc_hd__o211a_1 _13433_ (.A1(net1005),
    .A2(net756),
    .B1(_02336_),
    .C1(net710),
    .X(_02337_));
 sky130_fd_sc_hd__o211a_1 _13434_ (.A1(net998),
    .A2(net756),
    .B1(_02133_),
    .C1(_02315_),
    .X(_02338_));
 sky130_fd_sc_hd__nor2_1 _13435_ (.A(is_lui_auipc_jal),
    .B(_06069_),
    .Y(_02339_));
 sky130_fd_sc_hd__a211o_1 _13436_ (.A1(\reg_pc[28] ),
    .A2(_05079_),
    .B1(_02339_),
    .C1(_04880_),
    .X(_02340_));
 sky130_fd_sc_hd__o41a_1 _13437_ (.A1(_04879_),
    .A2(_02335_),
    .A3(_02337_),
    .A4(_02338_),
    .B1(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(net996),
    .A1(_02341_),
    .S(net398),
    .X(_01859_));
 sky130_fd_sc_hd__a21oi_1 _13439_ (.A1(_05031_),
    .A2(_05033_),
    .B1(net961),
    .Y(_02342_));
 sky130_fd_sc_hd__o21a_1 _13440_ (.A1(_05031_),
    .A2(_05033_),
    .B1(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__nor2_1 _13441_ (.A(net570),
    .B(_06105_),
    .Y(_02344_));
 sky130_fd_sc_hd__and3_1 _13442_ (.A(net710),
    .B(_02322_),
    .C(_02336_),
    .X(_02345_));
 sky130_fd_sc_hd__o211a_1 _13443_ (.A1(net996),
    .A2(net757),
    .B1(net558),
    .C1(_02321_),
    .X(_02346_));
 sky130_fd_sc_hd__a2111o_1 _13444_ (.A1(\reg_pc[29] ),
    .A2(net566),
    .B1(_02345_),
    .C1(_02346_),
    .D1(net393),
    .X(_02347_));
 sky130_fd_sc_hd__o32a_1 _13445_ (.A1(_02343_),
    .A2(_02344_),
    .A3(_02347_),
    .B1(net397),
    .B2(net994),
    .X(_01860_));
 sky130_fd_sc_hd__o21a_1 _13446_ (.A1(_04894_),
    .A2(_05032_),
    .B1(_04893_),
    .X(_02348_));
 sky130_fd_sc_hd__nor3_1 _13447_ (.A(net961),
    .B(_05034_),
    .C(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hd__o211a_1 _13448_ (.A1(net1000),
    .A2(net757),
    .B1(_02336_),
    .C1(_02501_),
    .X(_02350_));
 sky130_fd_sc_hd__o211a_1 _13449_ (.A1(net994),
    .A2(net756),
    .B1(net558),
    .C1(_02328_),
    .X(_02351_));
 sky130_fd_sc_hd__or4_1 _13450_ (.A(_04879_),
    .B(_02349_),
    .C(_02350_),
    .D(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__o2bb2a_1 _13451_ (.A1_N(\reg_pc[30] ),
    .A2_N(_05079_),
    .B1(_06143_),
    .B2(is_lui_auipc_jal),
    .X(_02353_));
 sky130_fd_sc_hd__a21oi_1 _13452_ (.A1(_04879_),
    .A2(_02353_),
    .B1(net394),
    .Y(_02354_));
 sky130_fd_sc_hd__a22o_1 _13453_ (.A1(net992),
    .A2(net394),
    .B1(_02352_),
    .B2(_02354_),
    .X(_01861_));
 sky130_fd_sc_hd__nor2_1 _13454_ (.A(_03745_),
    .B(_02127_),
    .Y(_02355_));
 sky130_fd_sc_hd__mux2_1 _13455_ (.A0(net1581),
    .A1(net587),
    .S(net426),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _13456_ (.A0(net1677),
    .A1(net583),
    .S(net425),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _13457_ (.A0(net1399),
    .A1(net579),
    .S(net426),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _13458_ (.A0(net1431),
    .A1(net575),
    .S(net423),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _13459_ (.A0(net1413),
    .A1(net571),
    .S(net426),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _13460_ (.A0(net1929),
    .A1(net544),
    .S(net423),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _13461_ (.A0(net1583),
    .A1(net537),
    .S(net424),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _13462_ (.A0(net1710),
    .A1(net526),
    .S(net424),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _13463_ (.A0(net1634),
    .A1(net520),
    .S(net424),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _13464_ (.A0(net1544),
    .A1(net407),
    .S(net424),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _13465_ (.A0(net1415),
    .A1(net404),
    .S(net424),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _13466_ (.A0(net2080),
    .A1(net356),
    .S(net424),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _13467_ (.A0(net1994),
    .A1(net352),
    .S(net423),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _13468_ (.A0(net1429),
    .A1(net348),
    .S(net423),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _13469_ (.A0(net1708),
    .A1(net345),
    .S(net424),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _13470_ (.A0(net1521),
    .A1(net341),
    .S(net423),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(net1694),
    .A1(net336),
    .S(net423),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _13472_ (.A0(net1595),
    .A1(net334),
    .S(net423),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(net1576),
    .A1(net329),
    .S(net423),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _13474_ (.A0(net1779),
    .A1(net324),
    .S(net425),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(net1693),
    .A1(net320),
    .S(net423),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _13476_ (.A0(net1445),
    .A1(net317),
    .S(net423),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _13477_ (.A0(net1420),
    .A1(net312),
    .S(net425),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _13478_ (.A0(net1551),
    .A1(net308),
    .S(net424),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _13479_ (.A0(net1742),
    .A1(net305),
    .S(net426),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _13480_ (.A0(net1560),
    .A1(net303),
    .S(net425),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _13481_ (.A0(net1554),
    .A1(net299),
    .S(net425),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_1 _13482_ (.A0(net1473),
    .A1(net295),
    .S(net425),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _13483_ (.A0(net1407),
    .A1(net290),
    .S(net425),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _13484_ (.A0(net1343),
    .A1(net287),
    .S(net425),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _13485_ (.A0(net1610),
    .A1(net282),
    .S(net425),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _13486_ (.A0(net1559),
    .A1(net280),
    .S(net425),
    .X(_01893_));
 sky130_fd_sc_hd__nor2_1 _13487_ (.A(_04283_),
    .B(_02127_),
    .Y(_02356_));
 sky130_fd_sc_hd__mux2_1 _13488_ (.A0(net2255),
    .A1(net586),
    .S(net422),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _13489_ (.A0(net2113),
    .A1(net583),
    .S(net421),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_1 _13490_ (.A0(net1775),
    .A1(net579),
    .S(net422),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _13491_ (.A0(net1771),
    .A1(net575),
    .S(net419),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _13492_ (.A0(net1485),
    .A1(net572),
    .S(net422),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _13493_ (.A0(net1856),
    .A1(net544),
    .S(net419),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _13494_ (.A0(net2188),
    .A1(net537),
    .S(net420),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _13495_ (.A0(net1657),
    .A1(net526),
    .S(net420),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _13496_ (.A0(net1943),
    .A1(net520),
    .S(net420),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _13497_ (.A0(net2165),
    .A1(net407),
    .S(net420),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _13498_ (.A0(net1533),
    .A1(net404),
    .S(net420),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _13499_ (.A0(net1483),
    .A1(net356),
    .S(net420),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _13500_ (.A0(net1975),
    .A1(net352),
    .S(net419),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _13501_ (.A0(net1519),
    .A1(net348),
    .S(net419),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _13502_ (.A0(net1707),
    .A1(net345),
    .S(net420),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _13503_ (.A0(net1776),
    .A1(net341),
    .S(net419),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _13504_ (.A0(net1885),
    .A1(net336),
    .S(net419),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(net1839),
    .A1(net334),
    .S(net419),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _13506_ (.A0(net1980),
    .A1(net329),
    .S(net419),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _13507_ (.A0(net1952),
    .A1(net324),
    .S(net421),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _13508_ (.A0(net1794),
    .A1(net320),
    .S(net419),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _13509_ (.A0(net1690),
    .A1(net317),
    .S(net419),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(net1855),
    .A1(net312),
    .S(net421),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _13511_ (.A0(net1678),
    .A1(net308),
    .S(net420),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _13512_ (.A0(net1947),
    .A1(net305),
    .S(net422),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _13513_ (.A0(net2013),
    .A1(net303),
    .S(net421),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _13514_ (.A0(net1726),
    .A1(net299),
    .S(net421),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_1 _13515_ (.A0(net2100),
    .A1(net295),
    .S(net421),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_1 _13516_ (.A0(net1787),
    .A1(net290),
    .S(net421),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _13517_ (.A0(net1586),
    .A1(net287),
    .S(net421),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(net1621),
    .A1(net282),
    .S(net421),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _13519_ (.A0(net2022),
    .A1(net280),
    .S(net421),
    .X(_01925_));
 sky130_fd_sc_hd__or2_4 _13520_ (.A(_03742_),
    .B(_04273_),
    .X(_02357_));
 sky130_fd_sc_hd__mux2_1 _13521_ (.A0(net587),
    .A1(net2459),
    .S(net417),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_1 _13522_ (.A0(net583),
    .A1(net1844),
    .S(net417),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _13523_ (.A0(net579),
    .A1(net1558),
    .S(net418),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(net576),
    .A1(net1661),
    .S(net415),
    .X(_01929_));
 sky130_fd_sc_hd__mux2_1 _13525_ (.A0(net574),
    .A1(net1795),
    .S(net418),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_1 _13526_ (.A0(net541),
    .A1(net2075),
    .S(net415),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _13527_ (.A0(net540),
    .A1(net1800),
    .S(net415),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(net524),
    .A1(net1722),
    .S(net416),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _13529_ (.A0(net520),
    .A1(net1443),
    .S(net416),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _13530_ (.A0(net407),
    .A1(net1870),
    .S(net416),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _13531_ (.A0(net404),
    .A1(net2019),
    .S(net416),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(net354),
    .A1(net1983),
    .S(net416),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _13533_ (.A0(net350),
    .A1(net1816),
    .S(net415),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _13534_ (.A0(net348),
    .A1(net2070),
    .S(net415),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _13535_ (.A0(net344),
    .A1(net1433),
    .S(net416),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _13536_ (.A0(net339),
    .A1(net1817),
    .S(net415),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _13537_ (.A0(net336),
    .A1(net1752),
    .S(net415),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _13538_ (.A0(net332),
    .A1(net1709),
    .S(net415),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _13539_ (.A0(net328),
    .A1(net1789),
    .S(net415),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(net324),
    .A1(net1904),
    .S(net417),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _13541_ (.A0(net320),
    .A1(net2044),
    .S(net415),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _13542_ (.A0(net316),
    .A1(net1757),
    .S(net417),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _13543_ (.A0(net312),
    .A1(net1878),
    .S(net417),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _13544_ (.A0(net310),
    .A1(net2111),
    .S(net417),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(net306),
    .A1(net2072),
    .S(net418),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _13546_ (.A0(net301),
    .A1(net1868),
    .S(net418),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _13547_ (.A0(net297),
    .A1(net1686),
    .S(net418),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _13548_ (.A0(net293),
    .A1(net2088),
    .S(net417),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _13549_ (.A0(net289),
    .A1(net2321),
    .S(net417),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _13550_ (.A0(net286),
    .A1(net2620),
    .S(net418),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _13551_ (.A0(net283),
    .A1(net2045),
    .S(net417),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _13552_ (.A0(net278),
    .A1(net2186),
    .S(net417),
    .X(_01957_));
 sky130_fd_sc_hd__or2_4 _13553_ (.A(_03742_),
    .B(_04275_),
    .X(_02358_));
 sky130_fd_sc_hd__mux2_1 _13554_ (.A0(net587),
    .A1(net2526),
    .S(net413),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _13555_ (.A0(net583),
    .A1(net2416),
    .S(net413),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _13556_ (.A0(net581),
    .A1(net2212),
    .S(net414),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _13557_ (.A0(net577),
    .A1(net2288),
    .S(net411),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(net574),
    .A1(net2436),
    .S(net414),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _13559_ (.A0(net542),
    .A1(net2417),
    .S(net411),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _13560_ (.A0(net540),
    .A1(net2439),
    .S(net411),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _13561_ (.A0(net524),
    .A1(net2396),
    .S(net412),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _13562_ (.A0(net520),
    .A1(net2232),
    .S(net412),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_1 _13563_ (.A0(net407),
    .A1(net2282),
    .S(net412),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _13564_ (.A0(net405),
    .A1(net2192),
    .S(net412),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _13565_ (.A0(net355),
    .A1(net2301),
    .S(net412),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _13566_ (.A0(net350),
    .A1(net2144),
    .S(net411),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _13567_ (.A0(net348),
    .A1(net2180),
    .S(net411),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(net343),
    .A1(net2358),
    .S(net412),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _13569_ (.A0(net339),
    .A1(net2171),
    .S(net411),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _13570_ (.A0(net336),
    .A1(net2214),
    .S(net411),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _13571_ (.A0(net332),
    .A1(net2228),
    .S(net411),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _13572_ (.A0(net328),
    .A1(net2325),
    .S(net411),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _13573_ (.A0(net324),
    .A1(net2494),
    .S(net413),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_1 _13574_ (.A0(net320),
    .A1(net2412),
    .S(net411),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _13575_ (.A0(net316),
    .A1(net2374),
    .S(net413),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(net312),
    .A1(net2407),
    .S(net413),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _13577_ (.A0(net310),
    .A1(net2230),
    .S(net413),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _13578_ (.A0(net306),
    .A1(net2359),
    .S(net414),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _13579_ (.A0(net301),
    .A1(net2272),
    .S(net414),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _13580_ (.A0(net297),
    .A1(net2251),
    .S(net414),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_1 _13581_ (.A0(net293),
    .A1(net2372),
    .S(net413),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _13582_ (.A0(net289),
    .A1(net2484),
    .S(net413),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _13583_ (.A0(net286),
    .A1(net2168),
    .S(net414),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _13584_ (.A0(net283),
    .A1(net2441),
    .S(net413),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _13585_ (.A0(net278),
    .A1(net2431),
    .S(net413),
    .X(_01989_));
 sky130_fd_sc_hd__clkbuf_1 _13586_ (.A(net1325),
    .X(_01598_));
 sky130_fd_sc_hd__clkbuf_1 _13587_ (.A(net1319),
    .X(_01599_));
 sky130_fd_sc_hd__clkbuf_1 _13588_ (.A(net1323),
    .X(_01600_));
 sky130_fd_sc_hd__clkbuf_1 _13589_ (.A(net1320),
    .X(_01601_));
 sky130_fd_sc_hd__clkbuf_1 _13590_ (.A(net1321),
    .X(_01602_));
 sky130_fd_sc_hd__clkbuf_1 _13591_ (.A(net1324),
    .X(_01603_));
 sky130_fd_sc_hd__clkbuf_1 _13592_ (.A(net1317),
    .X(_01604_));
 sky130_fd_sc_hd__clkbuf_1 _13593_ (.A(net1318),
    .X(_01605_));
 sky130_fd_sc_hd__clkbuf_1 _13594_ (.A(net1322),
    .X(_01606_));
 sky130_fd_sc_hd__dfxtp_1 _13595_ (.CLK(clknet_leaf_39_clk),
    .D(_00050_),
    .Q(\cpuregs[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13596_ (.CLK(clknet_leaf_45_clk),
    .D(_00051_),
    .Q(\cpuregs[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13597_ (.CLK(clknet_leaf_28_clk),
    .D(_00052_),
    .Q(\cpuregs[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13598_ (.CLK(clknet_leaf_21_clk),
    .D(_00053_),
    .Q(\cpuregs[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13599_ (.CLK(clknet_leaf_27_clk),
    .D(_00054_),
    .Q(\cpuregs[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13600_ (.CLK(clknet_leaf_24_clk),
    .D(_00055_),
    .Q(\cpuregs[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13601_ (.CLK(clknet_leaf_178_clk),
    .D(_00056_),
    .Q(\cpuregs[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13602_ (.CLK(clknet_leaf_192_clk),
    .D(_00057_),
    .Q(\cpuregs[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13603_ (.CLK(clknet_leaf_183_clk),
    .D(_00058_),
    .Q(\cpuregs[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13604_ (.CLK(clknet_leaf_184_clk),
    .D(_00059_),
    .Q(\cpuregs[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13605_ (.CLK(clknet_leaf_187_clk),
    .D(_00060_),
    .Q(\cpuregs[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13606_ (.CLK(clknet_leaf_191_clk),
    .D(_00061_),
    .Q(\cpuregs[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13607_ (.CLK(clknet_leaf_2_clk),
    .D(_00062_),
    .Q(\cpuregs[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13608_ (.CLK(clknet_leaf_195_clk),
    .D(_00063_),
    .Q(\cpuregs[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13609_ (.CLK(clknet_leaf_191_clk),
    .D(_00064_),
    .Q(\cpuregs[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13610_ (.CLK(clknet_leaf_199_clk),
    .D(_00065_),
    .Q(\cpuregs[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13611_ (.CLK(clknet_leaf_10_clk),
    .D(_00066_),
    .Q(\cpuregs[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13612_ (.CLK(clknet_leaf_0_clk),
    .D(_00067_),
    .Q(\cpuregs[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13613_ (.CLK(clknet_leaf_1_clk),
    .D(_00068_),
    .Q(\cpuregs[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13614_ (.CLK(clknet_leaf_42_clk),
    .D(_00069_),
    .Q(\cpuregs[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13615_ (.CLK(clknet_leaf_11_clk),
    .D(_00070_),
    .Q(\cpuregs[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13616_ (.CLK(clknet_leaf_13_clk),
    .D(_00071_),
    .Q(\cpuregs[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13617_ (.CLK(clknet_leaf_44_clk),
    .D(_00072_),
    .Q(\cpuregs[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13618_ (.CLK(clknet_leaf_23_clk),
    .D(_00073_),
    .Q(\cpuregs[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13619_ (.CLK(clknet_leaf_31_clk),
    .D(_00074_),
    .Q(\cpuregs[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13620_ (.CLK(clknet_leaf_72_clk),
    .D(_00075_),
    .Q(\cpuregs[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13621_ (.CLK(clknet_leaf_71_clk),
    .D(_00076_),
    .Q(\cpuregs[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13622_ (.CLK(clknet_leaf_49_clk),
    .D(_00077_),
    .Q(\cpuregs[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13623_ (.CLK(clknet_leaf_46_clk),
    .D(_00078_),
    .Q(\cpuregs[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13624_ (.CLK(clknet_leaf_73_clk),
    .D(_00079_),
    .Q(\cpuregs[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13625_ (.CLK(clknet_leaf_53_clk),
    .D(_00080_),
    .Q(\cpuregs[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13626_ (.CLK(clknet_leaf_49_clk),
    .D(_00081_),
    .Q(\cpuregs[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13627_ (.CLK(clknet_leaf_98_clk),
    .D(net945),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_ready ));
 sky130_fd_sc_hd__dfxtp_1 _13628_ (.CLK(clknet_leaf_102_clk),
    .D(_00082_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13629_ (.CLK(clknet_leaf_120_clk),
    .D(_00083_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13630_ (.CLK(clknet_leaf_120_clk),
    .D(_00084_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13631_ (.CLK(clknet_leaf_120_clk),
    .D(_00085_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_leaf_120_clk),
    .D(_00086_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_leaf_119_clk),
    .D(_00087_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_leaf_144_clk),
    .D(_00088_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_leaf_144_clk),
    .D(_00089_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_leaf_144_clk),
    .D(_00090_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_leaf_145_clk),
    .D(_00091_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_leaf_148_clk),
    .D(_00092_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_leaf_147_clk),
    .D(_00093_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_leaf_148_clk),
    .D(_00094_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_leaf_149_clk),
    .D(_00095_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_leaf_151_clk),
    .D(_00096_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_leaf_151_clk),
    .D(_00097_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_leaf_151_clk),
    .D(_00098_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_leaf_147_clk),
    .D(_00099_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_leaf_146_clk),
    .D(_00100_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_leaf_143_clk),
    .D(_00101_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_leaf_144_clk),
    .D(_00102_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_leaf_118_clk),
    .D(_00103_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13650_ (.CLK(clknet_leaf_116_clk),
    .D(_00104_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_leaf_116_clk),
    .D(_00105_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_leaf_116_clk),
    .D(_00106_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13653_ (.CLK(clknet_leaf_112_clk),
    .D(_00107_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13654_ (.CLK(clknet_leaf_112_clk),
    .D(_00108_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_leaf_113_clk),
    .D(_00109_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_leaf_113_clk),
    .D(_00110_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_leaf_107_clk),
    .D(_00111_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13658_ (.CLK(clknet_leaf_107_clk),
    .D(_00112_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_leaf_108_clk),
    .D(_00113_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_leaf_105_clk),
    .D(_00114_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_leaf_108_clk),
    .D(_00115_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13662_ (.CLK(clknet_leaf_116_clk),
    .D(_00116_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_leaf_120_clk),
    .D(_00117_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[33] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_leaf_119_clk),
    .D(_00118_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_leaf_119_clk),
    .D(_00119_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_leaf_118_clk),
    .D(_00120_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13667_ (.CLK(clknet_leaf_118_clk),
    .D(_00121_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13668_ (.CLK(clknet_leaf_144_clk),
    .D(_00122_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13669_ (.CLK(clknet_leaf_145_clk),
    .D(_00123_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13670_ (.CLK(clknet_leaf_148_clk),
    .D(_00124_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13671_ (.CLK(clknet_leaf_148_clk),
    .D(_00125_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13672_ (.CLK(clknet_leaf_148_clk),
    .D(_00126_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13673_ (.CLK(clknet_leaf_149_clk),
    .D(_00127_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13674_ (.CLK(clknet_leaf_150_clk),
    .D(_00128_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13675_ (.CLK(clknet_leaf_150_clk),
    .D(_00129_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13676_ (.CLK(clknet_leaf_150_clk),
    .D(_00130_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13677_ (.CLK(clknet_leaf_147_clk),
    .D(_00131_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13678_ (.CLK(clknet_leaf_146_clk),
    .D(_00132_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13679_ (.CLK(clknet_leaf_146_clk),
    .D(_00133_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13680_ (.CLK(clknet_leaf_144_clk),
    .D(_00134_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13681_ (.CLK(clknet_leaf_118_clk),
    .D(_00135_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13682_ (.CLK(clknet_leaf_117_clk),
    .D(_00136_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13683_ (.CLK(clknet_leaf_117_clk),
    .D(_00137_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13684_ (.CLK(clknet_leaf_115_clk),
    .D(_00138_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13685_ (.CLK(clknet_leaf_115_clk),
    .D(_00139_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13686_ (.CLK(clknet_leaf_114_clk),
    .D(_00140_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13687_ (.CLK(clknet_leaf_113_clk),
    .D(_00141_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13688_ (.CLK(clknet_leaf_113_clk),
    .D(_00142_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13689_ (.CLK(clknet_leaf_107_clk),
    .D(_00143_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13690_ (.CLK(clknet_leaf_106_clk),
    .D(_00144_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13691_ (.CLK(clknet_leaf_106_clk),
    .D(_00145_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13692_ (.CLK(clknet_leaf_106_clk),
    .D(_00146_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13693_ (.CLK(clknet_leaf_105_clk),
    .D(_00147_),
    .Q(\genblk1.genblk1.pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13694_ (.CLK(clknet_leaf_119_clk),
    .D(_00148_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13695_ (.CLK(clknet_leaf_147_clk),
    .D(_00149_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13696_ (.CLK(clknet_leaf_151_clk),
    .D(_00150_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13697_ (.CLK(clknet_leaf_146_clk),
    .D(_00151_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13698_ (.CLK(clknet_leaf_116_clk),
    .D(_00152_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13699_ (.CLK(clknet_leaf_112_clk),
    .D(_00153_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13700_ (.CLK(clknet_leaf_107_clk),
    .D(_00154_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13701_ (.CLK(clknet_leaf_112_clk),
    .D(_00155_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13702_ (.CLK(clknet_leaf_119_clk),
    .D(_00156_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13703_ (.CLK(clknet_leaf_147_clk),
    .D(_00157_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13704_ (.CLK(clknet_leaf_149_clk),
    .D(_00158_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13705_ (.CLK(clknet_leaf_146_clk),
    .D(_00159_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13706_ (.CLK(clknet_leaf_117_clk),
    .D(_00160_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13707_ (.CLK(clknet_leaf_115_clk),
    .D(_00161_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13708_ (.CLK(clknet_leaf_107_clk),
    .D(_00162_),
    .Q(\genblk1.genblk1.pcpi_mul.rdx[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_leaf_124_clk),
    .D(_00163_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13710_ (.CLK(clknet_leaf_120_clk),
    .D(_00164_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_leaf_120_clk),
    .D(_00165_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_leaf_122_clk),
    .D(_00166_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_leaf_119_clk),
    .D(_00167_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_leaf_121_clk),
    .D(_00168_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_leaf_144_clk),
    .D(_00169_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_leaf_140_clk),
    .D(_00170_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_leaf_151_clk),
    .D(_00171_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_leaf_138_clk),
    .D(_00172_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_leaf_151_clk),
    .D(_00173_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13720_ (.CLK(clknet_leaf_150_clk),
    .D(_00174_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_leaf_151_clk),
    .D(_00175_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_leaf_151_clk),
    .D(_00176_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_leaf_151_clk),
    .D(_00177_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_leaf_150_clk),
    .D(_00178_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_leaf_146_clk),
    .D(_00179_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_leaf_141_clk),
    .D(_00180_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_leaf_142_clk),
    .D(_00181_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_leaf_122_clk),
    .D(_00182_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13729_ (.CLK(clknet_leaf_116_clk),
    .D(_00183_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13730_ (.CLK(clknet_leaf_116_clk),
    .D(_00184_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13731_ (.CLK(clknet_leaf_112_clk),
    .D(_00185_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13732_ (.CLK(clknet_leaf_112_clk),
    .D(_00186_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13733_ (.CLK(clknet_leaf_112_clk),
    .D(_00187_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_leaf_113_clk),
    .D(_00188_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_leaf_113_clk),
    .D(_00189_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_leaf_107_clk),
    .D(_00190_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13737_ (.CLK(clknet_leaf_108_clk),
    .D(_00191_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_leaf_108_clk),
    .D(_00192_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13739_ (.CLK(clknet_leaf_105_clk),
    .D(_00193_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13740_ (.CLK(clknet_leaf_108_clk),
    .D(_00194_),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_rd[31] ));
 sky130_fd_sc_hd__dfxtp_4 _13741_ (.CLK(clknet_leaf_105_clk),
    .D(net2516),
    .Q(\genblk1.genblk1.pcpi_mul.mul_waiting ));
 sky130_fd_sc_hd__dfxtp_1 _13742_ (.CLK(clknet_leaf_36_clk),
    .D(_00196_),
    .Q(\cpuregs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13743_ (.CLK(clknet_leaf_44_clk),
    .D(_00197_),
    .Q(\cpuregs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13744_ (.CLK(clknet_leaf_31_clk),
    .D(_00198_),
    .Q(\cpuregs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13745_ (.CLK(clknet_leaf_17_clk),
    .D(_00199_),
    .Q(\cpuregs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13746_ (.CLK(clknet_leaf_29_clk),
    .D(_00200_),
    .Q(\cpuregs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13747_ (.CLK(clknet_leaf_21_clk),
    .D(_00201_),
    .Q(\cpuregs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13748_ (.CLK(clknet_leaf_21_clk),
    .D(_00202_),
    .Q(\cpuregs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13749_ (.CLK(clknet_leaf_19_clk),
    .D(_00203_),
    .Q(\cpuregs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13750_ (.CLK(clknet_leaf_182_clk),
    .D(_00204_),
    .Q(\cpuregs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13751_ (.CLK(clknet_leaf_181_clk),
    .D(_00205_),
    .Q(\cpuregs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13752_ (.CLK(clknet_leaf_193_clk),
    .D(_00206_),
    .Q(\cpuregs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13753_ (.CLK(clknet_leaf_194_clk),
    .D(_00207_),
    .Q(\cpuregs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13754_ (.CLK(clknet_leaf_3_clk),
    .D(_00208_),
    .Q(\cpuregs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13755_ (.CLK(clknet_leaf_4_clk),
    .D(_00209_),
    .Q(\cpuregs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13756_ (.CLK(clknet_leaf_4_clk),
    .D(_00210_),
    .Q(\cpuregs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13757_ (.CLK(clknet_leaf_1_clk),
    .D(_00211_),
    .Q(\cpuregs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13758_ (.CLK(clknet_leaf_11_clk),
    .D(_00212_),
    .Q(\cpuregs[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13759_ (.CLK(clknet_leaf_9_clk),
    .D(_00213_),
    .Q(\cpuregs[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13760_ (.CLK(clknet_leaf_8_clk),
    .D(_00214_),
    .Q(\cpuregs[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13761_ (.CLK(clknet_leaf_41_clk),
    .D(_00215_),
    .Q(\cpuregs[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13762_ (.CLK(clknet_leaf_14_clk),
    .D(_00216_),
    .Q(\cpuregs[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13763_ (.CLK(clknet_leaf_15_clk),
    .D(_00217_),
    .Q(\cpuregs[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13764_ (.CLK(clknet_leaf_40_clk),
    .D(_00218_),
    .Q(\cpuregs[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13765_ (.CLK(clknet_leaf_16_clk),
    .D(_00219_),
    .Q(\cpuregs[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13766_ (.CLK(clknet_leaf_35_clk),
    .D(_00220_),
    .Q(\cpuregs[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13767_ (.CLK(clknet_leaf_57_clk),
    .D(_00221_),
    .Q(\cpuregs[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13768_ (.CLK(clknet_leaf_57_clk),
    .D(_00222_),
    .Q(\cpuregs[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13769_ (.CLK(clknet_leaf_52_clk),
    .D(_00223_),
    .Q(\cpuregs[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13770_ (.CLK(clknet_leaf_52_clk),
    .D(_00224_),
    .Q(\cpuregs[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13771_ (.CLK(clknet_leaf_70_clk),
    .D(_00225_),
    .Q(\cpuregs[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13772_ (.CLK(clknet_leaf_52_clk),
    .D(_00226_),
    .Q(\cpuregs[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13773_ (.CLK(clknet_leaf_57_clk),
    .D(_00227_),
    .Q(\cpuregs[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13774_ (.CLK(clknet_leaf_37_clk),
    .D(_00228_),
    .Q(\cpuregs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13775_ (.CLK(clknet_leaf_47_clk),
    .D(_00229_),
    .Q(\cpuregs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13776_ (.CLK(clknet_leaf_32_clk),
    .D(_00230_),
    .Q(\cpuregs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13777_ (.CLK(clknet_leaf_22_clk),
    .D(_00231_),
    .Q(\cpuregs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13778_ (.CLK(clknet_leaf_23_clk),
    .D(_00232_),
    .Q(\cpuregs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13779_ (.CLK(clknet_leaf_22_clk),
    .D(_00233_),
    .Q(\cpuregs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13780_ (.CLK(clknet_leaf_179_clk),
    .D(_00234_),
    .Q(\cpuregs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13781_ (.CLK(clknet_leaf_20_clk),
    .D(_00235_),
    .Q(\cpuregs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13782_ (.CLK(clknet_leaf_180_clk),
    .D(_00236_),
    .Q(\cpuregs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13783_ (.CLK(clknet_leaf_181_clk),
    .D(_00237_),
    .Q(\cpuregs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13784_ (.CLK(clknet_leaf_181_clk),
    .D(_00238_),
    .Q(\cpuregs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13785_ (.CLK(clknet_leaf_5_clk),
    .D(_00239_),
    .Q(\cpuregs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13786_ (.CLK(clknet_leaf_6_clk),
    .D(_00240_),
    .Q(\cpuregs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13787_ (.CLK(clknet_leaf_5_clk),
    .D(_00241_),
    .Q(\cpuregs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13788_ (.CLK(clknet_leaf_19_clk),
    .D(_00242_),
    .Q(\cpuregs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13789_ (.CLK(clknet_leaf_7_clk),
    .D(_00243_),
    .Q(\cpuregs[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13790_ (.CLK(clknet_leaf_11_clk),
    .D(_00244_),
    .Q(\cpuregs[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13791_ (.CLK(clknet_leaf_7_clk),
    .D(_00245_),
    .Q(\cpuregs[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13792_ (.CLK(clknet_leaf_8_clk),
    .D(_00246_),
    .Q(\cpuregs[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13793_ (.CLK(clknet_leaf_41_clk),
    .D(_00247_),
    .Q(\cpuregs[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13794_ (.CLK(clknet_leaf_14_clk),
    .D(_00248_),
    .Q(\cpuregs[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13795_ (.CLK(clknet_leaf_16_clk),
    .D(_00249_),
    .Q(\cpuregs[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13796_ (.CLK(clknet_leaf_44_clk),
    .D(_00250_),
    .Q(\cpuregs[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13797_ (.CLK(clknet_leaf_17_clk),
    .D(_00251_),
    .Q(\cpuregs[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13798_ (.CLK(clknet_leaf_33_clk),
    .D(_00252_),
    .Q(\cpuregs[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13799_ (.CLK(clknet_leaf_71_clk),
    .D(_00253_),
    .Q(\cpuregs[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_34_clk),
    .D(_00254_),
    .Q(\cpuregs[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13801_ (.CLK(clknet_leaf_48_clk),
    .D(_00255_),
    .Q(\cpuregs[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_47_clk),
    .D(_00256_),
    .Q(\cpuregs[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13803_ (.CLK(clknet_leaf_72_clk),
    .D(_00257_),
    .Q(\cpuregs[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13804_ (.CLK(clknet_leaf_52_clk),
    .D(_00258_),
    .Q(\cpuregs[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13805_ (.CLK(clknet_leaf_49_clk),
    .D(_00259_),
    .Q(\cpuregs[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_36_clk),
    .D(_00260_),
    .Q(\cpuregs[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_45_clk),
    .D(_00261_),
    .Q(\cpuregs[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13808_ (.CLK(clknet_leaf_29_clk),
    .D(_00262_),
    .Q(\cpuregs[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13809_ (.CLK(clknet_leaf_21_clk),
    .D(_00263_),
    .Q(\cpuregs[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13810_ (.CLK(clknet_leaf_28_clk),
    .D(_00264_),
    .Q(\cpuregs[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13811_ (.CLK(clknet_leaf_24_clk),
    .D(_00265_),
    .Q(\cpuregs[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13812_ (.CLK(clknet_leaf_178_clk),
    .D(_00266_),
    .Q(\cpuregs[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13813_ (.CLK(clknet_leaf_190_clk),
    .D(_00267_),
    .Q(\cpuregs[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13814_ (.CLK(clknet_leaf_188_clk),
    .D(_00268_),
    .Q(\cpuregs[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13815_ (.CLK(clknet_leaf_182_clk),
    .D(_00269_),
    .Q(\cpuregs[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13816_ (.CLK(clknet_leaf_187_clk),
    .D(_00270_),
    .Q(\cpuregs[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13817_ (.CLK(clknet_leaf_191_clk),
    .D(_00271_),
    .Q(\cpuregs[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13818_ (.CLK(clknet_leaf_198_clk),
    .D(_00272_),
    .Q(\cpuregs[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13819_ (.CLK(clknet_leaf_196_clk),
    .D(_00273_),
    .Q(\cpuregs[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13820_ (.CLK(clknet_leaf_197_clk),
    .D(_00274_),
    .Q(\cpuregs[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13821_ (.CLK(clknet_leaf_198_clk),
    .D(_00275_),
    .Q(\cpuregs[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13822_ (.CLK(clknet_leaf_10_clk),
    .D(_00276_),
    .Q(\cpuregs[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13823_ (.CLK(clknet_leaf_0_clk),
    .D(_00277_),
    .Q(\cpuregs[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13824_ (.CLK(clknet_leaf_1_clk),
    .D(_00278_),
    .Q(\cpuregs[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13825_ (.CLK(clknet_leaf_42_clk),
    .D(_00279_),
    .Q(\cpuregs[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13826_ (.CLK(clknet_leaf_12_clk),
    .D(_00280_),
    .Q(\cpuregs[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13827_ (.CLK(clknet_leaf_13_clk),
    .D(_00281_),
    .Q(\cpuregs[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13828_ (.CLK(clknet_leaf_43_clk),
    .D(_00282_),
    .Q(\cpuregs[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13829_ (.CLK(clknet_leaf_23_clk),
    .D(_00283_),
    .Q(\cpuregs[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13830_ (.CLK(clknet_leaf_36_clk),
    .D(_00284_),
    .Q(\cpuregs[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13831_ (.CLK(clknet_leaf_71_clk),
    .D(_00285_),
    .Q(\cpuregs[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13832_ (.CLK(clknet_leaf_57_clk),
    .D(_00286_),
    .Q(\cpuregs[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13833_ (.CLK(clknet_leaf_48_clk),
    .D(_00287_),
    .Q(\cpuregs[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13834_ (.CLK(clknet_leaf_46_clk),
    .D(_00288_),
    .Q(\cpuregs[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13835_ (.CLK(clknet_leaf_68_clk),
    .D(_00289_),
    .Q(\cpuregs[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13836_ (.CLK(clknet_leaf_53_clk),
    .D(_00290_),
    .Q(\cpuregs[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_49_clk),
    .D(_00291_),
    .Q(\cpuregs[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_36_clk),
    .D(_00292_),
    .Q(\cpuregs[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_45_clk),
    .D(_00293_),
    .Q(\cpuregs[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_28_clk),
    .D(_00294_),
    .Q(\cpuregs[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_21_clk),
    .D(_00295_),
    .Q(\cpuregs[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_28_clk),
    .D(_00296_),
    .Q(\cpuregs[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13843_ (.CLK(clknet_leaf_24_clk),
    .D(_00297_),
    .Q(\cpuregs[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_178_clk),
    .D(_00298_),
    .Q(\cpuregs[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_190_clk),
    .D(_00299_),
    .Q(\cpuregs[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_187_clk),
    .D(_00300_),
    .Q(\cpuregs[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_182_clk),
    .D(_00301_),
    .Q(\cpuregs[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_188_clk),
    .D(_00302_),
    .Q(\cpuregs[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_191_clk),
    .D(_00303_),
    .Q(\cpuregs[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_198_clk),
    .D(_00304_),
    .Q(\cpuregs[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_196_clk),
    .D(_00305_),
    .Q(\cpuregs[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_197_clk),
    .D(_00306_),
    .Q(\cpuregs[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_199_clk),
    .D(_00307_),
    .Q(\cpuregs[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_10_clk),
    .D(_00308_),
    .Q(\cpuregs[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_0_clk),
    .D(_00309_),
    .Q(\cpuregs[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_1_clk),
    .D(_00310_),
    .Q(\cpuregs[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_42_clk),
    .D(_00311_),
    .Q(\cpuregs[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_12_clk),
    .D(_00312_),
    .Q(\cpuregs[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_12_clk),
    .D(_00313_),
    .Q(\cpuregs[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_43_clk),
    .D(_00314_),
    .Q(\cpuregs[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_23_clk),
    .D(_00315_),
    .Q(\cpuregs[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_36_clk),
    .D(_00316_),
    .Q(\cpuregs[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_72_clk),
    .D(_00317_),
    .Q(\cpuregs[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_57_clk),
    .D(_00318_),
    .Q(\cpuregs[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_48_clk),
    .D(_00319_),
    .Q(\cpuregs[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13866_ (.CLK(clknet_leaf_46_clk),
    .D(_00320_),
    .Q(\cpuregs[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_68_clk),
    .D(_00321_),
    .Q(\cpuregs[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_53_clk),
    .D(_00322_),
    .Q(\cpuregs[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_49_clk),
    .D(_00323_),
    .Q(\cpuregs[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13870_ (.CLK(clknet_leaf_38_clk),
    .D(_00324_),
    .Q(\cpuregs[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_47_clk),
    .D(_00325_),
    .Q(\cpuregs[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_73_clk),
    .D(_00326_),
    .Q(\cpuregs[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_176_clk),
    .D(_00327_),
    .Q(\cpuregs[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13874_ (.CLK(clknet_leaf_25_clk),
    .D(_00328_),
    .Q(\cpuregs[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13875_ (.CLK(clknet_leaf_25_clk),
    .D(_00329_),
    .Q(\cpuregs[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_178_clk),
    .D(_00330_),
    .Q(\cpuregs[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_188_clk),
    .D(_00331_),
    .Q(\cpuregs[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13878_ (.CLK(clknet_leaf_185_clk),
    .D(_00332_),
    .Q(\cpuregs[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_185_clk),
    .D(_00333_),
    .Q(\cpuregs[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_186_clk),
    .D(_00334_),
    .Q(\cpuregs[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_191_clk),
    .D(_00335_),
    .Q(\cpuregs[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_196_clk),
    .D(_00336_),
    .Q(\cpuregs[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_196_clk),
    .D(_00337_),
    .Q(\cpuregs[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_191_clk),
    .D(_00338_),
    .Q(\cpuregs[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13885_ (.CLK(clknet_leaf_199_clk),
    .D(_00339_),
    .Q(\cpuregs[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_7_clk),
    .D(_00340_),
    .Q(\cpuregs[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_2_clk),
    .D(_00341_),
    .Q(\cpuregs[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13888_ (.CLK(clknet_leaf_2_clk),
    .D(_00342_),
    .Q(\cpuregs[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_41_clk),
    .D(_00343_),
    .Q(\cpuregs[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_15_clk),
    .D(_00344_),
    .Q(\cpuregs[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_14_clk),
    .D(_00345_),
    .Q(\cpuregs[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_40_clk),
    .D(_00346_),
    .Q(\cpuregs[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_30_clk),
    .D(_00347_),
    .Q(\cpuregs[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_30_clk),
    .D(_00348_),
    .Q(\cpuregs[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_60_clk),
    .D(_00349_),
    .Q(\cpuregs[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_59_clk),
    .D(_00350_),
    .Q(\cpuregs[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_56_clk),
    .D(_00351_),
    .Q(\cpuregs[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_51_clk),
    .D(_00352_),
    .Q(\cpuregs[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_66_clk),
    .D(_00353_),
    .Q(\cpuregs[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_54_clk),
    .D(_00354_),
    .Q(\cpuregs[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13901_ (.CLK(clknet_leaf_56_clk),
    .D(_00355_),
    .Q(\cpuregs[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_37_clk),
    .D(_00356_),
    .Q(\cpuregs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13903_ (.CLK(clknet_leaf_47_clk),
    .D(_00357_),
    .Q(\cpuregs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13904_ (.CLK(clknet_leaf_32_clk),
    .D(_00358_),
    .Q(\cpuregs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13905_ (.CLK(clknet_leaf_22_clk),
    .D(_00359_),
    .Q(\cpuregs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_23_clk),
    .D(_00360_),
    .Q(\cpuregs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_23_clk),
    .D(_00361_),
    .Q(\cpuregs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_179_clk),
    .D(_00362_),
    .Q(\cpuregs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_20_clk),
    .D(_00363_),
    .Q(\cpuregs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_180_clk),
    .D(_00364_),
    .Q(\cpuregs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_181_clk),
    .D(_00365_),
    .Q(\cpuregs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13912_ (.CLK(clknet_leaf_181_clk),
    .D(_00366_),
    .Q(\cpuregs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_5_clk),
    .D(_00367_),
    .Q(\cpuregs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_6_clk),
    .D(_00368_),
    .Q(\cpuregs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_5_clk),
    .D(_00369_),
    .Q(\cpuregs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_19_clk),
    .D(_00370_),
    .Q(\cpuregs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_7_clk),
    .D(_00371_),
    .Q(\cpuregs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_18_clk),
    .D(_00372_),
    .Q(\cpuregs[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13919_ (.CLK(clknet_leaf_6_clk),
    .D(_00373_),
    .Q(\cpuregs[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_8_clk),
    .D(_00374_),
    .Q(\cpuregs[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_14_clk),
    .D(_00375_),
    .Q(\cpuregs[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_15_clk),
    .D(_00376_),
    .Q(\cpuregs[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13923_ (.CLK(clknet_leaf_16_clk),
    .D(_00377_),
    .Q(\cpuregs[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13924_ (.CLK(clknet_leaf_44_clk),
    .D(_00378_),
    .Q(\cpuregs[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13925_ (.CLK(clknet_leaf_23_clk),
    .D(_00379_),
    .Q(\cpuregs[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13926_ (.CLK(clknet_leaf_33_clk),
    .D(_00380_),
    .Q(\cpuregs[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13927_ (.CLK(clknet_leaf_32_clk),
    .D(_00381_),
    .Q(\cpuregs[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13928_ (.CLK(clknet_leaf_33_clk),
    .D(_00382_),
    .Q(\cpuregs[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13929_ (.CLK(clknet_leaf_48_clk),
    .D(_00383_),
    .Q(\cpuregs[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_46_clk),
    .D(_00384_),
    .Q(\cpuregs[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_72_clk),
    .D(_00385_),
    .Q(\cpuregs[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13932_ (.CLK(clknet_leaf_46_clk),
    .D(_00386_),
    .Q(\cpuregs[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_49_clk),
    .D(_00387_),
    .Q(\cpuregs[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13934_ (.CLK(clknet_leaf_39_clk),
    .D(_00388_),
    .Q(\cpuregs[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13935_ (.CLK(clknet_leaf_44_clk),
    .D(_00389_),
    .Q(\cpuregs[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_76_clk),
    .D(_00390_),
    .Q(\cpuregs[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_176_clk),
    .D(_00391_),
    .Q(\cpuregs[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_26_clk),
    .D(_00392_),
    .Q(\cpuregs[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_176_clk),
    .D(_00393_),
    .Q(\cpuregs[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_178_clk),
    .D(_00394_),
    .Q(\cpuregs[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_188_clk),
    .D(_00395_),
    .Q(\cpuregs[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_185_clk),
    .D(_00396_),
    .Q(\cpuregs[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_185_clk),
    .D(_00397_),
    .Q(\cpuregs[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_186_clk),
    .D(_00398_),
    .Q(\cpuregs[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_190_clk),
    .D(_00399_),
    .Q(\cpuregs[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_198_clk),
    .D(_00400_),
    .Q(\cpuregs[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_197_clk),
    .D(_00401_),
    .Q(\cpuregs[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13948_ (.CLK(clknet_leaf_191_clk),
    .D(_00402_),
    .Q(\cpuregs[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13949_ (.CLK(clknet_leaf_198_clk),
    .D(_00403_),
    .Q(\cpuregs[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13950_ (.CLK(clknet_leaf_11_clk),
    .D(_00404_),
    .Q(\cpuregs[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13951_ (.CLK(clknet_leaf_2_clk),
    .D(_00405_),
    .Q(\cpuregs[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13952_ (.CLK(clknet_leaf_2_clk),
    .D(_00406_),
    .Q(\cpuregs[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13953_ (.CLK(clknet_leaf_41_clk),
    .D(_00407_),
    .Q(\cpuregs[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13954_ (.CLK(clknet_leaf_15_clk),
    .D(_00408_),
    .Q(\cpuregs[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13955_ (.CLK(clknet_leaf_14_clk),
    .D(_00409_),
    .Q(\cpuregs[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13956_ (.CLK(clknet_leaf_40_clk),
    .D(_00410_),
    .Q(\cpuregs[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13957_ (.CLK(clknet_leaf_30_clk),
    .D(_00411_),
    .Q(\cpuregs[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13958_ (.CLK(clknet_leaf_30_clk),
    .D(_00412_),
    .Q(\cpuregs[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13959_ (.CLK(clknet_leaf_60_clk),
    .D(_00413_),
    .Q(\cpuregs[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13960_ (.CLK(clknet_leaf_59_clk),
    .D(_00414_),
    .Q(\cpuregs[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13961_ (.CLK(clknet_leaf_56_clk),
    .D(_00415_),
    .Q(\cpuregs[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13962_ (.CLK(clknet_leaf_52_clk),
    .D(_00416_),
    .Q(\cpuregs[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13963_ (.CLK(clknet_leaf_66_clk),
    .D(_00417_),
    .Q(\cpuregs[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13964_ (.CLK(clknet_leaf_51_clk),
    .D(_00418_),
    .Q(\cpuregs[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13965_ (.CLK(clknet_leaf_56_clk),
    .D(_00419_),
    .Q(\cpuregs[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13966_ (.CLK(clknet_leaf_36_clk),
    .D(_00420_),
    .Q(\cpuregs[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13967_ (.CLK(clknet_leaf_45_clk),
    .D(_00421_),
    .Q(\cpuregs[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13968_ (.CLK(clknet_leaf_28_clk),
    .D(_00422_),
    .Q(\cpuregs[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13969_ (.CLK(clknet_leaf_21_clk),
    .D(_00423_),
    .Q(\cpuregs[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13970_ (.CLK(clknet_leaf_29_clk),
    .D(_00424_),
    .Q(\cpuregs[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13971_ (.CLK(clknet_leaf_25_clk),
    .D(_00425_),
    .Q(\cpuregs[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13972_ (.CLK(clknet_leaf_178_clk),
    .D(_00426_),
    .Q(\cpuregs[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13973_ (.CLK(clknet_leaf_190_clk),
    .D(_00427_),
    .Q(\cpuregs[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13974_ (.CLK(clknet_leaf_190_clk),
    .D(_00428_),
    .Q(\cpuregs[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13975_ (.CLK(clknet_leaf_183_clk),
    .D(_00429_),
    .Q(\cpuregs[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13976_ (.CLK(clknet_leaf_190_clk),
    .D(_00430_),
    .Q(\cpuregs[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13977_ (.CLK(clknet_leaf_191_clk),
    .D(_00431_),
    .Q(\cpuregs[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13978_ (.CLK(clknet_leaf_198_clk),
    .D(_00432_),
    .Q(\cpuregs[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13979_ (.CLK(clknet_leaf_196_clk),
    .D(_00433_),
    .Q(\cpuregs[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13980_ (.CLK(clknet_leaf_197_clk),
    .D(_00434_),
    .Q(\cpuregs[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13981_ (.CLK(clknet_leaf_199_clk),
    .D(_00435_),
    .Q(\cpuregs[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13982_ (.CLK(clknet_leaf_10_clk),
    .D(_00436_),
    .Q(\cpuregs[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _13983_ (.CLK(clknet_leaf_0_clk),
    .D(_00437_),
    .Q(\cpuregs[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_0_clk),
    .D(_00438_),
    .Q(\cpuregs[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_42_clk),
    .D(_00439_),
    .Q(\cpuregs[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_12_clk),
    .D(_00440_),
    .Q(\cpuregs[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _13987_ (.CLK(clknet_leaf_13_clk),
    .D(_00441_),
    .Q(\cpuregs[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _13988_ (.CLK(clknet_leaf_43_clk),
    .D(_00442_),
    .Q(\cpuregs[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _13989_ (.CLK(clknet_leaf_22_clk),
    .D(_00443_),
    .Q(\cpuregs[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _13990_ (.CLK(clknet_leaf_35_clk),
    .D(_00444_),
    .Q(\cpuregs[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _13991_ (.CLK(clknet_leaf_71_clk),
    .D(_00445_),
    .Q(\cpuregs[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _13992_ (.CLK(clknet_leaf_71_clk),
    .D(_00446_),
    .Q(\cpuregs[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _13993_ (.CLK(clknet_leaf_49_clk),
    .D(_00447_),
    .Q(\cpuregs[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _13994_ (.CLK(clknet_leaf_45_clk),
    .D(_00448_),
    .Q(\cpuregs[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _13995_ (.CLK(clknet_leaf_68_clk),
    .D(_00449_),
    .Q(\cpuregs[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _13996_ (.CLK(clknet_leaf_53_clk),
    .D(_00450_),
    .Q(\cpuregs[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _13997_ (.CLK(clknet_leaf_50_clk),
    .D(_00451_),
    .Q(\cpuregs[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _13998_ (.CLK(clknet_leaf_36_clk),
    .D(_00452_),
    .Q(\cpuregs[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13999_ (.CLK(clknet_leaf_45_clk),
    .D(_00453_),
    .Q(\cpuregs[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14000_ (.CLK(clknet_leaf_29_clk),
    .D(_00454_),
    .Q(\cpuregs[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14001_ (.CLK(clknet_leaf_21_clk),
    .D(_00455_),
    .Q(\cpuregs[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14002_ (.CLK(clknet_leaf_29_clk),
    .D(_00456_),
    .Q(\cpuregs[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14003_ (.CLK(clknet_leaf_25_clk),
    .D(_00457_),
    .Q(\cpuregs[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14004_ (.CLK(clknet_leaf_178_clk),
    .D(_00458_),
    .Q(\cpuregs[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14005_ (.CLK(clknet_leaf_190_clk),
    .D(_00459_),
    .Q(\cpuregs[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14006_ (.CLK(clknet_leaf_190_clk),
    .D(_00460_),
    .Q(\cpuregs[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14007_ (.CLK(clknet_leaf_183_clk),
    .D(_00461_),
    .Q(\cpuregs[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14008_ (.CLK(clknet_leaf_190_clk),
    .D(_00462_),
    .Q(\cpuregs[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14009_ (.CLK(clknet_leaf_191_clk),
    .D(_00463_),
    .Q(\cpuregs[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14010_ (.CLK(clknet_leaf_198_clk),
    .D(_00464_),
    .Q(\cpuregs[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14011_ (.CLK(clknet_leaf_196_clk),
    .D(_00465_),
    .Q(\cpuregs[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14012_ (.CLK(clknet_leaf_197_clk),
    .D(_00466_),
    .Q(\cpuregs[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14013_ (.CLK(clknet_leaf_199_clk),
    .D(_00467_),
    .Q(\cpuregs[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14014_ (.CLK(clknet_leaf_10_clk),
    .D(_00468_),
    .Q(\cpuregs[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14015_ (.CLK(clknet_leaf_0_clk),
    .D(_00469_),
    .Q(\cpuregs[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14016_ (.CLK(clknet_leaf_1_clk),
    .D(_00470_),
    .Q(\cpuregs[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14017_ (.CLK(clknet_leaf_42_clk),
    .D(_00471_),
    .Q(\cpuregs[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14018_ (.CLK(clknet_leaf_12_clk),
    .D(_00472_),
    .Q(\cpuregs[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14019_ (.CLK(clknet_leaf_13_clk),
    .D(_00473_),
    .Q(\cpuregs[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14020_ (.CLK(clknet_leaf_43_clk),
    .D(_00474_),
    .Q(\cpuregs[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14021_ (.CLK(clknet_leaf_23_clk),
    .D(_00475_),
    .Q(\cpuregs[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14022_ (.CLK(clknet_leaf_36_clk),
    .D(_00476_),
    .Q(\cpuregs[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14023_ (.CLK(clknet_leaf_71_clk),
    .D(_00477_),
    .Q(\cpuregs[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14024_ (.CLK(clknet_leaf_71_clk),
    .D(_00478_),
    .Q(\cpuregs[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14025_ (.CLK(clknet_leaf_49_clk),
    .D(_00479_),
    .Q(\cpuregs[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14026_ (.CLK(clknet_leaf_45_clk),
    .D(_00480_),
    .Q(\cpuregs[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14027_ (.CLK(clknet_leaf_68_clk),
    .D(_00481_),
    .Q(\cpuregs[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14028_ (.CLK(clknet_leaf_53_clk),
    .D(_00482_),
    .Q(\cpuregs[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14029_ (.CLK(clknet_leaf_50_clk),
    .D(_00483_),
    .Q(\cpuregs[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14030_ (.CLK(clknet_leaf_39_clk),
    .D(_00484_),
    .Q(\cpuregs[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14031_ (.CLK(clknet_leaf_45_clk),
    .D(_00485_),
    .Q(\cpuregs[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14032_ (.CLK(clknet_leaf_32_clk),
    .D(_00486_),
    .Q(\cpuregs[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14033_ (.CLK(clknet_leaf_179_clk),
    .D(_00487_),
    .Q(\cpuregs[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14034_ (.CLK(clknet_leaf_23_clk),
    .D(_00488_),
    .Q(\cpuregs[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14035_ (.CLK(clknet_leaf_25_clk),
    .D(_00489_),
    .Q(\cpuregs[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14036_ (.CLK(clknet_leaf_179_clk),
    .D(_00490_),
    .Q(\cpuregs[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14037_ (.CLK(clknet_leaf_187_clk),
    .D(_00491_),
    .Q(\cpuregs[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14038_ (.CLK(clknet_leaf_185_clk),
    .D(_00492_),
    .Q(\cpuregs[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14039_ (.CLK(clknet_leaf_184_clk),
    .D(_00493_),
    .Q(\cpuregs[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14040_ (.CLK(clknet_leaf_186_clk),
    .D(_00494_),
    .Q(\cpuregs[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14041_ (.CLK(clknet_leaf_191_clk),
    .D(_00495_),
    .Q(\cpuregs[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14042_ (.CLK(clknet_leaf_196_clk),
    .D(_00496_),
    .Q(\cpuregs[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14043_ (.CLK(clknet_leaf_195_clk),
    .D(_00497_),
    .Q(\cpuregs[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14044_ (.CLK(clknet_leaf_195_clk),
    .D(_00498_),
    .Q(\cpuregs[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14045_ (.CLK(clknet_leaf_199_clk),
    .D(_00499_),
    .Q(\cpuregs[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14046_ (.CLK(clknet_leaf_10_clk),
    .D(_00500_),
    .Q(\cpuregs[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14047_ (.CLK(clknet_leaf_0_clk),
    .D(_00501_),
    .Q(\cpuregs[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14048_ (.CLK(clknet_leaf_1_clk),
    .D(_00502_),
    .Q(\cpuregs[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14049_ (.CLK(clknet_leaf_41_clk),
    .D(_00503_),
    .Q(\cpuregs[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14050_ (.CLK(clknet_leaf_11_clk),
    .D(_00504_),
    .Q(\cpuregs[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14051_ (.CLK(clknet_leaf_13_clk),
    .D(_00505_),
    .Q(\cpuregs[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14052_ (.CLK(clknet_leaf_44_clk),
    .D(_00506_),
    .Q(\cpuregs[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14053_ (.CLK(clknet_leaf_38_clk),
    .D(_00507_),
    .Q(\cpuregs[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14054_ (.CLK(clknet_leaf_37_clk),
    .D(_00508_),
    .Q(\cpuregs[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14055_ (.CLK(clknet_leaf_60_clk),
    .D(_00509_),
    .Q(\cpuregs[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14056_ (.CLK(clknet_leaf_58_clk),
    .D(_00510_),
    .Q(\cpuregs[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14057_ (.CLK(clknet_leaf_50_clk),
    .D(_00511_),
    .Q(\cpuregs[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14058_ (.CLK(clknet_leaf_52_clk),
    .D(_00512_),
    .Q(\cpuregs[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14059_ (.CLK(clknet_leaf_66_clk),
    .D(_00513_),
    .Q(\cpuregs[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14060_ (.CLK(clknet_leaf_54_clk),
    .D(_00514_),
    .Q(\cpuregs[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14061_ (.CLK(clknet_leaf_50_clk),
    .D(_00515_),
    .Q(\cpuregs[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14062_ (.CLK(clknet_leaf_39_clk),
    .D(_00516_),
    .Q(\cpuregs[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14063_ (.CLK(clknet_leaf_44_clk),
    .D(_00517_),
    .Q(\cpuregs[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14064_ (.CLK(clknet_leaf_76_clk),
    .D(_00518_),
    .Q(\cpuregs[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14065_ (.CLK(clknet_leaf_179_clk),
    .D(_00519_),
    .Q(\cpuregs[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14066_ (.CLK(clknet_leaf_26_clk),
    .D(_00520_),
    .Q(\cpuregs[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14067_ (.CLK(clknet_leaf_176_clk),
    .D(_00521_),
    .Q(\cpuregs[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14068_ (.CLK(clknet_leaf_185_clk),
    .D(_00522_),
    .Q(\cpuregs[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14069_ (.CLK(clknet_leaf_188_clk),
    .D(_00523_),
    .Q(\cpuregs[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14070_ (.CLK(clknet_leaf_185_clk),
    .D(_00524_),
    .Q(\cpuregs[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14071_ (.CLK(clknet_leaf_185_clk),
    .D(_00525_),
    .Q(\cpuregs[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14072_ (.CLK(clknet_leaf_186_clk),
    .D(_00526_),
    .Q(\cpuregs[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14073_ (.CLK(clknet_leaf_190_clk),
    .D(_00527_),
    .Q(\cpuregs[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14074_ (.CLK(clknet_leaf_198_clk),
    .D(_00528_),
    .Q(\cpuregs[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14075_ (.CLK(clknet_leaf_197_clk),
    .D(_00529_),
    .Q(\cpuregs[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14076_ (.CLK(clknet_leaf_191_clk),
    .D(_00530_),
    .Q(\cpuregs[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14077_ (.CLK(clknet_leaf_198_clk),
    .D(_00531_),
    .Q(\cpuregs[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14078_ (.CLK(clknet_leaf_7_clk),
    .D(_00532_),
    .Q(\cpuregs[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14079_ (.CLK(clknet_leaf_2_clk),
    .D(_00533_),
    .Q(\cpuregs[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14080_ (.CLK(clknet_leaf_2_clk),
    .D(_00534_),
    .Q(\cpuregs[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14081_ (.CLK(clknet_leaf_41_clk),
    .D(_00535_),
    .Q(\cpuregs[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14082_ (.CLK(clknet_leaf_18_clk),
    .D(_00536_),
    .Q(\cpuregs[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14083_ (.CLK(clknet_leaf_14_clk),
    .D(_00537_),
    .Q(\cpuregs[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14084_ (.CLK(clknet_leaf_40_clk),
    .D(_00538_),
    .Q(\cpuregs[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14085_ (.CLK(clknet_leaf_30_clk),
    .D(_00539_),
    .Q(\cpuregs[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14086_ (.CLK(clknet_leaf_30_clk),
    .D(_00540_),
    .Q(\cpuregs[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14087_ (.CLK(clknet_leaf_60_clk),
    .D(_00541_),
    .Q(\cpuregs[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14088_ (.CLK(clknet_leaf_59_clk),
    .D(_00542_),
    .Q(\cpuregs[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14089_ (.CLK(clknet_leaf_56_clk),
    .D(_00543_),
    .Q(\cpuregs[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14090_ (.CLK(clknet_leaf_52_clk),
    .D(_00544_),
    .Q(\cpuregs[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14091_ (.CLK(clknet_leaf_66_clk),
    .D(_00545_),
    .Q(\cpuregs[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14092_ (.CLK(clknet_leaf_51_clk),
    .D(_00546_),
    .Q(\cpuregs[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14093_ (.CLK(clknet_leaf_56_clk),
    .D(_00547_),
    .Q(\cpuregs[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14094_ (.CLK(clknet_leaf_39_clk),
    .D(_00548_),
    .Q(\cpuregs[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14095_ (.CLK(clknet_leaf_47_clk),
    .D(_00549_),
    .Q(\cpuregs[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14096_ (.CLK(clknet_leaf_32_clk),
    .D(_00550_),
    .Q(\cpuregs[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14097_ (.CLK(clknet_leaf_179_clk),
    .D(_00551_),
    .Q(\cpuregs[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14098_ (.CLK(clknet_leaf_24_clk),
    .D(_00552_),
    .Q(\cpuregs[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14099_ (.CLK(clknet_leaf_25_clk),
    .D(_00553_),
    .Q(\cpuregs[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14100_ (.CLK(clknet_leaf_178_clk),
    .D(_00554_),
    .Q(\cpuregs[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14101_ (.CLK(clknet_leaf_186_clk),
    .D(_00555_),
    .Q(\cpuregs[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14102_ (.CLK(clknet_leaf_185_clk),
    .D(_00556_),
    .Q(\cpuregs[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14103_ (.CLK(clknet_leaf_185_clk),
    .D(_00557_),
    .Q(\cpuregs[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14104_ (.CLK(clknet_leaf_186_clk),
    .D(_00558_),
    .Q(\cpuregs[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14105_ (.CLK(clknet_leaf_192_clk),
    .D(_00559_),
    .Q(\cpuregs[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14106_ (.CLK(clknet_leaf_196_clk),
    .D(_00560_),
    .Q(\cpuregs[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14107_ (.CLK(clknet_leaf_195_clk),
    .D(_00561_),
    .Q(\cpuregs[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14108_ (.CLK(clknet_leaf_195_clk),
    .D(_00562_),
    .Q(\cpuregs[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14109_ (.CLK(clknet_leaf_199_clk),
    .D(_00563_),
    .Q(\cpuregs[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14110_ (.CLK(clknet_leaf_11_clk),
    .D(_00564_),
    .Q(\cpuregs[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14111_ (.CLK(clknet_leaf_2_clk),
    .D(_00565_),
    .Q(\cpuregs[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14112_ (.CLK(clknet_leaf_2_clk),
    .D(_00566_),
    .Q(\cpuregs[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14113_ (.CLK(clknet_leaf_41_clk),
    .D(_00567_),
    .Q(\cpuregs[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14114_ (.CLK(clknet_leaf_11_clk),
    .D(_00568_),
    .Q(\cpuregs[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14115_ (.CLK(clknet_leaf_13_clk),
    .D(_00569_),
    .Q(\cpuregs[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14116_ (.CLK(clknet_leaf_44_clk),
    .D(_00570_),
    .Q(\cpuregs[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14117_ (.CLK(clknet_leaf_37_clk),
    .D(_00571_),
    .Q(\cpuregs[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14118_ (.CLK(clknet_leaf_30_clk),
    .D(_00572_),
    .Q(\cpuregs[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14119_ (.CLK(clknet_leaf_69_clk),
    .D(_00573_),
    .Q(\cpuregs[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14120_ (.CLK(clknet_leaf_58_clk),
    .D(_00574_),
    .Q(\cpuregs[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14121_ (.CLK(clknet_leaf_56_clk),
    .D(_00575_),
    .Q(\cpuregs[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14122_ (.CLK(clknet_leaf_52_clk),
    .D(_00576_),
    .Q(\cpuregs[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14123_ (.CLK(clknet_leaf_66_clk),
    .D(_00577_),
    .Q(\cpuregs[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14124_ (.CLK(clknet_leaf_54_clk),
    .D(_00578_),
    .Q(\cpuregs[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_50_clk),
    .D(_00579_),
    .Q(\cpuregs[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_98_clk),
    .D(_00580_),
    .Q(\genblk2.pcpi_div.instr_remu ));
 sky130_fd_sc_hd__dfxtp_2 _14127_ (.CLK(clknet_leaf_92_clk),
    .D(_00581_),
    .Q(net267));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_91_clk),
    .D(_00582_),
    .Q(net268));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_83_clk),
    .D(_00583_),
    .Q(\count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_83_clk),
    .D(_00584_),
    .Q(\count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_127_clk),
    .D(_00585_),
    .Q(\count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_127_clk),
    .D(_00586_),
    .Q(\count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_127_clk),
    .D(_00587_),
    .Q(\count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_127_clk),
    .D(_00588_),
    .Q(\count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_125_clk),
    .D(_00589_),
    .Q(\count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_125_clk),
    .D(_00590_),
    .Q(\count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_125_clk),
    .D(_00591_),
    .Q(\count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_126_clk),
    .D(_00592_),
    .Q(\count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_126_clk),
    .D(_00593_),
    .Q(\count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_126_clk),
    .D(_00594_),
    .Q(\count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_126_clk),
    .D(_00595_),
    .Q(\count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14142_ (.CLK(clknet_leaf_110_clk),
    .D(_00596_),
    .Q(\count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14143_ (.CLK(clknet_leaf_110_clk),
    .D(_00597_),
    .Q(\count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14144_ (.CLK(clknet_leaf_110_clk),
    .D(_00598_),
    .Q(\count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14145_ (.CLK(clknet_leaf_110_clk),
    .D(_00599_),
    .Q(\count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14146_ (.CLK(clknet_leaf_110_clk),
    .D(net2562),
    .Q(\count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_97_clk),
    .D(_00601_),
    .Q(\count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_97_clk),
    .D(_00602_),
    .Q(\count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14149_ (.CLK(clknet_leaf_97_clk),
    .D(_00603_),
    .Q(\count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14150_ (.CLK(clknet_leaf_97_clk),
    .D(_00604_),
    .Q(\count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_99_clk),
    .D(_00605_),
    .Q(\count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_100_clk),
    .D(net2616),
    .Q(\count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_100_clk),
    .D(_00607_),
    .Q(\count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_100_clk),
    .D(_00608_),
    .Q(\count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_100_clk),
    .D(_00609_),
    .Q(\count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_100_clk),
    .D(_00610_),
    .Q(\count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_100_clk),
    .D(_00611_),
    .Q(\count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_94_clk),
    .D(_00612_),
    .Q(\count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_94_clk),
    .D(_00613_),
    .Q(\count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_94_clk),
    .D(_00614_),
    .Q(\count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_126_clk),
    .D(_00615_),
    .Q(\count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_126_clk),
    .D(_00616_),
    .Q(\count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_126_clk),
    .D(net2583),
    .Q(\count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_126_clk),
    .D(_00618_),
    .Q(\count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_126_clk),
    .D(_00619_),
    .Q(\count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_126_clk),
    .D(_00620_),
    .Q(\count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_126_clk),
    .D(_00621_),
    .Q(\count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_126_clk),
    .D(_00622_),
    .Q(\count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_125_clk),
    .D(_00623_),
    .Q(\count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_125_clk),
    .D(_00624_),
    .Q(\count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_111_clk),
    .D(_00625_),
    .Q(\count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_111_clk),
    .D(_00626_),
    .Q(\count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_111_clk),
    .D(_00627_),
    .Q(\count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_111_clk),
    .D(_00628_),
    .Q(\count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_111_clk),
    .D(_00629_),
    .Q(\count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_111_clk),
    .D(_00630_),
    .Q(\count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_109_clk),
    .D(_00631_),
    .Q(\count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_109_clk),
    .D(net2585),
    .Q(\count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_109_clk),
    .D(_00633_),
    .Q(\count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_109_clk),
    .D(_00634_),
    .Q(\count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_109_clk),
    .D(_00635_),
    .Q(\count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_109_clk),
    .D(net2591),
    .Q(\count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_102_clk),
    .D(_00637_),
    .Q(\count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_102_clk),
    .D(_00638_),
    .Q(\count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_100_clk),
    .D(_00639_),
    .Q(\count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_100_clk),
    .D(_00640_),
    .Q(\count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_100_clk),
    .D(_00641_),
    .Q(\count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_100_clk),
    .D(_00642_),
    .Q(\count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_101_clk),
    .D(_00643_),
    .Q(\count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_94_clk),
    .D(_00644_),
    .Q(\count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_94_clk),
    .D(_00645_),
    .Q(\count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_94_clk),
    .D(_00646_),
    .Q(\count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_2 _14193_ (.CLK(clknet_leaf_132_clk),
    .D(_00647_),
    .Q(\reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14194_ (.CLK(clknet_leaf_132_clk),
    .D(_00648_),
    .Q(\reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14195_ (.CLK(clknet_leaf_132_clk),
    .D(_00649_),
    .Q(\reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_132_clk),
    .D(_00650_),
    .Q(\reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_133_clk),
    .D(_00651_),
    .Q(\reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_174_clk),
    .D(_00652_),
    .Q(\reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_174_clk),
    .D(_00653_),
    .Q(\reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_173_clk),
    .D(_00654_),
    .Q(\reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_173_clk),
    .D(_00655_),
    .Q(\reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14202_ (.CLK(clknet_leaf_177_clk),
    .D(_00656_),
    .Q(\reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_177_clk),
    .D(_00657_),
    .Q(\reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14204_ (.CLK(clknet_leaf_177_clk),
    .D(_00658_),
    .Q(\reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_177_clk),
    .D(_00659_),
    .Q(\reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14206_ (.CLK(clknet_leaf_176_clk),
    .D(_00660_),
    .Q(\reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_176_clk),
    .D(_00661_),
    .Q(\reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14208_ (.CLK(clknet_leaf_25_clk),
    .D(_00662_),
    .Q(\reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_26_clk),
    .D(_00663_),
    .Q(\reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14210_ (.CLK(clknet_leaf_27_clk),
    .D(_00664_),
    .Q(\reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _14211_ (.CLK(clknet_leaf_26_clk),
    .D(_00665_),
    .Q(\reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _14212_ (.CLK(clknet_leaf_77_clk),
    .D(_00666_),
    .Q(\reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_76_clk),
    .D(_00667_),
    .Q(\reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_76_clk),
    .D(_00668_),
    .Q(\reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _14215_ (.CLK(clknet_leaf_75_clk),
    .D(_00669_),
    .Q(\reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14216_ (.CLK(clknet_leaf_75_clk),
    .D(_00670_),
    .Q(\reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14217_ (.CLK(clknet_leaf_75_clk),
    .D(_00671_),
    .Q(\reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _14218_ (.CLK(clknet_leaf_68_clk),
    .D(_00672_),
    .Q(\reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14219_ (.CLK(clknet_leaf_67_clk),
    .D(_00673_),
    .Q(\reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14220_ (.CLK(clknet_leaf_67_clk),
    .D(_00674_),
    .Q(\reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14221_ (.CLK(clknet_leaf_66_clk),
    .D(_00675_),
    .Q(\reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14222_ (.CLK(clknet_leaf_67_clk),
    .D(_00676_),
    .Q(\reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14223_ (.CLK(clknet_leaf_87_clk),
    .D(_00677_),
    .Q(\reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14224_ (.CLK(clknet_leaf_78_clk),
    .D(_00678_),
    .Q(\reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14225_ (.CLK(clknet_leaf_132_clk),
    .D(_00679_),
    .Q(\reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14226_ (.CLK(clknet_leaf_132_clk),
    .D(_00680_),
    .Q(\reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_132_clk),
    .D(_00681_),
    .Q(\reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14228_ (.CLK(clknet_leaf_175_clk),
    .D(_00682_),
    .Q(\reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14229_ (.CLK(clknet_leaf_174_clk),
    .D(_00683_),
    .Q(\reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_174_clk),
    .D(_00684_),
    .Q(\reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_173_clk),
    .D(_00685_),
    .Q(\reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_173_clk),
    .D(_00686_),
    .Q(\reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_173_clk),
    .D(_00687_),
    .Q(\reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_177_clk),
    .D(_00688_),
    .Q(\reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_177_clk),
    .D(_00689_),
    .Q(\reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_177_clk),
    .D(_00690_),
    .Q(\reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_177_clk),
    .D(_00691_),
    .Q(\reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_176_clk),
    .D(_00692_),
    .Q(\reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_175_clk),
    .D(_00693_),
    .Q(\reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_26_clk),
    .D(_00694_),
    .Q(\reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_27_clk),
    .D(_00695_),
    .Q(\reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_27_clk),
    .D(_00696_),
    .Q(\reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_76_clk),
    .D(_00697_),
    .Q(\reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_76_clk),
    .D(_00698_),
    .Q(\reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_76_clk),
    .D(_00699_),
    .Q(\reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_75_clk),
    .D(_00700_),
    .Q(\reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_75_clk),
    .D(_00701_),
    .Q(\reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_75_clk),
    .D(_00702_),
    .Q(\reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_68_clk),
    .D(_00703_),
    .Q(\reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_68_clk),
    .D(_00704_),
    .Q(\reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_68_clk),
    .D(_00705_),
    .Q(\reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_66_clk),
    .D(_00706_),
    .Q(\reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_66_clk),
    .D(_00707_),
    .Q(\reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_87_clk),
    .D(_00708_),
    .Q(\reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_127_clk),
    .D(_00709_),
    .Q(\count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_127_clk),
    .D(net2907),
    .Q(\count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_127_clk),
    .D(_00711_),
    .Q(\count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_128_clk),
    .D(_00712_),
    .Q(\count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_128_clk),
    .D(_00713_),
    .Q(\count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_129_clk),
    .D(_00714_),
    .Q(\count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_123_clk),
    .D(_00715_),
    .Q(\count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_122_clk),
    .D(_00716_),
    .Q(\count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_122_clk),
    .D(_00717_),
    .Q(\count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_122_clk),
    .D(_00718_),
    .Q(\count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_122_clk),
    .D(_00719_),
    .Q(\count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_122_clk),
    .D(_00720_),
    .Q(\count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_122_clk),
    .D(_00721_),
    .Q(\count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_129_clk),
    .D(_00722_),
    .Q(\count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_129_clk),
    .D(_00723_),
    .Q(\count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_129_clk),
    .D(_00724_),
    .Q(\count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_84_clk),
    .D(_00725_),
    .Q(\count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_97_clk),
    .D(_00726_),
    .Q(\count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_97_clk),
    .D(_00727_),
    .Q(\count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_97_clk),
    .D(_00728_),
    .Q(\count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_97_clk),
    .D(_00729_),
    .Q(\count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_97_clk),
    .D(_00730_),
    .Q(\count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_98_clk),
    .D(_00731_),
    .Q(\count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_98_clk),
    .D(_00732_),
    .Q(\count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_98_clk),
    .D(_00733_),
    .Q(\count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_100_clk),
    .D(_00734_),
    .Q(\count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_100_clk),
    .D(_00735_),
    .Q(\count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_100_clk),
    .D(_00736_),
    .Q(\count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_96_clk),
    .D(_00737_),
    .Q(\count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_97_clk),
    .D(_00738_),
    .Q(\count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_97_clk),
    .D(_00739_),
    .Q(\count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_97_clk),
    .D(_00740_),
    .Q(\count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_84_clk),
    .D(_00741_),
    .Q(\count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_83_clk),
    .D(_00742_),
    .Q(\count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_126_clk),
    .D(_00743_),
    .Q(\count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_127_clk),
    .D(_00744_),
    .Q(\count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_128_clk),
    .D(_00745_),
    .Q(\count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_128_clk),
    .D(_00746_),
    .Q(\count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_123_clk),
    .D(_00747_),
    .Q(\count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_123_clk),
    .D(_00748_),
    .Q(\count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_123_clk),
    .D(_00749_),
    .Q(\count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_123_clk),
    .D(_00750_),
    .Q(\count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_124_clk),
    .D(_00751_),
    .Q(\count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_125_clk),
    .D(_00752_),
    .Q(\count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_126_clk),
    .D(_00753_),
    .Q(\count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_126_clk),
    .D(_00754_),
    .Q(\count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_126_clk),
    .D(_00755_),
    .Q(\count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_leaf_110_clk),
    .D(_00756_),
    .Q(\count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_110_clk),
    .D(_00757_),
    .Q(\count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_110_clk),
    .D(_00758_),
    .Q(\count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_110_clk),
    .D(_00759_),
    .Q(\count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_98_clk),
    .D(_00760_),
    .Q(\count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_98_clk),
    .D(_00761_),
    .Q(\count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_1 _14308_ (.CLK(clknet_leaf_98_clk),
    .D(_00762_),
    .Q(\count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_101_clk),
    .D(_00763_),
    .Q(\count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_101_clk),
    .D(_00764_),
    .Q(\count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_101_clk),
    .D(_00765_),
    .Q(\count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.CLK(clknet_leaf_101_clk),
    .D(_00766_),
    .Q(\count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_101_clk),
    .D(_00767_),
    .Q(\count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_101_clk),
    .D(_00768_),
    .Q(\count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_101_clk),
    .D(_00769_),
    .Q(\count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.CLK(clknet_leaf_93_clk),
    .D(_00770_),
    .Q(\count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_94_clk),
    .D(_00771_),
    .Q(\count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_93_clk),
    .D(_00772_),
    .Q(\count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.CLK(clknet_leaf_86_clk),
    .D(_00773_),
    .Q(net227));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.CLK(clknet_leaf_128_clk),
    .D(_06716_),
    .Q(\reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_131_clk),
    .D(_06727_),
    .Q(\reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_130_clk),
    .D(_06738_),
    .Q(\reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_133_clk),
    .D(_06741_),
    .Q(\reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_130_clk),
    .D(_06742_),
    .Q(\reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_134_clk),
    .D(_06743_),
    .Q(\reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_174_clk),
    .D(_06744_),
    .Q(\reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_174_clk),
    .D(_06745_),
    .Q(\reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_172_clk),
    .D(_06746_),
    .Q(\reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_171_clk),
    .D(_06747_),
    .Q(\reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_173_clk),
    .D(_06717_),
    .Q(\reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_177_clk),
    .D(_06718_),
    .Q(\reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_178_clk),
    .D(_06719_),
    .Q(\reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_177_clk),
    .D(_06720_),
    .Q(\reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_177_clk),
    .D(_06721_),
    .Q(\reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_176_clk),
    .D(_06722_),
    .Q(\reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_175_clk),
    .D(_06723_),
    .Q(\reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_26_clk),
    .D(_06724_),
    .Q(\reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14338_ (.CLK(clknet_leaf_27_clk),
    .D(_06725_),
    .Q(\reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.CLK(clknet_leaf_27_clk),
    .D(_06726_),
    .Q(\reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.CLK(clknet_leaf_76_clk),
    .D(_06728_),
    .Q(\reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_76_clk),
    .D(_06729_),
    .Q(\reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_76_clk),
    .D(_06730_),
    .Q(\reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.CLK(clknet_leaf_75_clk),
    .D(_06731_),
    .Q(\reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.CLK(clknet_leaf_82_clk),
    .D(_06732_),
    .Q(\reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14345_ (.CLK(clknet_leaf_82_clk),
    .D(_06733_),
    .Q(\reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_68_clk),
    .D(_06734_),
    .Q(\reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_67_clk),
    .D(_06735_),
    .Q(\reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_68_clk),
    .D(_06736_),
    .Q(\reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.CLK(clknet_leaf_66_clk),
    .D(_06737_),
    .Q(\reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.CLK(clknet_leaf_67_clk),
    .D(_06739_),
    .Q(\reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.CLK(clknet_leaf_87_clk),
    .D(_06740_),
    .Q(\reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.CLK(clknet_leaf_109_clk),
    .D(_00774_),
    .Q(\genblk2.pcpi_div.divisor[62] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_85_clk),
    .D(_00775_),
    .Q(mem_do_prefetch));
 sky130_fd_sc_hd__dfxtp_2 _14354_ (.CLK(clknet_leaf_85_clk),
    .D(_00776_),
    .Q(mem_do_rinst));
 sky130_fd_sc_hd__dfxtp_2 _14355_ (.CLK(clknet_leaf_85_clk),
    .D(_00777_),
    .Q(mem_do_rdata));
 sky130_fd_sc_hd__dfxtp_2 _14356_ (.CLK(clknet_leaf_85_clk),
    .D(_00778_),
    .Q(mem_do_wdata));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_87_clk),
    .D(_00000_),
    .Q(decoder_trigger));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_131_clk),
    .D(_00779_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_80_clk),
    .D(_00780_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_2 _14360_ (.CLK(clknet_leaf_80_clk),
    .D(_00781_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_2 _14361_ (.CLK(clknet_leaf_131_clk),
    .D(_00782_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_82_clk),
    .D(_00783_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_133_clk),
    .D(_00784_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_2 _14364_ (.CLK(clknet_leaf_136_clk),
    .D(_00785_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_171_clk),
    .D(_00786_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_2 _14366_ (.CLK(clknet_leaf_170_clk),
    .D(_00787_),
    .Q(net265));
 sky130_fd_sc_hd__dfxtp_2 _14367_ (.CLK(clknet_leaf_169_clk),
    .D(_00788_),
    .Q(net266));
 sky130_fd_sc_hd__dfxtp_4 _14368_ (.CLK(clknet_leaf_172_clk),
    .D(_00789_),
    .Q(net236));
 sky130_fd_sc_hd__dfxtp_2 _14369_ (.CLK(clknet_4_4_0_clk),
    .D(_00790_),
    .Q(net237));
 sky130_fd_sc_hd__dfxtp_4 _14370_ (.CLK(clknet_leaf_167_clk),
    .D(_00791_),
    .Q(net238));
 sky130_fd_sc_hd__dfxtp_4 _14371_ (.CLK(clknet_leaf_167_clk),
    .D(_00792_),
    .Q(net239));
 sky130_fd_sc_hd__dfxtp_4 _14372_ (.CLK(clknet_leaf_136_clk),
    .D(_00793_),
    .Q(net240));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_171_clk),
    .D(_00794_),
    .Q(net241));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_136_clk),
    .D(_00795_),
    .Q(net242));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_134_clk),
    .D(_00796_),
    .Q(net243));
 sky130_fd_sc_hd__dfxtp_4 _14376_ (.CLK(clknet_leaf_132_clk),
    .D(_00797_),
    .Q(net244));
 sky130_fd_sc_hd__dfxtp_2 _14377_ (.CLK(clknet_leaf_78_clk),
    .D(_00798_),
    .Q(net245));
 sky130_fd_sc_hd__dfxtp_2 _14378_ (.CLK(clknet_leaf_131_clk),
    .D(_00799_),
    .Q(net247));
 sky130_fd_sc_hd__dfxtp_4 _14379_ (.CLK(clknet_leaf_131_clk),
    .D(_00800_),
    .Q(net248));
 sky130_fd_sc_hd__dfxtp_4 _14380_ (.CLK(clknet_leaf_79_clk),
    .D(_00801_),
    .Q(net249));
 sky130_fd_sc_hd__dfxtp_4 _14381_ (.CLK(clknet_leaf_128_clk),
    .D(_00802_),
    .Q(net250));
 sky130_fd_sc_hd__dfxtp_2 _14382_ (.CLK(clknet_leaf_83_clk),
    .D(_00803_),
    .Q(net251));
 sky130_fd_sc_hd__dfxtp_2 _14383_ (.CLK(clknet_leaf_83_clk),
    .D(_00804_),
    .Q(net252));
 sky130_fd_sc_hd__dfxtp_4 _14384_ (.CLK(clknet_leaf_84_clk),
    .D(_00805_),
    .Q(net253));
 sky130_fd_sc_hd__dfxtp_2 _14385_ (.CLK(clknet_leaf_84_clk),
    .D(_00806_),
    .Q(net254));
 sky130_fd_sc_hd__dfxtp_2 _14386_ (.CLK(clknet_leaf_85_clk),
    .D(_00807_),
    .Q(net255));
 sky130_fd_sc_hd__dfxtp_2 _14387_ (.CLK(clknet_leaf_84_clk),
    .D(_00808_),
    .Q(net256));
 sky130_fd_sc_hd__dfxtp_4 _14388_ (.CLK(clknet_leaf_85_clk),
    .D(_00809_),
    .Q(net258));
 sky130_fd_sc_hd__dfxtp_1 _14389_ (.CLK(clknet_leaf_84_clk),
    .D(_00810_),
    .Q(net259));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.CLK(clknet_leaf_87_clk),
    .D(_00811_),
    .Q(latched_store));
 sky130_fd_sc_hd__dfxtp_1 _14391_ (.CLK(clknet_leaf_86_clk),
    .D(_00812_),
    .Q(latched_stalu));
 sky130_fd_sc_hd__dfxtp_1 _14392_ (.CLK(clknet_leaf_86_clk),
    .D(_00813_),
    .Q(latched_branch));
 sky130_fd_sc_hd__dfxtp_1 _14393_ (.CLK(clknet_leaf_87_clk),
    .D(_00814_),
    .Q(decoder_pseudo_trigger));
 sky130_fd_sc_hd__dfxtp_1 _14394_ (.CLK(clknet_leaf_85_clk),
    .D(_00815_),
    .Q(latched_is_lh));
 sky130_fd_sc_hd__dfxtp_1 _14395_ (.CLK(clknet_leaf_84_clk),
    .D(_00816_),
    .Q(latched_is_lb));
 sky130_fd_sc_hd__dfxtp_1 _14396_ (.CLK(clknet_leaf_102_clk),
    .D(_00817_),
    .Q(\pcpi_timeout_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14397_ (.CLK(clknet_leaf_102_clk),
    .D(_00818_),
    .Q(\pcpi_timeout_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14398_ (.CLK(clknet_leaf_99_clk),
    .D(_00819_),
    .Q(\pcpi_timeout_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14399_ (.CLK(clknet_leaf_99_clk),
    .D(_00820_),
    .Q(\pcpi_timeout_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14400_ (.CLK(clknet_leaf_127_clk),
    .D(\alu_out[0] ),
    .Q(\alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14401_ (.CLK(clknet_leaf_131_clk),
    .D(\alu_out[1] ),
    .Q(\alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14402_ (.CLK(clknet_leaf_130_clk),
    .D(\alu_out[2] ),
    .Q(\alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.CLK(clknet_leaf_134_clk),
    .D(\alu_out[3] ),
    .Q(\alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.CLK(clknet_leaf_134_clk),
    .D(\alu_out[4] ),
    .Q(\alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.CLK(clknet_leaf_135_clk),
    .D(\alu_out[5] ),
    .Q(\alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.CLK(clknet_leaf_136_clk),
    .D(\alu_out[6] ),
    .Q(\alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.CLK(clknet_leaf_136_clk),
    .D(\alu_out[7] ),
    .Q(\alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.CLK(clknet_leaf_171_clk),
    .D(\alu_out[8] ),
    .Q(\alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.CLK(clknet_leaf_170_clk),
    .D(\alu_out[9] ),
    .Q(\alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14410_ (.CLK(clknet_leaf_171_clk),
    .D(\alu_out[10] ),
    .Q(\alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.CLK(clknet_leaf_177_clk),
    .D(\alu_out[11] ),
    .Q(\alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.CLK(clknet_leaf_178_clk),
    .D(\alu_out[12] ),
    .Q(\alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.CLK(clknet_leaf_177_clk),
    .D(\alu_out[13] ),
    .Q(\alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.CLK(clknet_leaf_177_clk),
    .D(\alu_out[14] ),
    .Q(\alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_176_clk),
    .D(\alu_out[15] ),
    .Q(\alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_175_clk),
    .D(\alu_out[16] ),
    .Q(\alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.CLK(clknet_leaf_26_clk),
    .D(\alu_out[17] ),
    .Q(\alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.CLK(clknet_leaf_77_clk),
    .D(\alu_out[18] ),
    .Q(\alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.CLK(clknet_leaf_27_clk),
    .D(\alu_out[19] ),
    .Q(\alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.CLK(clknet_leaf_77_clk),
    .D(\alu_out[20] ),
    .Q(\alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.CLK(clknet_leaf_76_clk),
    .D(\alu_out[21] ),
    .Q(\alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.CLK(clknet_leaf_76_clk),
    .D(\alu_out[22] ),
    .Q(\alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_76_clk),
    .D(\alu_out[23] ),
    .Q(\alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_83_clk),
    .D(\alu_out[24] ),
    .Q(\alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_83_clk),
    .D(\alu_out[25] ),
    .Q(\alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.CLK(clknet_leaf_67_clk),
    .D(\alu_out[26] ),
    .Q(\alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.CLK(clknet_leaf_67_clk),
    .D(\alu_out[27] ),
    .Q(\alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.CLK(clknet_leaf_67_clk),
    .D(\alu_out[28] ),
    .Q(\alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.CLK(clknet_leaf_67_clk),
    .D(\alu_out[29] ),
    .Q(\alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14430_ (.CLK(clknet_leaf_67_clk),
    .D(\alu_out[30] ),
    .Q(\alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.CLK(clknet_leaf_87_clk),
    .D(\alu_out[31] ),
    .Q(\alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.CLK(clknet_leaf_100_clk),
    .D(_00821_),
    .Q(pcpi_timeout));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_91_clk),
    .D(net2555),
    .Q(net171));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.CLK(clknet_leaf_91_clk),
    .D(_00823_),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_65_clk),
    .D(_00824_),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.CLK(clknet_leaf_89_clk),
    .D(net2613),
    .Q(net196));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_64_clk),
    .D(net2637),
    .Q(net197));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_64_clk),
    .D(net2981),
    .Q(net198));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_64_clk),
    .D(net2738),
    .Q(net199));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.CLK(clknet_leaf_64_clk),
    .D(_00829_),
    .Q(net200));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_64_clk),
    .D(_00830_),
    .Q(net201));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_89_clk),
    .D(_00831_),
    .Q(net202));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_90_clk),
    .D(_00832_),
    .Q(net172));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_90_clk),
    .D(_00833_),
    .Q(net173));
 sky130_fd_sc_hd__dfxtp_2 _14445_ (.CLK(clknet_leaf_98_clk),
    .D(_00834_),
    .Q(net174));
 sky130_fd_sc_hd__dfxtp_2 _14446_ (.CLK(clknet_leaf_98_clk),
    .D(_00835_),
    .Q(net175));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_98_clk),
    .D(_00836_),
    .Q(net176));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_42_clk),
    .D(_00837_),
    .Q(net177));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_55_clk),
    .D(_00838_),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_55_clk),
    .D(_00839_),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.CLK(clknet_4_11_0_clk),
    .D(_00840_),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.CLK(clknet_leaf_64_clk),
    .D(_00841_),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.CLK(clknet_leaf_64_clk),
    .D(_00842_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_55_clk),
    .D(_00843_),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_64_clk),
    .D(_00844_),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_90_clk),
    .D(_00845_),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_90_clk),
    .D(_00846_),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_64_clk),
    .D(_00847_),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_64_clk),
    .D(_00848_),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_65_clk),
    .D(_00849_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_65_clk),
    .D(_00850_),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_64_clk),
    .D(_00851_),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_64_clk),
    .D(_00852_),
    .Q(net194));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_64_clk),
    .D(_00853_),
    .Q(net195));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_89_clk),
    .D(_00854_),
    .Q(instr_lui));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_89_clk),
    .D(_00855_),
    .Q(instr_auipc));
 sky130_fd_sc_hd__dfxtp_2 _14467_ (.CLK(clknet_leaf_89_clk),
    .D(_00856_),
    .Q(instr_jal));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_93_clk),
    .D(_00857_),
    .Q(instr_beq));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_95_clk),
    .D(_00858_),
    .Q(instr_bne));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_95_clk),
    .D(_00859_),
    .Q(instr_blt));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_95_clk),
    .D(_00860_),
    .Q(instr_bge));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_95_clk),
    .D(_00861_),
    .Q(instr_bltu));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_94_clk),
    .D(_00862_),
    .Q(instr_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _14474_ (.CLK(clknet_leaf_88_clk),
    .D(_00863_),
    .Q(instr_jalr));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_96_clk),
    .D(_00864_),
    .Q(instr_lb));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_95_clk),
    .D(_00865_),
    .Q(instr_lh));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_95_clk),
    .D(_00866_),
    .Q(instr_lw));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_96_clk),
    .D(_00867_),
    .Q(instr_lbu));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_96_clk),
    .D(_00868_),
    .Q(instr_lhu));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_96_clk),
    .D(_00869_),
    .Q(instr_sb));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_95_clk),
    .D(_00870_),
    .Q(instr_sh));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_93_clk),
    .D(_00871_),
    .Q(instr_addi));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_94_clk),
    .D(_00872_),
    .Q(instr_slti));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_95_clk),
    .D(_00873_),
    .Q(instr_sltiu));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_95_clk),
    .D(_00874_),
    .Q(instr_xori));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_95_clk),
    .D(_00875_),
    .Q(instr_ori));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_94_clk),
    .D(_00876_),
    .Q(instr_andi));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_95_clk),
    .D(_00877_),
    .Q(instr_sw));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.CLK(clknet_leaf_92_clk),
    .D(_00878_),
    .Q(instr_slli));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.CLK(clknet_leaf_92_clk),
    .D(_00879_),
    .Q(instr_srli));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.CLK(clknet_leaf_93_clk),
    .D(_00880_),
    .Q(instr_add));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_93_clk),
    .D(_00881_),
    .Q(instr_sub));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_95_clk),
    .D(_00882_),
    .Q(instr_sll));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_94_clk),
    .D(_00883_),
    .Q(instr_slt));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_94_clk),
    .D(_00884_),
    .Q(instr_sltu));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_95_clk),
    .D(_00885_),
    .Q(instr_xor));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_95_clk),
    .D(_00886_),
    .Q(instr_srl));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_93_clk),
    .D(_00887_),
    .Q(instr_sra));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_96_clk),
    .D(_00888_),
    .Q(instr_or));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_94_clk),
    .D(_00889_),
    .Q(instr_and));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_93_clk),
    .D(_00890_),
    .Q(instr_srai));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_91_clk),
    .D(_00891_),
    .Q(instr_rdcycle));
 sky130_fd_sc_hd__dfxtp_2 _14503_ (.CLK(clknet_leaf_91_clk),
    .D(_00892_),
    .Q(instr_rdcycleh));
 sky130_fd_sc_hd__dfxtp_2 _14504_ (.CLK(clknet_leaf_91_clk),
    .D(_00893_),
    .Q(instr_rdinstr));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_91_clk),
    .D(_00894_),
    .Q(instr_rdinstrh));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_93_clk),
    .D(_00895_),
    .Q(instr_fence));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_92_clk),
    .D(_00896_),
    .Q(instr_ecall_ebreak));
 sky130_fd_sc_hd__dfxtp_2 _14508_ (.CLK(clknet_leaf_80_clk),
    .D(_00897_),
    .Q(\decoded_imm_j[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_80_clk),
    .D(_00898_),
    .Q(\decoded_imm_j[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_80_clk),
    .D(_00899_),
    .Q(\decoded_imm_j[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_80_clk),
    .D(_00900_),
    .Q(\decoded_imm_j[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_78_clk),
    .D(_00901_),
    .Q(\decoded_imm_j[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_79_clk),
    .D(_00902_),
    .Q(\decoded_imm_j[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_79_clk),
    .D(_00903_),
    .Q(\decoded_imm_j[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_77_clk),
    .D(_00904_),
    .Q(\decoded_imm_j[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_77_clk),
    .D(_00905_),
    .Q(\decoded_imm_j[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_77_clk),
    .D(_00906_),
    .Q(\decoded_imm_j[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_28_clk),
    .D(_00907_),
    .Q(\decoded_imm_j[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_65_clk),
    .D(_00908_),
    .Q(\decoded_imm_j[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_69_clk),
    .D(_00909_),
    .Q(\decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_69_clk),
    .D(_00910_),
    .Q(\decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_69_clk),
    .D(_00911_),
    .Q(\decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_69_clk),
    .D(_00912_),
    .Q(\decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_69_clk),
    .D(_00913_),
    .Q(\decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_76_clk),
    .D(_00914_),
    .Q(\decoded_imm_j[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_28_clk),
    .D(_00915_),
    .Q(\decoded_imm_j[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_28_clk),
    .D(_00916_),
    .Q(\decoded_imm_j[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_28_clk),
    .D(_00917_),
    .Q(\decoded_imm_j[18] ));
 sky130_fd_sc_hd__dfxtp_2 _14529_ (.CLK(clknet_leaf_80_clk),
    .D(_00918_),
    .Q(\decoded_imm_j[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14530_ (.CLK(clknet_leaf_73_clk),
    .D(_00919_),
    .Q(\decoded_imm_j[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14531_ (.CLK(clknet_leaf_73_clk),
    .D(_00920_),
    .Q(\decoded_imm_j[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14532_ (.CLK(clknet_leaf_81_clk),
    .D(_00921_),
    .Q(\decoded_imm_j[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14533_ (.CLK(clknet_leaf_82_clk),
    .D(_00922_),
    .Q(\decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14534_ (.CLK(clknet_leaf_87_clk),
    .D(_00001_),
    .Q(is_lui_auipc_jal));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_88_clk),
    .D(_00923_),
    .Q(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_92_clk),
    .D(net2672),
    .Q(is_slli_srli_srai));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_88_clk),
    .D(_00925_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
 sky130_fd_sc_hd__dfxtp_2 _14538_ (.CLK(clknet_leaf_88_clk),
    .D(_00926_),
    .Q(is_sb_sh_sw));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_91_clk),
    .D(_00927_),
    .Q(is_sll_srl_sra));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_96_clk),
    .D(net2655),
    .Q(is_slti_blt_slt));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_96_clk),
    .D(_00003_),
    .Q(is_sltiu_bltu_sltu));
 sky130_fd_sc_hd__dfxtp_2 _14542_ (.CLK(clknet_leaf_88_clk),
    .D(_00928_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_39_clk),
    .D(_00929_),
    .Q(\cpuregs[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_46_clk),
    .D(_00930_),
    .Q(\cpuregs[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_73_clk),
    .D(_00931_),
    .Q(\cpuregs[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_21_clk),
    .D(_00932_),
    .Q(\cpuregs[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_24_clk),
    .D(_00933_),
    .Q(\cpuregs[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_24_clk),
    .D(_00934_),
    .Q(\cpuregs[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_179_clk),
    .D(_00935_),
    .Q(\cpuregs[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_187_clk),
    .D(_00936_),
    .Q(\cpuregs[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_184_clk),
    .D(_00937_),
    .Q(\cpuregs[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_184_clk),
    .D(_00938_),
    .Q(\cpuregs[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_187_clk),
    .D(_00939_),
    .Q(\cpuregs[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_192_clk),
    .D(_00940_),
    .Q(\cpuregs[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_3_clk),
    .D(_00941_),
    .Q(\cpuregs[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_195_clk),
    .D(_00942_),
    .Q(\cpuregs[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_195_clk),
    .D(_00943_),
    .Q(\cpuregs[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_199_clk),
    .D(_00944_),
    .Q(\cpuregs[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_11_clk),
    .D(_00945_),
    .Q(\cpuregs[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_0_clk),
    .D(_00946_),
    .Q(\cpuregs[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_1_clk),
    .D(_00947_),
    .Q(\cpuregs[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_41_clk),
    .D(_00948_),
    .Q(\cpuregs[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_14_clk),
    .D(_00949_),
    .Q(\cpuregs[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_13_clk),
    .D(_00950_),
    .Q(\cpuregs[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_43_clk),
    .D(_00951_),
    .Q(\cpuregs[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_37_clk),
    .D(_00952_),
    .Q(\cpuregs[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_31_clk),
    .D(_00953_),
    .Q(\cpuregs[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_60_clk),
    .D(_00954_),
    .Q(\cpuregs[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_57_clk),
    .D(_00955_),
    .Q(\cpuregs[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_56_clk),
    .D(_00956_),
    .Q(\cpuregs[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_51_clk),
    .D(_00957_),
    .Q(\cpuregs[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_69_clk),
    .D(_00958_),
    .Q(\cpuregs[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_54_clk),
    .D(_00959_),
    .Q(\cpuregs[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_50_clk),
    .D(_00960_),
    .Q(\cpuregs[27][31] ));
 sky130_fd_sc_hd__dfxtp_2 _14575_ (.CLK(clknet_leaf_89_clk),
    .D(_00961_),
    .Q(is_alu_reg_imm));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_88_clk),
    .D(_00962_),
    .Q(is_alu_reg_reg));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_96_clk),
    .D(_00963_),
    .Q(is_compare));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_93_clk),
    .D(_00964_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_2 _14579_ (.CLK(clknet_leaf_69_clk),
    .D(_00965_),
    .Q(\latched_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _14580_ (.CLK(clknet_leaf_69_clk),
    .D(net1466),
    .Q(\latched_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _14581_ (.CLK(clknet_leaf_69_clk),
    .D(_00967_),
    .Q(\latched_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _14582_ (.CLK(clknet_leaf_69_clk),
    .D(_00968_),
    .Q(\latched_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14583_ (.CLK(clknet_leaf_69_clk),
    .D(_00969_),
    .Q(\latched_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_117_clk),
    .D(_00970_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_104_clk),
    .D(_00971_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.CLK(clknet_leaf_115_clk),
    .D(_00972_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_114_clk),
    .D(net1877),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.CLK(clknet_leaf_104_clk),
    .D(_00974_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_106_clk),
    .D(_00975_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_114_clk),
    .D(_00976_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_104_clk),
    .D(_00977_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_159_clk),
    .D(_00978_),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_156_clk),
    .D(_00979_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_115_clk),
    .D(_00980_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_159_clk),
    .D(_00981_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_159_clk),
    .D(_00982_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.CLK(clknet_leaf_115_clk),
    .D(_00983_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.CLK(clknet_leaf_117_clk),
    .D(_00984_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_115_clk),
    .D(_00985_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_118_clk),
    .D(_00986_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.CLK(clknet_leaf_145_clk),
    .D(_00987_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_156_clk),
    .D(_00988_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_117_clk),
    .D(_00989_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_118_clk),
    .D(_00990_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_118_clk),
    .D(_00991_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_156_clk),
    .D(_00992_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.CLK(clknet_leaf_114_clk),
    .D(_00993_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.CLK(clknet_leaf_104_clk),
    .D(_00994_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_104_clk),
    .D(_00995_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_106_clk),
    .D(_00996_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_106_clk),
    .D(_00997_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_104_clk),
    .D(_00998_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.CLK(clknet_leaf_104_clk),
    .D(_00999_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.CLK(clknet_leaf_114_clk),
    .D(_01000_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_115_clk),
    .D(_01001_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_93_clk),
    .D(_01002_),
    .Q(net167));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_93_clk),
    .D(_01003_),
    .Q(net168));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_117_clk),
    .D(_01004_),
    .Q(net169));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_107_clk),
    .D(_01005_),
    .Q(net170));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_93_clk),
    .D(_01006_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_109_clk),
    .D(_01007_),
    .Q(\genblk2.pcpi_div.instr_div ));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.CLK(clknet_leaf_108_clk),
    .D(_01008_),
    .Q(\genblk2.pcpi_div.outsign ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_109_clk),
    .D(net1371),
    .Q(\genblk2.pcpi_div.pcpi_wait ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_122_clk),
    .D(_01009_),
    .Q(\genblk2.pcpi_div.dividend[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_129_clk),
    .D(_01010_),
    .Q(\genblk2.pcpi_div.dividend[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_135_clk),
    .D(_01011_),
    .Q(\genblk2.pcpi_div.dividend[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_135_clk),
    .D(_01012_),
    .Q(\genblk2.pcpi_div.dividend[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_135_clk),
    .D(_01013_),
    .Q(\genblk2.pcpi_div.dividend[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_139_clk),
    .D(_01014_),
    .Q(\genblk2.pcpi_div.dividend[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_137_clk),
    .D(_01015_),
    .Q(\genblk2.pcpi_div.dividend[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.CLK(clknet_leaf_137_clk),
    .D(_01016_),
    .Q(\genblk2.pcpi_div.dividend[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_170_clk),
    .D(_01017_),
    .Q(\genblk2.pcpi_div.dividend[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_170_clk),
    .D(_01018_),
    .Q(\genblk2.pcpi_div.dividend[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_170_clk),
    .D(_01019_),
    .Q(\genblk2.pcpi_div.dividend[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_169_clk),
    .D(_01020_),
    .Q(\genblk2.pcpi_div.dividend[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_169_clk),
    .D(_01021_),
    .Q(\genblk2.pcpi_div.dividend[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_163_clk),
    .D(_01022_),
    .Q(\genblk2.pcpi_div.dividend[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14638_ (.CLK(clknet_leaf_169_clk),
    .D(_01023_),
    .Q(\genblk2.pcpi_div.dividend[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_164_clk),
    .D(_01024_),
    .Q(\genblk2.pcpi_div.dividend[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_164_clk),
    .D(_01025_),
    .Q(\genblk2.pcpi_div.dividend[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.CLK(clknet_leaf_165_clk),
    .D(_01026_),
    .Q(\genblk2.pcpi_div.dividend[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_165_clk),
    .D(_01027_),
    .Q(\genblk2.pcpi_div.dividend[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_161_clk),
    .D(_01028_),
    .Q(\genblk2.pcpi_div.dividend[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_161_clk),
    .D(_01029_),
    .Q(\genblk2.pcpi_div.dividend[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.CLK(clknet_leaf_161_clk),
    .D(_01030_),
    .Q(\genblk2.pcpi_div.dividend[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.CLK(clknet_leaf_161_clk),
    .D(_01031_),
    .Q(\genblk2.pcpi_div.dividend[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_161_clk),
    .D(_01032_),
    .Q(\genblk2.pcpi_div.dividend[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_160_clk),
    .D(_01033_),
    .Q(\genblk2.pcpi_div.dividend[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_158_clk),
    .D(_01034_),
    .Q(\genblk2.pcpi_div.dividend[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_157_clk),
    .D(_01035_),
    .Q(\genblk2.pcpi_div.dividend[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_157_clk),
    .D(_01036_),
    .Q(\genblk2.pcpi_div.dividend[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_155_clk),
    .D(_01037_),
    .Q(\genblk2.pcpi_div.dividend[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_153_clk),
    .D(_01038_),
    .Q(\genblk2.pcpi_div.dividend[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_155_clk),
    .D(_01039_),
    .Q(\genblk2.pcpi_div.dividend[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_150_clk),
    .D(_01040_),
    .Q(\genblk2.pcpi_div.dividend[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_153_clk),
    .D(_01041_),
    .Q(\genblk2.pcpi_div.running ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_143_clk),
    .D(net2603),
    .Q(\genblk2.pcpi_div.quotient_msk[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_141_clk),
    .D(net2751),
    .Q(\genblk2.pcpi_div.quotient_msk[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_141_clk),
    .D(_01044_),
    .Q(\genblk2.pcpi_div.quotient_msk[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_139_clk),
    .D(_01045_),
    .Q(\genblk2.pcpi_div.quotient_msk[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_152_clk),
    .D(net2530),
    .Q(\genblk2.pcpi_div.quotient_msk[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_138_clk),
    .D(_01047_),
    .Q(\genblk2.pcpi_div.quotient_msk[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_151_clk),
    .D(_01048_),
    .Q(\genblk2.pcpi_div.quotient_msk[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_152_clk),
    .D(_01049_),
    .Q(\genblk2.pcpi_div.quotient_msk[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_152_clk),
    .D(net2757),
    .Q(\genblk2.pcpi_div.quotient_msk[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_152_clk),
    .D(_01051_),
    .Q(\genblk2.pcpi_div.quotient_msk[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_152_clk),
    .D(_01052_),
    .Q(\genblk2.pcpi_div.quotient_msk[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_152_clk),
    .D(net2804),
    .Q(\genblk2.pcpi_div.quotient_msk[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_153_clk),
    .D(_01054_),
    .Q(\genblk2.pcpi_div.quotient_msk[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_153_clk),
    .D(_01055_),
    .Q(\genblk2.pcpi_div.quotient_msk[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_153_clk),
    .D(net2786),
    .Q(\genblk2.pcpi_div.quotient_msk[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_162_clk),
    .D(net2777),
    .Q(\genblk2.pcpi_div.quotient_msk[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_162_clk),
    .D(_01058_),
    .Q(\genblk2.pcpi_div.quotient_msk[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_162_clk),
    .D(_01059_),
    .Q(\genblk2.pcpi_div.quotient_msk[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_162_clk),
    .D(net2840),
    .Q(\genblk2.pcpi_div.quotient_msk[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_162_clk),
    .D(net2795),
    .Q(\genblk2.pcpi_div.quotient_msk[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_162_clk),
    .D(_01062_),
    .Q(\genblk2.pcpi_div.quotient_msk[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_162_clk),
    .D(_01063_),
    .Q(\genblk2.pcpi_div.quotient_msk[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_153_clk),
    .D(_01064_),
    .Q(\genblk2.pcpi_div.quotient_msk[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_153_clk),
    .D(net2868),
    .Q(\genblk2.pcpi_div.quotient_msk[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_153_clk),
    .D(net2792),
    .Q(\genblk2.pcpi_div.quotient_msk[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_153_clk),
    .D(_01067_),
    .Q(\genblk2.pcpi_div.quotient_msk[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_153_clk),
    .D(_01068_),
    .Q(\genblk2.pcpi_div.quotient_msk[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_156_clk),
    .D(net2844),
    .Q(\genblk2.pcpi_div.quotient_msk[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_156_clk),
    .D(net2733),
    .Q(\genblk2.pcpi_div.quotient_msk[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_156_clk),
    .D(_01071_),
    .Q(\genblk2.pcpi_div.quotient_msk[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_155_clk),
    .D(_01072_),
    .Q(\genblk2.pcpi_div.quotient_msk[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_155_clk),
    .D(_01073_),
    .Q(\genblk2.pcpi_div.quotient_msk[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_143_clk),
    .D(_01074_),
    .Q(\genblk2.pcpi_div.quotient[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_142_clk),
    .D(_01075_),
    .Q(\genblk2.pcpi_div.quotient[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_141_clk),
    .D(_01076_),
    .Q(\genblk2.pcpi_div.quotient[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_141_clk),
    .D(_01077_),
    .Q(\genblk2.pcpi_div.quotient[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.CLK(clknet_leaf_139_clk),
    .D(_01078_),
    .Q(\genblk2.pcpi_div.quotient[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.CLK(clknet_leaf_138_clk),
    .D(_01079_),
    .Q(\genblk2.pcpi_div.quotient[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_138_clk),
    .D(_01080_),
    .Q(\genblk2.pcpi_div.quotient[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.CLK(clknet_leaf_152_clk),
    .D(_01081_),
    .Q(\genblk2.pcpi_div.quotient[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_152_clk),
    .D(_01082_),
    .Q(\genblk2.pcpi_div.quotient[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.CLK(clknet_leaf_152_clk),
    .D(_01083_),
    .Q(\genblk2.pcpi_div.quotient[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_152_clk),
    .D(_01084_),
    .Q(\genblk2.pcpi_div.quotient[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_152_clk),
    .D(_01085_),
    .Q(\genblk2.pcpi_div.quotient[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_163_clk),
    .D(_01086_),
    .Q(\genblk2.pcpi_div.quotient[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.CLK(clknet_leaf_153_clk),
    .D(_01087_),
    .Q(\genblk2.pcpi_div.quotient[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_153_clk),
    .D(_01088_),
    .Q(\genblk2.pcpi_div.quotient[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_153_clk),
    .D(_01089_),
    .Q(\genblk2.pcpi_div.quotient[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_162_clk),
    .D(_01090_),
    .Q(\genblk2.pcpi_div.quotient[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_162_clk),
    .D(_01091_),
    .Q(\genblk2.pcpi_div.quotient[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_162_clk),
    .D(_01092_),
    .Q(\genblk2.pcpi_div.quotient[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_162_clk),
    .D(_01093_),
    .Q(\genblk2.pcpi_div.quotient[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_162_clk),
    .D(_01094_),
    .Q(\genblk2.pcpi_div.quotient[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_162_clk),
    .D(_01095_),
    .Q(\genblk2.pcpi_div.quotient[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_153_clk),
    .D(_01096_),
    .Q(\genblk2.pcpi_div.quotient[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_162_clk),
    .D(_01097_),
    .Q(\genblk2.pcpi_div.quotient[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_154_clk),
    .D(_01098_),
    .Q(\genblk2.pcpi_div.quotient[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_153_clk),
    .D(_01099_),
    .Q(\genblk2.pcpi_div.quotient[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_154_clk),
    .D(_01100_),
    .Q(\genblk2.pcpi_div.quotient[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_156_clk),
    .D(_01101_),
    .Q(\genblk2.pcpi_div.quotient[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.CLK(clknet_leaf_156_clk),
    .D(_01102_),
    .Q(\genblk2.pcpi_div.quotient[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.CLK(clknet_leaf_156_clk),
    .D(_01103_),
    .Q(\genblk2.pcpi_div.quotient[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_155_clk),
    .D(_01104_),
    .Q(\genblk2.pcpi_div.quotient[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_155_clk),
    .D(_01105_),
    .Q(\genblk2.pcpi_div.quotient[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_142_clk),
    .D(net2580),
    .Q(\genblk2.pcpi_div.divisor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.CLK(clknet_leaf_142_clk),
    .D(net2965),
    .Q(\genblk2.pcpi_div.divisor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_141_clk),
    .D(net2899),
    .Q(\genblk2.pcpi_div.divisor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_141_clk),
    .D(net2718),
    .Q(\genblk2.pcpi_div.divisor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_141_clk),
    .D(_01110_),
    .Q(\genblk2.pcpi_div.divisor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_138_clk),
    .D(_01111_),
    .Q(\genblk2.pcpi_div.divisor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_138_clk),
    .D(net2716),
    .Q(\genblk2.pcpi_div.divisor[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_170_clk),
    .D(_01113_),
    .Q(\genblk2.pcpi_div.divisor[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14729_ (.CLK(clknet_leaf_170_clk),
    .D(_01114_),
    .Q(\genblk2.pcpi_div.divisor[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.CLK(clknet_leaf_170_clk),
    .D(_01115_),
    .Q(\genblk2.pcpi_div.divisor[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_170_clk),
    .D(_01116_),
    .Q(\genblk2.pcpi_div.divisor[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.CLK(clknet_leaf_163_clk),
    .D(net2705),
    .Q(\genblk2.pcpi_div.divisor[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_163_clk),
    .D(net2678),
    .Q(\genblk2.pcpi_div.divisor[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_164_clk),
    .D(_01119_),
    .Q(\genblk2.pcpi_div.divisor[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.CLK(clknet_leaf_164_clk),
    .D(_01120_),
    .Q(\genblk2.pcpi_div.divisor[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_164_clk),
    .D(_01121_),
    .Q(\genblk2.pcpi_div.divisor[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.CLK(clknet_leaf_165_clk),
    .D(_01122_),
    .Q(\genblk2.pcpi_div.divisor[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.CLK(clknet_leaf_165_clk),
    .D(net2770),
    .Q(\genblk2.pcpi_div.divisor[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_161_clk),
    .D(_01124_),
    .Q(\genblk2.pcpi_div.divisor[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14740_ (.CLK(clknet_leaf_161_clk),
    .D(_01125_),
    .Q(\genblk2.pcpi_div.divisor[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.CLK(clknet_leaf_160_clk),
    .D(_01126_),
    .Q(\genblk2.pcpi_div.divisor[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.CLK(clknet_leaf_160_clk),
    .D(_01127_),
    .Q(\genblk2.pcpi_div.divisor[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_160_clk),
    .D(_01128_),
    .Q(\genblk2.pcpi_div.divisor[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.CLK(clknet_leaf_160_clk),
    .D(net2693),
    .Q(\genblk2.pcpi_div.divisor[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_158_clk),
    .D(_01130_),
    .Q(\genblk2.pcpi_div.divisor[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_158_clk),
    .D(_01131_),
    .Q(\genblk2.pcpi_div.divisor[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_158_clk),
    .D(net2744),
    .Q(\genblk2.pcpi_div.divisor[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14748_ (.CLK(clknet_leaf_157_clk),
    .D(_01133_),
    .Q(\genblk2.pcpi_div.divisor[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.CLK(clknet_leaf_155_clk),
    .D(net2874),
    .Q(\genblk2.pcpi_div.divisor[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.CLK(clknet_leaf_153_clk),
    .D(_01135_),
    .Q(\genblk2.pcpi_div.divisor[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14751_ (.CLK(clknet_leaf_153_clk),
    .D(net2174),
    .Q(\genblk2.pcpi_div.divisor[30] ));
 sky130_fd_sc_hd__dfxtp_2 _14752_ (.CLK(clknet_leaf_152_clk),
    .D(_01137_),
    .Q(\genblk2.pcpi_div.pcpi_ready ));
 sky130_fd_sc_hd__dfxtp_1 _14753_ (.CLK(clknet_leaf_123_clk),
    .D(_00016_),
    .Q(\genblk2.pcpi_div.pcpi_rd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14754_ (.CLK(clknet_leaf_124_clk),
    .D(_00027_),
    .Q(\genblk2.pcpi_div.pcpi_rd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14755_ (.CLK(clknet_leaf_122_clk),
    .D(_00038_),
    .Q(\genblk2.pcpi_div.pcpi_rd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14756_ (.CLK(clknet_leaf_122_clk),
    .D(_00041_),
    .Q(\genblk2.pcpi_div.pcpi_rd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14757_ (.CLK(clknet_leaf_141_clk),
    .D(_00042_),
    .Q(\genblk2.pcpi_div.pcpi_rd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14758_ (.CLK(clknet_leaf_141_clk),
    .D(_00043_),
    .Q(\genblk2.pcpi_div.pcpi_rd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14759_ (.CLK(clknet_leaf_139_clk),
    .D(_00044_),
    .Q(\genblk2.pcpi_div.pcpi_rd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14760_ (.CLK(clknet_leaf_137_clk),
    .D(_00045_),
    .Q(\genblk2.pcpi_div.pcpi_rd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.CLK(clknet_leaf_137_clk),
    .D(_00046_),
    .Q(\genblk2.pcpi_div.pcpi_rd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14762_ (.CLK(clknet_leaf_137_clk),
    .D(_00047_),
    .Q(\genblk2.pcpi_div.pcpi_rd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.CLK(clknet_leaf_152_clk),
    .D(_00017_),
    .Q(\genblk2.pcpi_div.pcpi_rd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.CLK(clknet_leaf_170_clk),
    .D(_00018_),
    .Q(\genblk2.pcpi_div.pcpi_rd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.CLK(clknet_leaf_163_clk),
    .D(_00019_),
    .Q(\genblk2.pcpi_div.pcpi_rd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.CLK(clknet_leaf_163_clk),
    .D(_00020_),
    .Q(\genblk2.pcpi_div.pcpi_rd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.CLK(clknet_leaf_163_clk),
    .D(_00021_),
    .Q(\genblk2.pcpi_div.pcpi_rd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_163_clk),
    .D(_00022_),
    .Q(\genblk2.pcpi_div.pcpi_rd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_164_clk),
    .D(_00023_),
    .Q(\genblk2.pcpi_div.pcpi_rd[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_164_clk),
    .D(_00024_),
    .Q(\genblk2.pcpi_div.pcpi_rd[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_164_clk),
    .D(_00025_),
    .Q(\genblk2.pcpi_div.pcpi_rd[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_161_clk),
    .D(_00026_),
    .Q(\genblk2.pcpi_div.pcpi_rd[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_162_clk),
    .D(_00028_),
    .Q(\genblk2.pcpi_div.pcpi_rd[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_153_clk),
    .D(_00029_),
    .Q(\genblk2.pcpi_div.pcpi_rd[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14775_ (.CLK(clknet_leaf_153_clk),
    .D(_00030_),
    .Q(\genblk2.pcpi_div.pcpi_rd[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_154_clk),
    .D(_00031_),
    .Q(\genblk2.pcpi_div.pcpi_rd[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.CLK(clknet_leaf_154_clk),
    .D(_00032_),
    .Q(\genblk2.pcpi_div.pcpi_rd[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_154_clk),
    .D(_00033_),
    .Q(\genblk2.pcpi_div.pcpi_rd[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_154_clk),
    .D(_00034_),
    .Q(\genblk2.pcpi_div.pcpi_rd[26] ));
 sky130_fd_sc_hd__dfxtp_2 _14780_ (.CLK(clknet_leaf_157_clk),
    .D(_00035_),
    .Q(\genblk2.pcpi_div.pcpi_rd[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_155_clk),
    .D(_00036_),
    .Q(\genblk2.pcpi_div.pcpi_rd[28] ));
 sky130_fd_sc_hd__dfxtp_2 _14782_ (.CLK(clknet_leaf_155_clk),
    .D(_00037_),
    .Q(\genblk2.pcpi_div.pcpi_rd[29] ));
 sky130_fd_sc_hd__dfxtp_2 _14783_ (.CLK(clknet_leaf_149_clk),
    .D(_00039_),
    .Q(\genblk2.pcpi_div.pcpi_rd[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_149_clk),
    .D(_00040_),
    .Q(\genblk2.pcpi_div.pcpi_rd[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_98_clk),
    .D(_01138_),
    .Q(\genblk1.genblk1.pcpi_mul.instr_mulhu ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_91_clk),
    .D(_01139_),
    .Q(\mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.CLK(clknet_leaf_91_clk),
    .D(_01140_),
    .Q(\mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.CLK(clknet_leaf_109_clk),
    .D(_01141_),
    .Q(\genblk2.pcpi_div.instr_divu ));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.CLK(clknet_leaf_109_clk),
    .D(_01142_),
    .Q(\genblk2.pcpi_div.instr_rem ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_109_clk),
    .D(_00049_),
    .Q(\genblk2.pcpi_div.pcpi_wait_q ));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.CLK(clknet_leaf_67_clk),
    .D(_01143_),
    .Q(\decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.CLK(clknet_leaf_86_clk),
    .D(_01144_),
    .Q(\decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.CLK(clknet_leaf_67_clk),
    .D(_01145_),
    .Q(\decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.CLK(clknet_leaf_67_clk),
    .D(_01146_),
    .Q(\decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_67_clk),
    .D(_01147_),
    .Q(\decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.CLK(clknet_leaf_67_clk),
    .D(_01148_),
    .Q(\decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.CLK(clknet_leaf_75_clk),
    .D(_01149_),
    .Q(\decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.CLK(clknet_leaf_81_clk),
    .D(_01150_),
    .Q(\decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_2 _14799_ (.CLK(clknet_leaf_81_clk),
    .D(_01151_),
    .Q(\decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_75_clk),
    .D(_01152_),
    .Q(\decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_75_clk),
    .D(_01153_),
    .Q(\decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.CLK(clknet_leaf_75_clk),
    .D(_01154_),
    .Q(\decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_2 _14803_ (.CLK(clknet_leaf_77_clk),
    .D(_01155_),
    .Q(\decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_77_clk),
    .D(_01156_),
    .Q(\decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_2 _14805_ (.CLK(clknet_leaf_77_clk),
    .D(_01157_),
    .Q(\decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_2 _14806_ (.CLK(clknet_leaf_77_clk),
    .D(_01158_),
    .Q(\decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_2 _14807_ (.CLK(clknet_leaf_77_clk),
    .D(_01159_),
    .Q(\decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_2 _14808_ (.CLK(clknet_leaf_78_clk),
    .D(_01160_),
    .Q(\decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_2 _14809_ (.CLK(clknet_leaf_77_clk),
    .D(_01161_),
    .Q(\decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_2 _14810_ (.CLK(clknet_leaf_77_clk),
    .D(_01162_),
    .Q(\decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 _14811_ (.CLK(clknet_leaf_81_clk),
    .D(_01163_),
    .Q(\decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_2 _14812_ (.CLK(clknet_leaf_131_clk),
    .D(_01164_),
    .Q(\decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_2 _14813_ (.CLK(clknet_leaf_79_clk),
    .D(_01165_),
    .Q(\decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_2 _14814_ (.CLK(clknet_leaf_78_clk),
    .D(_01166_),
    .Q(\decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_2 _14815_ (.CLK(clknet_leaf_79_clk),
    .D(_01167_),
    .Q(\decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_2 _14816_ (.CLK(clknet_leaf_79_clk),
    .D(_01168_),
    .Q(\decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_2 _14817_ (.CLK(clknet_leaf_79_clk),
    .D(_01169_),
    .Q(\decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_2 _14818_ (.CLK(clknet_leaf_82_clk),
    .D(_01170_),
    .Q(\decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.CLK(clknet_leaf_82_clk),
    .D(_01171_),
    .Q(\decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_2 _14820_ (.CLK(clknet_leaf_82_clk),
    .D(_01172_),
    .Q(\decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_82_clk),
    .D(_01173_),
    .Q(\decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_105_clk),
    .D(_01174_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_39_clk),
    .D(_01175_),
    .Q(\cpuregs[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_46_clk),
    .D(_01176_),
    .Q(\cpuregs[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_32_clk),
    .D(_01177_),
    .Q(\cpuregs[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_21_clk),
    .D(_01178_),
    .Q(\cpuregs[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_23_clk),
    .D(_01179_),
    .Q(\cpuregs[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.CLK(clknet_leaf_24_clk),
    .D(_01180_),
    .Q(\cpuregs[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.CLK(clknet_leaf_179_clk),
    .D(_01181_),
    .Q(\cpuregs[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14830_ (.CLK(clknet_leaf_187_clk),
    .D(_01182_),
    .Q(\cpuregs[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14831_ (.CLK(clknet_leaf_184_clk),
    .D(_01183_),
    .Q(\cpuregs[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.CLK(clknet_leaf_184_clk),
    .D(_01184_),
    .Q(\cpuregs[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.CLK(clknet_leaf_187_clk),
    .D(_01185_),
    .Q(\cpuregs[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.CLK(clknet_leaf_192_clk),
    .D(_01186_),
    .Q(\cpuregs[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14835_ (.CLK(clknet_leaf_3_clk),
    .D(_01187_),
    .Q(\cpuregs[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.CLK(clknet_leaf_195_clk),
    .D(_01188_),
    .Q(\cpuregs[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.CLK(clknet_leaf_195_clk),
    .D(_01189_),
    .Q(\cpuregs[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_0_clk),
    .D(_01190_),
    .Q(\cpuregs[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.CLK(clknet_leaf_11_clk),
    .D(_01191_),
    .Q(\cpuregs[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_0_clk),
    .D(_01192_),
    .Q(\cpuregs[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_1_clk),
    .D(_01193_),
    .Q(\cpuregs[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_41_clk),
    .D(_01194_),
    .Q(\cpuregs[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14843_ (.CLK(clknet_leaf_11_clk),
    .D(_01195_),
    .Q(\cpuregs[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14844_ (.CLK(clknet_leaf_13_clk),
    .D(_01196_),
    .Q(\cpuregs[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14845_ (.CLK(clknet_leaf_43_clk),
    .D(_01197_),
    .Q(\cpuregs[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14846_ (.CLK(clknet_leaf_38_clk),
    .D(_01198_),
    .Q(\cpuregs[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14847_ (.CLK(clknet_leaf_31_clk),
    .D(_01199_),
    .Q(\cpuregs[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.CLK(clknet_leaf_60_clk),
    .D(_01200_),
    .Q(\cpuregs[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.CLK(clknet_leaf_57_clk),
    .D(_01201_),
    .Q(\cpuregs[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14850_ (.CLK(clknet_leaf_56_clk),
    .D(_01202_),
    .Q(\cpuregs[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14851_ (.CLK(clknet_leaf_51_clk),
    .D(_01203_),
    .Q(\cpuregs[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.CLK(clknet_leaf_69_clk),
    .D(_01204_),
    .Q(\cpuregs[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14853_ (.CLK(clknet_leaf_54_clk),
    .D(_01205_),
    .Q(\cpuregs[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14854_ (.CLK(clknet_leaf_50_clk),
    .D(_01206_),
    .Q(\cpuregs[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14855_ (.CLK(clknet_leaf_30_clk),
    .D(_01207_),
    .Q(\cpuregs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.CLK(clknet_leaf_48_clk),
    .D(_01208_),
    .Q(\cpuregs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.CLK(clknet_leaf_32_clk),
    .D(_01209_),
    .Q(\cpuregs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.CLK(clknet_leaf_17_clk),
    .D(_01210_),
    .Q(\cpuregs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.CLK(clknet_leaf_23_clk),
    .D(_01211_),
    .Q(\cpuregs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_23_clk),
    .D(_01212_),
    .Q(\cpuregs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_179_clk),
    .D(_01213_),
    .Q(\cpuregs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_19_clk),
    .D(_01214_),
    .Q(\cpuregs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.CLK(clknet_leaf_180_clk),
    .D(_01215_),
    .Q(\cpuregs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.CLK(clknet_leaf_182_clk),
    .D(_01216_),
    .Q(\cpuregs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.CLK(clknet_leaf_181_clk),
    .D(_01217_),
    .Q(\cpuregs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.CLK(clknet_leaf_20_clk),
    .D(_01218_),
    .Q(\cpuregs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.CLK(clknet_leaf_6_clk),
    .D(_01219_),
    .Q(\cpuregs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_6_clk),
    .D(_01220_),
    .Q(\cpuregs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_19_clk),
    .D(_01221_),
    .Q(\cpuregs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_7_clk),
    .D(_01222_),
    .Q(\cpuregs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_18_clk),
    .D(_01223_),
    .Q(\cpuregs[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_6_clk),
    .D(_01224_),
    .Q(\cpuregs[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_6_clk),
    .D(_01225_),
    .Q(\cpuregs[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_39_clk),
    .D(_01226_),
    .Q(\cpuregs[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_18_clk),
    .D(_01227_),
    .Q(\cpuregs[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.CLK(clknet_leaf_38_clk),
    .D(_01228_),
    .Q(\cpuregs[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.CLK(clknet_leaf_36_clk),
    .D(_01229_),
    .Q(\cpuregs[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.CLK(clknet_leaf_17_clk),
    .D(_01230_),
    .Q(\cpuregs[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.CLK(clknet_leaf_35_clk),
    .D(_01231_),
    .Q(\cpuregs[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_72_clk),
    .D(_01232_),
    .Q(\cpuregs[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_33_clk),
    .D(_01233_),
    .Q(\cpuregs[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_34_clk),
    .D(_01234_),
    .Q(\cpuregs[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_47_clk),
    .D(_01235_),
    .Q(\cpuregs[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_72_clk),
    .D(_01236_),
    .Q(\cpuregs[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_48_clk),
    .D(_01237_),
    .Q(\cpuregs[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_49_clk),
    .D(_01238_),
    .Q(\cpuregs[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_104_clk),
    .D(_01239_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_105_clk),
    .D(_01240_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_105_clk),
    .D(_01241_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_105_clk),
    .D(_01242_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_105_clk),
    .D(_01243_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_151_clk),
    .D(_01244_),
    .Q(\genblk2.pcpi_div.divisor[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_140_clk),
    .D(_01245_),
    .Q(\genblk2.pcpi_div.divisor[32] ));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_140_clk),
    .D(_01246_),
    .Q(\genblk2.pcpi_div.divisor[33] ));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_140_clk),
    .D(_01247_),
    .Q(\genblk2.pcpi_div.divisor[34] ));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.CLK(clknet_leaf_140_clk),
    .D(_01248_),
    .Q(\genblk2.pcpi_div.divisor[35] ));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_143_clk),
    .D(_01249_),
    .Q(\genblk2.pcpi_div.divisor[36] ));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_143_clk),
    .D(_01250_),
    .Q(\genblk2.pcpi_div.divisor[37] ));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.CLK(clknet_leaf_143_clk),
    .D(_01251_),
    .Q(\genblk2.pcpi_div.divisor[38] ));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.CLK(clknet_leaf_143_clk),
    .D(_01252_),
    .Q(\genblk2.pcpi_div.divisor[39] ));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_143_clk),
    .D(_01253_),
    .Q(\genblk2.pcpi_div.divisor[40] ));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_143_clk),
    .D(_01254_),
    .Q(\genblk2.pcpi_div.divisor[41] ));
 sky130_fd_sc_hd__dfxtp_1 _14903_ (.CLK(clknet_leaf_143_clk),
    .D(_01255_),
    .Q(\genblk2.pcpi_div.divisor[42] ));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.CLK(clknet_leaf_144_clk),
    .D(_01256_),
    .Q(\genblk2.pcpi_div.divisor[43] ));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.CLK(clknet_leaf_142_clk),
    .D(_01257_),
    .Q(\genblk2.pcpi_div.divisor[44] ));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.CLK(clknet_leaf_121_clk),
    .D(_01258_),
    .Q(\genblk2.pcpi_div.divisor[45] ));
 sky130_fd_sc_hd__dfxtp_1 _14907_ (.CLK(clknet_leaf_142_clk),
    .D(_01259_),
    .Q(\genblk2.pcpi_div.divisor[46] ));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.CLK(clknet_leaf_142_clk),
    .D(_01260_),
    .Q(\genblk2.pcpi_div.divisor[47] ));
 sky130_fd_sc_hd__dfxtp_1 _14909_ (.CLK(clknet_leaf_121_clk),
    .D(_01261_),
    .Q(\genblk2.pcpi_div.divisor[48] ));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.CLK(clknet_leaf_121_clk),
    .D(_01262_),
    .Q(\genblk2.pcpi_div.divisor[49] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_122_clk),
    .D(_01263_),
    .Q(\genblk2.pcpi_div.divisor[50] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_121_clk),
    .D(_01264_),
    .Q(\genblk2.pcpi_div.divisor[51] ));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.CLK(clknet_leaf_124_clk),
    .D(_01265_),
    .Q(\genblk2.pcpi_div.divisor[52] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_124_clk),
    .D(_01266_),
    .Q(\genblk2.pcpi_div.divisor[53] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_125_clk),
    .D(_01267_),
    .Q(\genblk2.pcpi_div.divisor[54] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_111_clk),
    .D(_01268_),
    .Q(\genblk2.pcpi_div.divisor[55] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_111_clk),
    .D(_01269_),
    .Q(\genblk2.pcpi_div.divisor[56] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_111_clk),
    .D(_01270_),
    .Q(\genblk2.pcpi_div.divisor[57] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_113_clk),
    .D(_01271_),
    .Q(\genblk2.pcpi_div.divisor[58] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_109_clk),
    .D(_01272_),
    .Q(\genblk2.pcpi_div.divisor[59] ));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.CLK(clknet_leaf_109_clk),
    .D(_01273_),
    .Q(\genblk2.pcpi_div.divisor[60] ));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.CLK(clknet_leaf_108_clk),
    .D(_01274_),
    .Q(\genblk2.pcpi_div.divisor[61] ));
 sky130_fd_sc_hd__dfxtp_1 _14923_ (.CLK(clknet_leaf_30_clk),
    .D(_01275_),
    .Q(\cpuregs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.CLK(clknet_leaf_48_clk),
    .D(_01276_),
    .Q(\cpuregs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.CLK(clknet_leaf_31_clk),
    .D(_01277_),
    .Q(\cpuregs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.CLK(clknet_leaf_17_clk),
    .D(_01278_),
    .Q(\cpuregs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14927_ (.CLK(clknet_leaf_23_clk),
    .D(_01279_),
    .Q(\cpuregs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14928_ (.CLK(clknet_leaf_23_clk),
    .D(_01280_),
    .Q(\cpuregs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14929_ (.CLK(clknet_leaf_179_clk),
    .D(_01281_),
    .Q(\cpuregs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14930_ (.CLK(clknet_leaf_19_clk),
    .D(_01282_),
    .Q(\cpuregs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.CLK(clknet_leaf_180_clk),
    .D(_01283_),
    .Q(\cpuregs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.CLK(clknet_leaf_182_clk),
    .D(_01284_),
    .Q(\cpuregs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.CLK(clknet_leaf_181_clk),
    .D(_01285_),
    .Q(\cpuregs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.CLK(clknet_leaf_20_clk),
    .D(_01286_),
    .Q(\cpuregs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.CLK(clknet_leaf_6_clk),
    .D(_01287_),
    .Q(\cpuregs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.CLK(clknet_leaf_5_clk),
    .D(_01288_),
    .Q(\cpuregs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.CLK(clknet_leaf_19_clk),
    .D(_01289_),
    .Q(\cpuregs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.CLK(clknet_leaf_7_clk),
    .D(_01290_),
    .Q(\cpuregs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.CLK(clknet_leaf_18_clk),
    .D(_01291_),
    .Q(\cpuregs[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.CLK(clknet_leaf_6_clk),
    .D(_01292_),
    .Q(\cpuregs[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14941_ (.CLK(clknet_leaf_8_clk),
    .D(_01293_),
    .Q(\cpuregs[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14942_ (.CLK(clknet_leaf_38_clk),
    .D(_01294_),
    .Q(\cpuregs[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.CLK(clknet_leaf_15_clk),
    .D(_01295_),
    .Q(\cpuregs[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14944_ (.CLK(clknet_leaf_38_clk),
    .D(_01296_),
    .Q(\cpuregs[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.CLK(clknet_leaf_36_clk),
    .D(_01297_),
    .Q(\cpuregs[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.CLK(clknet_leaf_17_clk),
    .D(_01298_),
    .Q(\cpuregs[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14947_ (.CLK(clknet_leaf_35_clk),
    .D(_01299_),
    .Q(\cpuregs[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.CLK(clknet_leaf_72_clk),
    .D(_01300_),
    .Q(\cpuregs[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.CLK(clknet_leaf_33_clk),
    .D(_01301_),
    .Q(\cpuregs[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14950_ (.CLK(clknet_leaf_34_clk),
    .D(_01302_),
    .Q(\cpuregs[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.CLK(clknet_leaf_47_clk),
    .D(_01303_),
    .Q(\cpuregs[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_72_clk),
    .D(_01304_),
    .Q(\cpuregs[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.CLK(clknet_leaf_48_clk),
    .D(_01305_),
    .Q(\cpuregs[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.CLK(clknet_leaf_34_clk),
    .D(_01306_),
    .Q(\cpuregs[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.CLK(clknet_leaf_120_clk),
    .D(_01307_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _14956_ (.CLK(clknet_leaf_120_clk),
    .D(_01308_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14957_ (.CLK(clknet_leaf_121_clk),
    .D(_01309_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.CLK(clknet_leaf_144_clk),
    .D(net2951),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.CLK(clknet_leaf_144_clk),
    .D(_01311_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _14960_ (.CLK(clknet_leaf_144_clk),
    .D(_01312_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _14961_ (.CLK(clknet_leaf_145_clk),
    .D(_01313_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _14962_ (.CLK(clknet_leaf_147_clk),
    .D(_01314_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _14963_ (.CLK(clknet_leaf_147_clk),
    .D(_01315_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _14964_ (.CLK(clknet_leaf_147_clk),
    .D(_01316_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _14965_ (.CLK(clknet_leaf_149_clk),
    .D(_01317_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _14966_ (.CLK(clknet_leaf_149_clk),
    .D(_01318_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _14967_ (.CLK(clknet_leaf_151_clk),
    .D(_01319_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _14968_ (.CLK(clknet_leaf_151_clk),
    .D(_01320_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _14969_ (.CLK(clknet_leaf_150_clk),
    .D(_01321_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _14970_ (.CLK(clknet_leaf_146_clk),
    .D(_01322_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _14971_ (.CLK(clknet_leaf_143_clk),
    .D(_01323_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _14972_ (.CLK(clknet_leaf_143_clk),
    .D(_01324_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.CLK(clknet_leaf_118_clk),
    .D(_01325_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.CLK(clknet_leaf_118_clk),
    .D(_01326_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.CLK(clknet_leaf_116_clk),
    .D(_01327_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _14976_ (.CLK(clknet_leaf_116_clk),
    .D(_01328_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _14977_ (.CLK(clknet_leaf_116_clk),
    .D(_01329_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.CLK(clknet_leaf_112_clk),
    .D(_01330_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _14979_ (.CLK(clknet_leaf_112_clk),
    .D(_01331_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _14980_ (.CLK(clknet_leaf_108_clk),
    .D(_01332_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _14981_ (.CLK(clknet_leaf_107_clk),
    .D(_01333_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _14982_ (.CLK(clknet_leaf_108_clk),
    .D(_01334_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _14983_ (.CLK(clknet_leaf_108_clk),
    .D(_01335_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _14984_ (.CLK(clknet_leaf_108_clk),
    .D(_01336_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _14985_ (.CLK(clknet_leaf_108_clk),
    .D(_01337_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[32] ));
 sky130_fd_sc_hd__dfxtp_1 _14986_ (.CLK(clknet_leaf_112_clk),
    .D(_01338_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[33] ));
 sky130_fd_sc_hd__dfxtp_1 _14987_ (.CLK(clknet_leaf_116_clk),
    .D(_01339_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[34] ));
 sky130_fd_sc_hd__dfxtp_1 _14988_ (.CLK(clknet_leaf_119_clk),
    .D(_01340_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[35] ));
 sky130_fd_sc_hd__dfxtp_1 _14989_ (.CLK(clknet_leaf_119_clk),
    .D(_01341_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[36] ));
 sky130_fd_sc_hd__dfxtp_1 _14990_ (.CLK(clknet_leaf_119_clk),
    .D(_01342_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[37] ));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.CLK(clknet_leaf_118_clk),
    .D(net2895),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[38] ));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.CLK(clknet_leaf_118_clk),
    .D(_01344_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[39] ));
 sky130_fd_sc_hd__dfxtp_1 _14993_ (.CLK(clknet_leaf_145_clk),
    .D(_01345_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[40] ));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.CLK(clknet_leaf_148_clk),
    .D(_01346_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[41] ));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.CLK(clknet_leaf_148_clk),
    .D(net2943),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[42] ));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.CLK(clknet_leaf_148_clk),
    .D(_01348_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[43] ));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.CLK(clknet_leaf_148_clk),
    .D(_01349_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[44] ));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.CLK(clknet_leaf_149_clk),
    .D(net2827),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[45] ));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.CLK(clknet_leaf_150_clk),
    .D(_01351_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[46] ));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.CLK(clknet_leaf_147_clk),
    .D(_01352_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[47] ));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.CLK(clknet_leaf_147_clk),
    .D(net2916),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[48] ));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.CLK(clknet_leaf_147_clk),
    .D(_01354_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[49] ));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.CLK(clknet_leaf_146_clk),
    .D(net2929),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[50] ));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.CLK(clknet_leaf_145_clk),
    .D(_01356_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[51] ));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.CLK(clknet_leaf_118_clk),
    .D(net2846),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[52] ));
 sky130_fd_sc_hd__dfxtp_1 _15006_ (.CLK(clknet_leaf_117_clk),
    .D(_01358_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[53] ));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.CLK(clknet_leaf_117_clk),
    .D(_01359_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[54] ));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.CLK(clknet_leaf_115_clk),
    .D(_01360_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[55] ));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.CLK(clknet_leaf_115_clk),
    .D(_01361_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[56] ));
 sky130_fd_sc_hd__dfxtp_1 _15010_ (.CLK(clknet_leaf_114_clk),
    .D(_01362_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[57] ));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.CLK(clknet_leaf_114_clk),
    .D(net2901),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[58] ));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.CLK(clknet_leaf_113_clk),
    .D(_01364_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[59] ));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.CLK(clknet_leaf_107_clk),
    .D(net2959),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[60] ));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.CLK(clknet_leaf_107_clk),
    .D(_01366_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[61] ));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.CLK(clknet_leaf_106_clk),
    .D(net2946),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[62] ));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.CLK(clknet_leaf_106_clk),
    .D(net2957),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs2[63] ));
 sky130_fd_sc_hd__dfxtp_1 _15017_ (.CLK(clknet_leaf_106_clk),
    .D(net2528),
    .Q(\genblk1.genblk1.pcpi_mul.rs2[63] ));
 sky130_fd_sc_hd__dfxtp_1 _15018_ (.CLK(clknet_leaf_121_clk),
    .D(_01370_),
    .Q(\genblk1.genblk1.pcpi_mul.rs1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15019_ (.CLK(clknet_leaf_122_clk),
    .D(net2410),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15020_ (.CLK(clknet_leaf_122_clk),
    .D(net1492),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15021_ (.CLK(clknet_leaf_122_clk),
    .D(_01373_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15022_ (.CLK(clknet_leaf_140_clk),
    .D(_01374_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15023_ (.CLK(clknet_leaf_140_clk),
    .D(_01375_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15024_ (.CLK(clknet_leaf_139_clk),
    .D(net1365),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15025_ (.CLK(clknet_leaf_140_clk),
    .D(net1355),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15026_ (.CLK(clknet_leaf_139_clk),
    .D(_01378_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15027_ (.CLK(clknet_leaf_138_clk),
    .D(net1543),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15028_ (.CLK(clknet_leaf_137_clk),
    .D(net1336),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15029_ (.CLK(clknet_leaf_137_clk),
    .D(_01381_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15030_ (.CLK(clknet_leaf_137_clk),
    .D(_01382_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _15031_ (.CLK(clknet_leaf_137_clk),
    .D(_01383_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15032_ (.CLK(clknet_leaf_136_clk),
    .D(net1332),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _15033_ (.CLK(clknet_leaf_136_clk),
    .D(net1327),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _15034_ (.CLK(clknet_leaf_135_clk),
    .D(_01386_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _15035_ (.CLK(clknet_leaf_135_clk),
    .D(_01387_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _15036_ (.CLK(clknet_leaf_135_clk),
    .D(net1338),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _15037_ (.CLK(clknet_leaf_135_clk),
    .D(_01389_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _15038_ (.CLK(clknet_leaf_135_clk),
    .D(_01390_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _15039_ (.CLK(clknet_leaf_129_clk),
    .D(net2106),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _15040_ (.CLK(clknet_leaf_129_clk),
    .D(net1329),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _15041_ (.CLK(clknet_leaf_129_clk),
    .D(_01393_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _15042_ (.CLK(clknet_leaf_124_clk),
    .D(_01394_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _15043_ (.CLK(clknet_leaf_125_clk),
    .D(_01395_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _15044_ (.CLK(clknet_leaf_112_clk),
    .D(_01396_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _15045_ (.CLK(clknet_leaf_112_clk),
    .D(net1579),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _15046_ (.CLK(clknet_leaf_112_clk),
    .D(_01398_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _15047_ (.CLK(clknet_leaf_108_clk),
    .D(_01399_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _15048_ (.CLK(clknet_leaf_108_clk),
    .D(_01400_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _15049_ (.CLK(clknet_leaf_105_clk),
    .D(_01401_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _15050_ (.CLK(clknet_leaf_102_clk),
    .D(net2338),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15051_ (.CLK(clknet_leaf_102_clk),
    .D(_01403_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _15052_ (.CLK(clknet_leaf_102_clk),
    .D(net2502),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _15053_ (.CLK(clknet_leaf_102_clk),
    .D(net2479),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _15054_ (.CLK(clknet_leaf_102_clk),
    .D(net2473),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _15055_ (.CLK(clknet_leaf_102_clk),
    .D(net2433),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _15056_ (.CLK(clknet_leaf_102_clk),
    .D(_01408_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _15057_ (.CLK(clknet_leaf_105_clk),
    .D(net2481),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _15058_ (.CLK(clknet_leaf_105_clk),
    .D(net2290),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _15059_ (.CLK(clknet_leaf_104_clk),
    .D(_01411_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _15060_ (.CLK(clknet_leaf_104_clk),
    .D(_01412_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _15061_ (.CLK(clknet_leaf_105_clk),
    .D(net2505),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _15062_ (.CLK(clknet_leaf_105_clk),
    .D(net2108),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _15063_ (.CLK(clknet_leaf_104_clk),
    .D(_01415_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _15064_ (.CLK(clknet_leaf_104_clk),
    .D(net2518),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _15065_ (.CLK(clknet_leaf_104_clk),
    .D(net2234),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _15066_ (.CLK(clknet_leaf_104_clk),
    .D(_01418_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _15067_ (.CLK(clknet_leaf_104_clk),
    .D(net2470),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _15068_ (.CLK(clknet_leaf_104_clk),
    .D(net2265),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _15069_ (.CLK(clknet_leaf_103_clk),
    .D(_01421_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _15070_ (.CLK(clknet_leaf_103_clk),
    .D(_01422_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _15071_ (.CLK(clknet_leaf_103_clk),
    .D(net2376),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _15072_ (.CLK(clknet_leaf_103_clk),
    .D(_01424_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _15073_ (.CLK(clknet_leaf_103_clk),
    .D(net2237),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _15074_ (.CLK(clknet_leaf_103_clk),
    .D(_01426_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _15075_ (.CLK(clknet_leaf_103_clk),
    .D(_01427_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _15076_ (.CLK(clknet_leaf_103_clk),
    .D(net2368),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _15077_ (.CLK(clknet_leaf_103_clk),
    .D(_01429_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _15078_ (.CLK(clknet_leaf_102_clk),
    .D(_01430_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _15079_ (.CLK(clknet_leaf_102_clk),
    .D(net1962),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _15080_ (.CLK(clknet_leaf_103_clk),
    .D(_01432_),
    .Q(\genblk1.genblk1.pcpi_mul.next_rs1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _15081_ (.CLK(clknet_leaf_105_clk),
    .D(_01433_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15082_ (.CLK(clknet_leaf_37_clk),
    .D(_01434_),
    .Q(\cpuregs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15083_ (.CLK(clknet_leaf_48_clk),
    .D(_01435_),
    .Q(\cpuregs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15084_ (.CLK(clknet_leaf_32_clk),
    .D(_01436_),
    .Q(\cpuregs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15085_ (.CLK(clknet_leaf_17_clk),
    .D(_01437_),
    .Q(\cpuregs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15086_ (.CLK(clknet_leaf_29_clk),
    .D(_01438_),
    .Q(\cpuregs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15087_ (.CLK(clknet_leaf_24_clk),
    .D(_01439_),
    .Q(\cpuregs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15088_ (.CLK(clknet_leaf_179_clk),
    .D(_01440_),
    .Q(\cpuregs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15089_ (.CLK(clknet_leaf_19_clk),
    .D(_01441_),
    .Q(\cpuregs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15090_ (.CLK(clknet_leaf_179_clk),
    .D(_01442_),
    .Q(\cpuregs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15091_ (.CLK(clknet_leaf_182_clk),
    .D(_01443_),
    .Q(\cpuregs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15092_ (.CLK(clknet_leaf_181_clk),
    .D(_01444_),
    .Q(\cpuregs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15093_ (.CLK(clknet_leaf_194_clk),
    .D(_01445_),
    .Q(\cpuregs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15094_ (.CLK(clknet_leaf_4_clk),
    .D(_01446_),
    .Q(\cpuregs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15095_ (.CLK(clknet_leaf_4_clk),
    .D(_01447_),
    .Q(\cpuregs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15096_ (.CLK(clknet_leaf_19_clk),
    .D(_01448_),
    .Q(\cpuregs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15097_ (.CLK(clknet_leaf_6_clk),
    .D(_01449_),
    .Q(\cpuregs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15098_ (.CLK(clknet_leaf_18_clk),
    .D(_01450_),
    .Q(\cpuregs[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15099_ (.CLK(clknet_leaf_6_clk),
    .D(_01451_),
    .Q(\cpuregs[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15100_ (.CLK(clknet_leaf_3_clk),
    .D(_01452_),
    .Q(\cpuregs[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15101_ (.CLK(clknet_leaf_38_clk),
    .D(_01453_),
    .Q(\cpuregs[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15102_ (.CLK(clknet_leaf_15_clk),
    .D(_01454_),
    .Q(\cpuregs[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15103_ (.CLK(clknet_leaf_16_clk),
    .D(_01455_),
    .Q(\cpuregs[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15104_ (.CLK(clknet_leaf_36_clk),
    .D(_01456_),
    .Q(\cpuregs[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15105_ (.CLK(clknet_leaf_22_clk),
    .D(_01457_),
    .Q(\cpuregs[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15106_ (.CLK(clknet_leaf_33_clk),
    .D(_01458_),
    .Q(\cpuregs[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15107_ (.CLK(clknet_leaf_73_clk),
    .D(_01459_),
    .Q(\cpuregs[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15108_ (.CLK(clknet_leaf_33_clk),
    .D(_01460_),
    .Q(\cpuregs[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15109_ (.CLK(clknet_leaf_34_clk),
    .D(_01461_),
    .Q(\cpuregs[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15110_ (.CLK(clknet_leaf_48_clk),
    .D(_01462_),
    .Q(\cpuregs[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15111_ (.CLK(clknet_leaf_72_clk),
    .D(_01463_),
    .Q(\cpuregs[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15112_ (.CLK(clknet_leaf_49_clk),
    .D(_01464_),
    .Q(\cpuregs[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15113_ (.CLK(clknet_leaf_49_clk),
    .D(_01465_),
    .Q(\cpuregs[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15114_ (.CLK(clknet_leaf_39_clk),
    .D(_01466_),
    .Q(\cpuregs[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15115_ (.CLK(clknet_leaf_46_clk),
    .D(_01467_),
    .Q(\cpuregs[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15116_ (.CLK(clknet_leaf_28_clk),
    .D(_01468_),
    .Q(\cpuregs[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15117_ (.CLK(clknet_leaf_21_clk),
    .D(_01469_),
    .Q(\cpuregs[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15118_ (.CLK(clknet_leaf_27_clk),
    .D(_01470_),
    .Q(\cpuregs[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15119_ (.CLK(clknet_leaf_24_clk),
    .D(_01471_),
    .Q(\cpuregs[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15120_ (.CLK(clknet_leaf_184_clk),
    .D(_01472_),
    .Q(\cpuregs[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15121_ (.CLK(clknet_leaf_182_clk),
    .D(_01473_),
    .Q(\cpuregs[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15122_ (.CLK(clknet_leaf_183_clk),
    .D(_01474_),
    .Q(\cpuregs[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15123_ (.CLK(clknet_leaf_184_clk),
    .D(_01475_),
    .Q(\cpuregs[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15124_ (.CLK(clknet_leaf_187_clk),
    .D(_01476_),
    .Q(\cpuregs[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15125_ (.CLK(clknet_leaf_192_clk),
    .D(_01477_),
    .Q(\cpuregs[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15126_ (.CLK(clknet_leaf_3_clk),
    .D(_01478_),
    .Q(\cpuregs[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15127_ (.CLK(clknet_leaf_195_clk),
    .D(_01479_),
    .Q(\cpuregs[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15128_ (.CLK(clknet_leaf_192_clk),
    .D(_01480_),
    .Q(\cpuregs[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15129_ (.CLK(clknet_leaf_0_clk),
    .D(_01481_),
    .Q(\cpuregs[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15130_ (.CLK(clknet_leaf_9_clk),
    .D(_01482_),
    .Q(\cpuregs[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15131_ (.CLK(clknet_leaf_0_clk),
    .D(_01483_),
    .Q(\cpuregs[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15132_ (.CLK(clknet_leaf_1_clk),
    .D(_01484_),
    .Q(\cpuregs[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15133_ (.CLK(clknet_leaf_41_clk),
    .D(_01485_),
    .Q(\cpuregs[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15134_ (.CLK(clknet_leaf_12_clk),
    .D(_01486_),
    .Q(\cpuregs[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15135_ (.CLK(clknet_leaf_13_clk),
    .D(_01487_),
    .Q(\cpuregs[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15136_ (.CLK(clknet_leaf_43_clk),
    .D(_01488_),
    .Q(\cpuregs[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15137_ (.CLK(clknet_leaf_16_clk),
    .D(_01489_),
    .Q(\cpuregs[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15138_ (.CLK(clknet_leaf_31_clk),
    .D(_01490_),
    .Q(\cpuregs[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15139_ (.CLK(clknet_leaf_72_clk),
    .D(_01491_),
    .Q(\cpuregs[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15140_ (.CLK(clknet_leaf_71_clk),
    .D(_01492_),
    .Q(\cpuregs[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15141_ (.CLK(clknet_leaf_49_clk),
    .D(_01493_),
    .Q(\cpuregs[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15142_ (.CLK(clknet_leaf_46_clk),
    .D(_01494_),
    .Q(\cpuregs[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15143_ (.CLK(clknet_leaf_73_clk),
    .D(_01495_),
    .Q(\cpuregs[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15144_ (.CLK(clknet_leaf_53_clk),
    .D(_01496_),
    .Q(\cpuregs[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15145_ (.CLK(clknet_leaf_49_clk),
    .D(_01497_),
    .Q(\cpuregs[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15146_ (.CLK(clknet_leaf_80_clk),
    .D(_06748_),
    .Q(\reg_sh[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15147_ (.CLK(clknet_leaf_80_clk),
    .D(_06749_),
    .Q(\reg_sh[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15148_ (.CLK(clknet_leaf_80_clk),
    .D(_06750_),
    .Q(\reg_sh[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15149_ (.CLK(clknet_leaf_91_clk),
    .D(_01498_),
    .Q(\mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15150_ (.CLK(clknet_leaf_91_clk),
    .D(_01499_),
    .Q(\mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15151_ (.CLK(clknet_leaf_90_clk),
    .D(_01500_),
    .Q(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15152_ (.CLK(clknet_leaf_89_clk),
    .D(_01501_),
    .Q(\mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15153_ (.CLK(clknet_leaf_89_clk),
    .D(_01502_),
    .Q(\mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15154_ (.CLK(clknet_leaf_89_clk),
    .D(_01503_),
    .Q(\mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15155_ (.CLK(clknet_leaf_89_clk),
    .D(_01504_),
    .Q(\mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _15156_ (.CLK(clknet_leaf_65_clk),
    .D(_01505_),
    .Q(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15157_ (.CLK(clknet_leaf_65_clk),
    .D(_01506_),
    .Q(\mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_1 _15158_ (.CLK(clknet_leaf_89_clk),
    .D(_01507_),
    .Q(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_1 _15159_ (.CLK(clknet_leaf_89_clk),
    .D(_01508_),
    .Q(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_1 _15160_ (.CLK(clknet_leaf_89_clk),
    .D(_01509_),
    .Q(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_4 _15161_ (.CLK(clknet_leaf_65_clk),
    .D(_01510_),
    .Q(\mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_4 _15162_ (.CLK(clknet_leaf_65_clk),
    .D(_01511_),
    .Q(\mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_4 _15163_ (.CLK(clknet_leaf_65_clk),
    .D(_01512_),
    .Q(\mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _15164_ (.CLK(clknet_leaf_64_clk),
    .D(_01513_),
    .Q(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _15165_ (.CLK(clknet_leaf_65_clk),
    .D(_01514_),
    .Q(\mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _15166_ (.CLK(clknet_leaf_65_clk),
    .D(_01515_),
    .Q(\mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _15167_ (.CLK(clknet_leaf_64_clk),
    .D(_01516_),
    .Q(\mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _15168_ (.CLK(clknet_leaf_65_clk),
    .D(_01517_),
    .Q(\mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _15169_ (.CLK(clknet_leaf_90_clk),
    .D(_01518_),
    .Q(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _15170_ (.CLK(clknet_leaf_65_clk),
    .D(_01519_),
    .Q(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _15171_ (.CLK(clknet_leaf_66_clk),
    .D(_01520_),
    .Q(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _15172_ (.CLK(clknet_leaf_90_clk),
    .D(_01521_),
    .Q(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _15173_ (.CLK(clknet_leaf_91_clk),
    .D(_01522_),
    .Q(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _15174_ (.CLK(clknet_leaf_90_clk),
    .D(_01523_),
    .Q(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 _15175_ (.CLK(clknet_leaf_90_clk),
    .D(_01524_),
    .Q(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_2 _15176_ (.CLK(clknet_leaf_90_clk),
    .D(_01525_),
    .Q(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _15177_ (.CLK(clknet_leaf_89_clk),
    .D(_01526_),
    .Q(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _15178_ (.CLK(clknet_leaf_89_clk),
    .D(_01527_),
    .Q(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_4 _15179_ (.CLK(clknet_leaf_91_clk),
    .D(_01528_),
    .Q(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _15180_ (.CLK(clknet_leaf_65_clk),
    .D(_01529_),
    .Q(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _15181_ (.CLK(clknet_leaf_37_clk),
    .D(_01530_),
    .Q(\cpuregs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15182_ (.CLK(clknet_leaf_35_clk),
    .D(_01531_),
    .Q(\cpuregs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15183_ (.CLK(clknet_leaf_32_clk),
    .D(_01532_),
    .Q(\cpuregs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15184_ (.CLK(clknet_leaf_17_clk),
    .D(_01533_),
    .Q(\cpuregs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15185_ (.CLK(clknet_leaf_29_clk),
    .D(_01534_),
    .Q(\cpuregs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15186_ (.CLK(clknet_leaf_24_clk),
    .D(_01535_),
    .Q(\cpuregs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15187_ (.CLK(clknet_leaf_179_clk),
    .D(_01536_),
    .Q(\cpuregs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15188_ (.CLK(clknet_leaf_19_clk),
    .D(_01537_),
    .Q(\cpuregs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15189_ (.CLK(clknet_leaf_179_clk),
    .D(_01538_),
    .Q(\cpuregs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15190_ (.CLK(clknet_leaf_184_clk),
    .D(_01539_),
    .Q(\cpuregs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15191_ (.CLK(clknet_leaf_181_clk),
    .D(_01540_),
    .Q(\cpuregs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15192_ (.CLK(clknet_leaf_5_clk),
    .D(_01541_),
    .Q(\cpuregs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15193_ (.CLK(clknet_leaf_4_clk),
    .D(_01542_),
    .Q(\cpuregs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15194_ (.CLK(clknet_leaf_5_clk),
    .D(_01543_),
    .Q(\cpuregs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15195_ (.CLK(clknet_leaf_19_clk),
    .D(_01544_),
    .Q(\cpuregs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15196_ (.CLK(clknet_leaf_6_clk),
    .D(_01545_),
    .Q(\cpuregs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15197_ (.CLK(clknet_leaf_18_clk),
    .D(_01546_),
    .Q(\cpuregs[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15198_ (.CLK(clknet_leaf_6_clk),
    .D(_01547_),
    .Q(\cpuregs[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15199_ (.CLK(clknet_leaf_6_clk),
    .D(_01548_),
    .Q(\cpuregs[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15200_ (.CLK(clknet_leaf_38_clk),
    .D(_01549_),
    .Q(\cpuregs[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15201_ (.CLK(clknet_leaf_15_clk),
    .D(_01550_),
    .Q(\cpuregs[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15202_ (.CLK(clknet_leaf_38_clk),
    .D(_01551_),
    .Q(\cpuregs[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15203_ (.CLK(clknet_leaf_36_clk),
    .D(_01552_),
    .Q(\cpuregs[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15204_ (.CLK(clknet_leaf_22_clk),
    .D(_01553_),
    .Q(\cpuregs[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15205_ (.CLK(clknet_leaf_33_clk),
    .D(_01554_),
    .Q(\cpuregs[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15206_ (.CLK(clknet_leaf_72_clk),
    .D(_01555_),
    .Q(\cpuregs[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15207_ (.CLK(clknet_leaf_33_clk),
    .D(_01556_),
    .Q(\cpuregs[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15208_ (.CLK(clknet_leaf_34_clk),
    .D(_01557_),
    .Q(\cpuregs[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15209_ (.CLK(clknet_leaf_48_clk),
    .D(_01558_),
    .Q(\cpuregs[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15210_ (.CLK(clknet_leaf_72_clk),
    .D(_01559_),
    .Q(\cpuregs[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15211_ (.CLK(clknet_leaf_50_clk),
    .D(_01560_),
    .Q(\cpuregs[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15212_ (.CLK(clknet_leaf_49_clk),
    .D(_01561_),
    .Q(\cpuregs[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15213_ (.CLK(clknet_leaf_98_clk),
    .D(_01562_),
    .Q(\genblk1.genblk1.pcpi_mul.instr_mulhsu ));
 sky130_fd_sc_hd__dfxtp_1 _15214_ (.CLK(clknet_leaf_99_clk),
    .D(_01563_),
    .Q(\genblk1.genblk1.pcpi_mul.instr_mulh ));
 sky130_fd_sc_hd__dfxtp_1 _15215_ (.CLK(clknet_leaf_88_clk),
    .D(_00004_),
    .Q(\cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15216_ (.CLK(clknet_leaf_87_clk),
    .D(_00005_),
    .Q(\cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15217_ (.CLK(clknet_leaf_86_clk),
    .D(_00006_),
    .Q(\cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _15218_ (.CLK(clknet_leaf_88_clk),
    .D(_00007_),
    .Q(\cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _15219_ (.CLK(clknet_leaf_87_clk),
    .D(_00008_),
    .Q(\cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_1 _15220_ (.CLK(clknet_leaf_88_clk),
    .D(_00009_),
    .Q(\cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_1 _15221_ (.CLK(clknet_leaf_85_clk),
    .D(_00010_),
    .Q(\cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_1 _15222_ (.CLK(clknet_leaf_87_clk),
    .D(_00011_),
    .Q(\cpu_state[7] ));
 sky130_fd_sc_hd__dfxtp_1 _15223_ (.CLK(clknet_leaf_79_clk),
    .D(_01564_),
    .Q(\reg_sh[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15224_ (.CLK(clknet_leaf_79_clk),
    .D(_01565_),
    .Q(\reg_sh[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15225_ (.CLK(clknet_leaf_37_clk),
    .D(_01566_),
    .Q(\cpuregs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15226_ (.CLK(clknet_leaf_47_clk),
    .D(_01567_),
    .Q(\cpuregs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15227_ (.CLK(clknet_leaf_32_clk),
    .D(_01568_),
    .Q(\cpuregs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15228_ (.CLK(clknet_leaf_22_clk),
    .D(_01569_),
    .Q(\cpuregs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15229_ (.CLK(clknet_leaf_23_clk),
    .D(_01570_),
    .Q(\cpuregs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15230_ (.CLK(clknet_leaf_22_clk),
    .D(_01571_),
    .Q(\cpuregs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15231_ (.CLK(clknet_leaf_180_clk),
    .D(_01572_),
    .Q(\cpuregs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15232_ (.CLK(clknet_leaf_20_clk),
    .D(_01573_),
    .Q(\cpuregs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15233_ (.CLK(clknet_leaf_180_clk),
    .D(_01574_),
    .Q(\cpuregs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15234_ (.CLK(clknet_leaf_181_clk),
    .D(_01575_),
    .Q(\cpuregs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15235_ (.CLK(clknet_leaf_20_clk),
    .D(_01576_),
    .Q(\cpuregs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15236_ (.CLK(clknet_leaf_5_clk),
    .D(_01577_),
    .Q(\cpuregs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15237_ (.CLK(clknet_leaf_6_clk),
    .D(_01578_),
    .Q(\cpuregs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15238_ (.CLK(clknet_leaf_5_clk),
    .D(_01579_),
    .Q(\cpuregs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15239_ (.CLK(clknet_leaf_19_clk),
    .D(_01580_),
    .Q(\cpuregs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15240_ (.CLK(clknet_leaf_7_clk),
    .D(_01581_),
    .Q(\cpuregs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15241_ (.CLK(clknet_leaf_18_clk),
    .D(_01582_),
    .Q(\cpuregs[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15242_ (.CLK(clknet_leaf_7_clk),
    .D(_01583_),
    .Q(\cpuregs[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15243_ (.CLK(clknet_leaf_7_clk),
    .D(_01584_),
    .Q(\cpuregs[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15244_ (.CLK(clknet_leaf_41_clk),
    .D(_01585_),
    .Q(\cpuregs[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15245_ (.CLK(clknet_leaf_14_clk),
    .D(_01586_),
    .Q(\cpuregs[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15246_ (.CLK(clknet_leaf_16_clk),
    .D(_01587_),
    .Q(\cpuregs[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15247_ (.CLK(clknet_leaf_40_clk),
    .D(_01588_),
    .Q(\cpuregs[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15248_ (.CLK(clknet_leaf_16_clk),
    .D(_01589_),
    .Q(\cpuregs[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15249_ (.CLK(clknet_leaf_32_clk),
    .D(_01590_),
    .Q(\cpuregs[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15250_ (.CLK(clknet_leaf_32_clk),
    .D(_01591_),
    .Q(\cpuregs[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15251_ (.CLK(clknet_leaf_34_clk),
    .D(_01592_),
    .Q(\cpuregs[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15252_ (.CLK(clknet_leaf_48_clk),
    .D(_01593_),
    .Q(\cpuregs[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15253_ (.CLK(clknet_leaf_47_clk),
    .D(_01594_),
    .Q(\cpuregs[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15254_ (.CLK(clknet_leaf_72_clk),
    .D(_01595_),
    .Q(\cpuregs[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15255_ (.CLK(clknet_leaf_46_clk),
    .D(_01596_),
    .Q(\cpuregs[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15256_ (.CLK(clknet_leaf_49_clk),
    .D(_01597_),
    .Q(\cpuregs[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15257_ (.CLK(clknet_leaf_37_clk),
    .D(_01598_),
    .Q(\cpuregs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15258_ (.CLK(clknet_leaf_32_clk),
    .D(_01599_),
    .Q(\cpuregs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15259_ (.CLK(clknet_leaf_20_clk),
    .D(_01600_),
    .Q(\cpuregs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15260_ (.CLK(clknet_leaf_11_clk),
    .D(_01601_),
    .Q(\cpuregs[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15261_ (.CLK(clknet_leaf_7_clk),
    .D(_01602_),
    .Q(\cpuregs[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15262_ (.CLK(clknet_leaf_41_clk),
    .D(_01603_),
    .Q(\cpuregs[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15263_ (.CLK(clknet_leaf_33_clk),
    .D(_01604_),
    .Q(\cpuregs[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15264_ (.CLK(clknet_leaf_52_clk),
    .D(_01605_),
    .Q(\cpuregs[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15265_ (.CLK(clknet_leaf_57_clk),
    .D(_01606_),
    .Q(\cpuregs[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15266_ (.CLK(clknet_leaf_38_clk),
    .D(_01607_),
    .Q(\cpuregs[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15267_ (.CLK(clknet_leaf_47_clk),
    .D(_01608_),
    .Q(\cpuregs[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15268_ (.CLK(clknet_leaf_73_clk),
    .D(_01609_),
    .Q(\cpuregs[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15269_ (.CLK(clknet_leaf_176_clk),
    .D(_01610_),
    .Q(\cpuregs[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15270_ (.CLK(clknet_leaf_25_clk),
    .D(_01611_),
    .Q(\cpuregs[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15271_ (.CLK(clknet_leaf_25_clk),
    .D(_01612_),
    .Q(\cpuregs[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15272_ (.CLK(clknet_leaf_178_clk),
    .D(_01613_),
    .Q(\cpuregs[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15273_ (.CLK(clknet_leaf_188_clk),
    .D(_01614_),
    .Q(\cpuregs[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15274_ (.CLK(clknet_leaf_185_clk),
    .D(_01615_),
    .Q(\cpuregs[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15275_ (.CLK(clknet_leaf_185_clk),
    .D(_01616_),
    .Q(\cpuregs[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15276_ (.CLK(clknet_leaf_185_clk),
    .D(_01617_),
    .Q(\cpuregs[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15277_ (.CLK(clknet_leaf_191_clk),
    .D(_01618_),
    .Q(\cpuregs[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15278_ (.CLK(clknet_leaf_198_clk),
    .D(_01619_),
    .Q(\cpuregs[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15279_ (.CLK(clknet_leaf_196_clk),
    .D(_01620_),
    .Q(\cpuregs[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15280_ (.CLK(clknet_leaf_191_clk),
    .D(_01621_),
    .Q(\cpuregs[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15281_ (.CLK(clknet_leaf_199_clk),
    .D(_01622_),
    .Q(\cpuregs[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15282_ (.CLK(clknet_leaf_7_clk),
    .D(_01623_),
    .Q(\cpuregs[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15283_ (.CLK(clknet_leaf_2_clk),
    .D(_01624_),
    .Q(\cpuregs[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15284_ (.CLK(clknet_leaf_2_clk),
    .D(_01625_),
    .Q(\cpuregs[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15285_ (.CLK(clknet_leaf_41_clk),
    .D(_01626_),
    .Q(\cpuregs[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15286_ (.CLK(clknet_leaf_15_clk),
    .D(_01627_),
    .Q(\cpuregs[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15287_ (.CLK(clknet_leaf_14_clk),
    .D(_01628_),
    .Q(\cpuregs[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15288_ (.CLK(clknet_leaf_40_clk),
    .D(_01629_),
    .Q(\cpuregs[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15289_ (.CLK(clknet_leaf_30_clk),
    .D(_01630_),
    .Q(\cpuregs[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15290_ (.CLK(clknet_leaf_30_clk),
    .D(_01631_),
    .Q(\cpuregs[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15291_ (.CLK(clknet_leaf_60_clk),
    .D(_01632_),
    .Q(\cpuregs[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15292_ (.CLK(clknet_4_10_0_clk),
    .D(_01633_),
    .Q(\cpuregs[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15293_ (.CLK(clknet_leaf_56_clk),
    .D(_01634_),
    .Q(\cpuregs[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15294_ (.CLK(clknet_leaf_51_clk),
    .D(_01635_),
    .Q(\cpuregs[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15295_ (.CLK(clknet_leaf_66_clk),
    .D(_01636_),
    .Q(\cpuregs[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15296_ (.CLK(clknet_leaf_54_clk),
    .D(_01637_),
    .Q(\cpuregs[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15297_ (.CLK(clknet_leaf_56_clk),
    .D(_01638_),
    .Q(\cpuregs[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15298_ (.CLK(clknet_leaf_99_clk),
    .D(_01639_),
    .Q(\genblk1.genblk1.pcpi_mul.instr_mul ));
 sky130_fd_sc_hd__dfxtp_1 _15299_ (.CLK(clknet_leaf_105_clk),
    .D(_01640_),
    .Q(\genblk1.genblk1.pcpi_mul.mul_finish ));
 sky130_fd_sc_hd__dfxtp_1 _15300_ (.CLK(clknet_leaf_102_clk),
    .D(net1315),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_wait_q ));
 sky130_fd_sc_hd__dfxtp_1 _15301_ (.CLK(clknet_leaf_36_clk),
    .D(_01641_),
    .Q(\cpuregs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15302_ (.CLK(clknet_leaf_44_clk),
    .D(_01642_),
    .Q(\cpuregs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15303_ (.CLK(clknet_leaf_31_clk),
    .D(_01643_),
    .Q(\cpuregs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15304_ (.CLK(clknet_leaf_17_clk),
    .D(_01644_),
    .Q(\cpuregs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15305_ (.CLK(clknet_leaf_30_clk),
    .D(_01645_),
    .Q(\cpuregs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15306_ (.CLK(clknet_leaf_21_clk),
    .D(_01646_),
    .Q(\cpuregs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15307_ (.CLK(clknet_leaf_21_clk),
    .D(_01647_),
    .Q(\cpuregs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15308_ (.CLK(clknet_leaf_19_clk),
    .D(_01648_),
    .Q(\cpuregs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15309_ (.CLK(clknet_leaf_182_clk),
    .D(_01649_),
    .Q(\cpuregs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15310_ (.CLK(clknet_leaf_181_clk),
    .D(_01650_),
    .Q(\cpuregs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15311_ (.CLK(clknet_leaf_193_clk),
    .D(_01651_),
    .Q(\cpuregs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15312_ (.CLK(clknet_leaf_194_clk),
    .D(_01652_),
    .Q(\cpuregs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15313_ (.CLK(clknet_leaf_3_clk),
    .D(_01653_),
    .Q(\cpuregs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15314_ (.CLK(clknet_leaf_4_clk),
    .D(_01654_),
    .Q(\cpuregs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15315_ (.CLK(clknet_leaf_4_clk),
    .D(_01655_),
    .Q(\cpuregs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15316_ (.CLK(clknet_leaf_8_clk),
    .D(_01656_),
    .Q(\cpuregs[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15317_ (.CLK(clknet_leaf_11_clk),
    .D(_01657_),
    .Q(\cpuregs[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15318_ (.CLK(clknet_leaf_9_clk),
    .D(_01658_),
    .Q(\cpuregs[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15319_ (.CLK(clknet_leaf_7_clk),
    .D(_01659_),
    .Q(\cpuregs[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15320_ (.CLK(clknet_leaf_40_clk),
    .D(_01660_),
    .Q(\cpuregs[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15321_ (.CLK(clknet_leaf_14_clk),
    .D(_01661_),
    .Q(\cpuregs[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15322_ (.CLK(clknet_leaf_15_clk),
    .D(_01662_),
    .Q(\cpuregs[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15323_ (.CLK(clknet_leaf_43_clk),
    .D(_01663_),
    .Q(\cpuregs[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15324_ (.CLK(clknet_leaf_16_clk),
    .D(_01664_),
    .Q(\cpuregs[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15325_ (.CLK(clknet_leaf_35_clk),
    .D(_01665_),
    .Q(\cpuregs[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15326_ (.CLK(clknet_leaf_58_clk),
    .D(_01666_),
    .Q(\cpuregs[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15327_ (.CLK(clknet_leaf_57_clk),
    .D(_01667_),
    .Q(\cpuregs[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15328_ (.CLK(clknet_leaf_50_clk),
    .D(_01668_),
    .Q(\cpuregs[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15329_ (.CLK(clknet_leaf_52_clk),
    .D(_01669_),
    .Q(\cpuregs[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15330_ (.CLK(clknet_leaf_70_clk),
    .D(_01670_),
    .Q(\cpuregs[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15331_ (.CLK(clknet_leaf_54_clk),
    .D(_01671_),
    .Q(\cpuregs[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15332_ (.CLK(clknet_leaf_57_clk),
    .D(_01672_),
    .Q(\cpuregs[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15333_ (.CLK(clknet_leaf_159_clk),
    .D(_01673_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _15334_ (.CLK(clknet_leaf_156_clk),
    .D(_01674_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _15335_ (.CLK(clknet_leaf_145_clk),
    .D(_01675_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _15336_ (.CLK(clknet_leaf_149_clk),
    .D(_01676_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _15337_ (.CLK(clknet_leaf_166_clk),
    .D(_01677_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _15338_ (.CLK(clknet_leaf_166_clk),
    .D(_01678_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _15339_ (.CLK(clknet_leaf_166_clk),
    .D(_01679_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _15340_ (.CLK(clknet_leaf_166_clk),
    .D(_01680_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _15341_ (.CLK(clknet_leaf_166_clk),
    .D(_01681_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _15342_ (.CLK(clknet_leaf_189_clk),
    .D(_01682_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _15343_ (.CLK(clknet_leaf_189_clk),
    .D(_01683_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _15344_ (.CLK(clknet_leaf_189_clk),
    .D(_01684_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _15345_ (.CLK(clknet_leaf_189_clk),
    .D(_01685_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _15346_ (.CLK(clknet_leaf_12_clk),
    .D(_01686_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _15347_ (.CLK(clknet_leaf_12_clk),
    .D(_01687_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _15348_ (.CLK(clknet_leaf_13_clk),
    .D(_01688_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _15349_ (.CLK(clknet_leaf_42_clk),
    .D(_01689_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _15350_ (.CLK(clknet_leaf_42_clk),
    .D(_01690_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _15351_ (.CLK(clknet_leaf_43_clk),
    .D(_01691_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _15352_ (.CLK(clknet_leaf_62_clk),
    .D(_01692_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _15353_ (.CLK(clknet_leaf_55_clk),
    .D(_01693_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _15354_ (.CLK(clknet_leaf_62_clk),
    .D(_01694_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _15355_ (.CLK(clknet_leaf_93_clk),
    .D(_01695_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _15356_ (.CLK(clknet_leaf_93_clk),
    .D(_01696_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _15357_ (.CLK(clknet_leaf_55_clk),
    .D(_01697_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _15358_ (.CLK(clknet_leaf_55_clk),
    .D(_01698_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _15359_ (.CLK(clknet_leaf_55_clk),
    .D(_01699_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _15360_ (.CLK(clknet_leaf_64_clk),
    .D(_01700_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _15361_ (.CLK(clknet_leaf_62_clk),
    .D(_01701_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _15362_ (.CLK(clknet_leaf_64_clk),
    .D(_01702_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _15363_ (.CLK(clknet_leaf_102_clk),
    .D(\genblk1.genblk1.pcpi_mul.instr_any_mul ),
    .Q(\genblk1.genblk1.pcpi_mul.pcpi_wait ));
 sky130_fd_sc_hd__dfxtp_1 _15364_ (.CLK(clknet_leaf_38_clk),
    .D(_01703_),
    .Q(\cpuregs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15365_ (.CLK(clknet_leaf_45_clk),
    .D(_01704_),
    .Q(\cpuregs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15366_ (.CLK(clknet_leaf_31_clk),
    .D(_01705_),
    .Q(\cpuregs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15367_ (.CLK(clknet_leaf_17_clk),
    .D(_01706_),
    .Q(\cpuregs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15368_ (.CLK(clknet_leaf_30_clk),
    .D(_01707_),
    .Q(\cpuregs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15369_ (.CLK(clknet_leaf_22_clk),
    .D(_01708_),
    .Q(\cpuregs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15370_ (.CLK(clknet_leaf_180_clk),
    .D(_01709_),
    .Q(\cpuregs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15371_ (.CLK(clknet_leaf_20_clk),
    .D(_01710_),
    .Q(\cpuregs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15372_ (.CLK(clknet_leaf_182_clk),
    .D(_01711_),
    .Q(\cpuregs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15373_ (.CLK(clknet_leaf_181_clk),
    .D(_01712_),
    .Q(\cpuregs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15374_ (.CLK(clknet_leaf_193_clk),
    .D(_01713_),
    .Q(\cpuregs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15375_ (.CLK(clknet_leaf_194_clk),
    .D(_01714_),
    .Q(\cpuregs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15376_ (.CLK(clknet_leaf_2_clk),
    .D(_01715_),
    .Q(\cpuregs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15377_ (.CLK(clknet_leaf_3_clk),
    .D(_01716_),
    .Q(\cpuregs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15378_ (.CLK(clknet_leaf_4_clk),
    .D(_01717_),
    .Q(\cpuregs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15379_ (.CLK(clknet_leaf_1_clk),
    .D(_01718_),
    .Q(\cpuregs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15380_ (.CLK(clknet_leaf_10_clk),
    .D(_01719_),
    .Q(\cpuregs[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15381_ (.CLK(clknet_leaf_9_clk),
    .D(_01720_),
    .Q(\cpuregs[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15382_ (.CLK(clknet_leaf_8_clk),
    .D(_01721_),
    .Q(\cpuregs[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15383_ (.CLK(clknet_leaf_41_clk),
    .D(_01722_),
    .Q(\cpuregs[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15384_ (.CLK(clknet_leaf_12_clk),
    .D(_01723_),
    .Q(\cpuregs[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15385_ (.CLK(clknet_leaf_15_clk),
    .D(_01724_),
    .Q(\cpuregs[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15386_ (.CLK(clknet_leaf_43_clk),
    .D(_01725_),
    .Q(\cpuregs[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15387_ (.CLK(clknet_leaf_16_clk),
    .D(_01726_),
    .Q(\cpuregs[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15388_ (.CLK(clknet_leaf_36_clk),
    .D(_01727_),
    .Q(\cpuregs[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15389_ (.CLK(clknet_leaf_57_clk),
    .D(_01728_),
    .Q(\cpuregs[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15390_ (.CLK(clknet_leaf_57_clk),
    .D(_01729_),
    .Q(\cpuregs[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15391_ (.CLK(clknet_leaf_50_clk),
    .D(_01730_),
    .Q(\cpuregs[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15392_ (.CLK(clknet_leaf_52_clk),
    .D(_01731_),
    .Q(\cpuregs[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15393_ (.CLK(clknet_leaf_71_clk),
    .D(_01732_),
    .Q(\cpuregs[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15394_ (.CLK(clknet_leaf_53_clk),
    .D(_01733_),
    .Q(\cpuregs[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15395_ (.CLK(clknet_leaf_49_clk),
    .D(_01734_),
    .Q(\cpuregs[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15396_ (.CLK(clknet_leaf_37_clk),
    .D(_01735_),
    .Q(\cpuregs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15397_ (.CLK(clknet_leaf_45_clk),
    .D(_01736_),
    .Q(\cpuregs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15398_ (.CLK(clknet_leaf_31_clk),
    .D(_01737_),
    .Q(\cpuregs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15399_ (.CLK(clknet_leaf_17_clk),
    .D(_01738_),
    .Q(\cpuregs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15400_ (.CLK(clknet_leaf_30_clk),
    .D(_01739_),
    .Q(\cpuregs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15401_ (.CLK(clknet_leaf_24_clk),
    .D(_01740_),
    .Q(\cpuregs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15402_ (.CLK(clknet_leaf_179_clk),
    .D(_01741_),
    .Q(\cpuregs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15403_ (.CLK(clknet_leaf_20_clk),
    .D(_01742_),
    .Q(\cpuregs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15404_ (.CLK(clknet_leaf_182_clk),
    .D(_01743_),
    .Q(\cpuregs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15405_ (.CLK(clknet_leaf_181_clk),
    .D(_01744_),
    .Q(\cpuregs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15406_ (.CLK(clknet_leaf_193_clk),
    .D(_01745_),
    .Q(\cpuregs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15407_ (.CLK(clknet_leaf_194_clk),
    .D(_01746_),
    .Q(\cpuregs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15408_ (.CLK(clknet_leaf_3_clk),
    .D(_01747_),
    .Q(\cpuregs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15409_ (.CLK(clknet_leaf_4_clk),
    .D(_01748_),
    .Q(\cpuregs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15410_ (.CLK(clknet_leaf_4_clk),
    .D(_01749_),
    .Q(\cpuregs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15411_ (.CLK(clknet_leaf_9_clk),
    .D(_01750_),
    .Q(\cpuregs[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15412_ (.CLK(clknet_leaf_10_clk),
    .D(_01751_),
    .Q(\cpuregs[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15413_ (.CLK(clknet_leaf_9_clk),
    .D(_01752_),
    .Q(\cpuregs[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15414_ (.CLK(clknet_leaf_9_clk),
    .D(_01753_),
    .Q(\cpuregs[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15415_ (.CLK(clknet_leaf_41_clk),
    .D(_01754_),
    .Q(\cpuregs[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15416_ (.CLK(clknet_leaf_11_clk),
    .D(_01755_),
    .Q(\cpuregs[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15417_ (.CLK(clknet_leaf_16_clk),
    .D(_01756_),
    .Q(\cpuregs[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15418_ (.CLK(clknet_leaf_43_clk),
    .D(_01757_),
    .Q(\cpuregs[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15419_ (.CLK(clknet_leaf_16_clk),
    .D(_01758_),
    .Q(\cpuregs[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15420_ (.CLK(clknet_leaf_35_clk),
    .D(_01759_),
    .Q(\cpuregs[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15421_ (.CLK(clknet_leaf_57_clk),
    .D(_01760_),
    .Q(\cpuregs[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15422_ (.CLK(clknet_leaf_57_clk),
    .D(_01761_),
    .Q(\cpuregs[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15423_ (.CLK(clknet_leaf_50_clk),
    .D(_01762_),
    .Q(\cpuregs[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15424_ (.CLK(clknet_leaf_52_clk),
    .D(_01763_),
    .Q(\cpuregs[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15425_ (.CLK(clknet_leaf_71_clk),
    .D(_01764_),
    .Q(\cpuregs[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15426_ (.CLK(clknet_leaf_53_clk),
    .D(_01765_),
    .Q(\cpuregs[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15427_ (.CLK(clknet_leaf_57_clk),
    .D(_01766_),
    .Q(\cpuregs[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15428_ (.CLK(clknet_leaf_38_clk),
    .D(_01767_),
    .Q(\cpuregs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15429_ (.CLK(clknet_leaf_45_clk),
    .D(_01768_),
    .Q(\cpuregs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15430_ (.CLK(clknet_leaf_29_clk),
    .D(_01769_),
    .Q(\cpuregs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15431_ (.CLK(clknet_leaf_18_clk),
    .D(_01770_),
    .Q(\cpuregs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15432_ (.CLK(clknet_leaf_29_clk),
    .D(_01771_),
    .Q(\cpuregs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15433_ (.CLK(clknet_leaf_22_clk),
    .D(_01772_),
    .Q(\cpuregs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15434_ (.CLK(clknet_leaf_181_clk),
    .D(_01773_),
    .Q(\cpuregs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15435_ (.CLK(clknet_leaf_20_clk),
    .D(_01774_),
    .Q(\cpuregs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15436_ (.CLK(clknet_leaf_192_clk),
    .D(_01775_),
    .Q(\cpuregs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15437_ (.CLK(clknet_leaf_192_clk),
    .D(_01776_),
    .Q(\cpuregs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15438_ (.CLK(clknet_leaf_193_clk),
    .D(_01777_),
    .Q(\cpuregs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15439_ (.CLK(clknet_leaf_194_clk),
    .D(_01778_),
    .Q(\cpuregs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15440_ (.CLK(clknet_leaf_3_clk),
    .D(_01779_),
    .Q(\cpuregs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15441_ (.CLK(clknet_leaf_195_clk),
    .D(_01780_),
    .Q(\cpuregs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15442_ (.CLK(clknet_leaf_195_clk),
    .D(_01781_),
    .Q(\cpuregs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15443_ (.CLK(clknet_leaf_1_clk),
    .D(_01782_),
    .Q(\cpuregs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15444_ (.CLK(clknet_leaf_10_clk),
    .D(_01783_),
    .Q(\cpuregs[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15445_ (.CLK(clknet_leaf_9_clk),
    .D(_01784_),
    .Q(\cpuregs[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15446_ (.CLK(clknet_leaf_9_clk),
    .D(_01785_),
    .Q(\cpuregs[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15447_ (.CLK(clknet_leaf_41_clk),
    .D(_01786_),
    .Q(\cpuregs[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15448_ (.CLK(clknet_leaf_12_clk),
    .D(_01787_),
    .Q(\cpuregs[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15449_ (.CLK(clknet_leaf_15_clk),
    .D(_01788_),
    .Q(\cpuregs[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15450_ (.CLK(clknet_leaf_42_clk),
    .D(_01789_),
    .Q(\cpuregs[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15451_ (.CLK(clknet_leaf_17_clk),
    .D(_01790_),
    .Q(\cpuregs[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15452_ (.CLK(clknet_leaf_35_clk),
    .D(_01791_),
    .Q(\cpuregs[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15453_ (.CLK(clknet_leaf_59_clk),
    .D(_01792_),
    .Q(\cpuregs[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15454_ (.CLK(clknet_leaf_56_clk),
    .D(_01793_),
    .Q(\cpuregs[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15455_ (.CLK(clknet_leaf_51_clk),
    .D(_01794_),
    .Q(\cpuregs[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15456_ (.CLK(clknet_leaf_53_clk),
    .D(_01795_),
    .Q(\cpuregs[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15457_ (.CLK(clknet_leaf_59_clk),
    .D(_01796_),
    .Q(\cpuregs[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15458_ (.CLK(clknet_leaf_54_clk),
    .D(_01797_),
    .Q(\cpuregs[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15459_ (.CLK(clknet_leaf_56_clk),
    .D(_01798_),
    .Q(\cpuregs[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15460_ (.CLK(clknet_leaf_85_clk),
    .D(_00012_),
    .Q(\mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_1 _15461_ (.CLK(clknet_leaf_85_clk),
    .D(_00013_),
    .Q(\mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_1 _15462_ (.CLK(clknet_leaf_85_clk),
    .D(_00014_),
    .Q(\mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_1 _15463_ (.CLK(clknet_leaf_38_clk),
    .D(_01799_),
    .Q(\cpuregs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15464_ (.CLK(clknet_leaf_45_clk),
    .D(_01800_),
    .Q(\cpuregs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15465_ (.CLK(clknet_leaf_31_clk),
    .D(_01801_),
    .Q(\cpuregs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15466_ (.CLK(clknet_leaf_18_clk),
    .D(_01802_),
    .Q(\cpuregs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15467_ (.CLK(clknet_leaf_29_clk),
    .D(_01803_),
    .Q(\cpuregs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15468_ (.CLK(clknet_leaf_22_clk),
    .D(_01804_),
    .Q(\cpuregs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15469_ (.CLK(clknet_leaf_20_clk),
    .D(_01805_),
    .Q(\cpuregs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15470_ (.CLK(clknet_leaf_20_clk),
    .D(_01806_),
    .Q(\cpuregs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15471_ (.CLK(clknet_leaf_192_clk),
    .D(_01807_),
    .Q(\cpuregs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15472_ (.CLK(clknet_leaf_192_clk),
    .D(_01808_),
    .Q(\cpuregs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15473_ (.CLK(clknet_leaf_192_clk),
    .D(_01809_),
    .Q(\cpuregs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15474_ (.CLK(clknet_leaf_194_clk),
    .D(_01810_),
    .Q(\cpuregs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15475_ (.CLK(clknet_leaf_3_clk),
    .D(_01811_),
    .Q(\cpuregs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15476_ (.CLK(clknet_leaf_195_clk),
    .D(_01812_),
    .Q(\cpuregs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15477_ (.CLK(clknet_leaf_195_clk),
    .D(_01813_),
    .Q(\cpuregs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15478_ (.CLK(clknet_leaf_9_clk),
    .D(_01814_),
    .Q(\cpuregs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15479_ (.CLK(clknet_leaf_10_clk),
    .D(_01815_),
    .Q(\cpuregs[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15480_ (.CLK(clknet_leaf_9_clk),
    .D(_01816_),
    .Q(\cpuregs[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15481_ (.CLK(clknet_leaf_9_clk),
    .D(_01817_),
    .Q(\cpuregs[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15482_ (.CLK(clknet_leaf_42_clk),
    .D(_01818_),
    .Q(\cpuregs[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15483_ (.CLK(clknet_leaf_12_clk),
    .D(_01819_),
    .Q(\cpuregs[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15484_ (.CLK(clknet_leaf_15_clk),
    .D(_01820_),
    .Q(\cpuregs[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15485_ (.CLK(clknet_leaf_42_clk),
    .D(_01821_),
    .Q(\cpuregs[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15486_ (.CLK(clknet_leaf_17_clk),
    .D(_01822_),
    .Q(\cpuregs[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15487_ (.CLK(clknet_leaf_35_clk),
    .D(_01823_),
    .Q(\cpuregs[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15488_ (.CLK(clknet_leaf_59_clk),
    .D(_01824_),
    .Q(\cpuregs[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15489_ (.CLK(clknet_leaf_56_clk),
    .D(_01825_),
    .Q(\cpuregs[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15490_ (.CLK(clknet_leaf_51_clk),
    .D(_01826_),
    .Q(\cpuregs[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15491_ (.CLK(clknet_leaf_53_clk),
    .D(_01827_),
    .Q(\cpuregs[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15492_ (.CLK(clknet_leaf_59_clk),
    .D(_01828_),
    .Q(\cpuregs[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15493_ (.CLK(clknet_leaf_54_clk),
    .D(_01829_),
    .Q(\cpuregs[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15494_ (.CLK(clknet_leaf_56_clk),
    .D(_01830_),
    .Q(\cpuregs[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _15495_ (.CLK(clknet_leaf_131_clk),
    .D(_01831_),
    .Q(net203));
 sky130_fd_sc_hd__dfxtp_1 _15496_ (.CLK(clknet_leaf_131_clk),
    .D(_01832_),
    .Q(net214));
 sky130_fd_sc_hd__dfxtp_2 _15497_ (.CLK(clknet_leaf_132_clk),
    .D(_01833_),
    .Q(net225));
 sky130_fd_sc_hd__dfxtp_2 _15498_ (.CLK(clknet_leaf_132_clk),
    .D(_01834_),
    .Q(net228));
 sky130_fd_sc_hd__dfxtp_2 _15499_ (.CLK(clknet_leaf_133_clk),
    .D(_01835_),
    .Q(net229));
 sky130_fd_sc_hd__dfxtp_1 _15500_ (.CLK(clknet_leaf_133_clk),
    .D(_01836_),
    .Q(net230));
 sky130_fd_sc_hd__dfxtp_2 _15501_ (.CLK(clknet_leaf_174_clk),
    .D(_01837_),
    .Q(net231));
 sky130_fd_sc_hd__dfxtp_1 _15502_ (.CLK(clknet_leaf_171_clk),
    .D(_01838_),
    .Q(net232));
 sky130_fd_sc_hd__dfxtp_1 _15503_ (.CLK(clknet_leaf_171_clk),
    .D(_01839_),
    .Q(net233));
 sky130_fd_sc_hd__dfxtp_1 _15504_ (.CLK(clknet_leaf_167_clk),
    .D(_01840_),
    .Q(net234));
 sky130_fd_sc_hd__dfxtp_1 _15505_ (.CLK(clknet_leaf_172_clk),
    .D(_01841_),
    .Q(net204));
 sky130_fd_sc_hd__dfxtp_1 _15506_ (.CLK(clknet_leaf_167_clk),
    .D(_01842_),
    .Q(net205));
 sky130_fd_sc_hd__dfxtp_1 _15507_ (.CLK(clknet_leaf_167_clk),
    .D(_01843_),
    .Q(net206));
 sky130_fd_sc_hd__dfxtp_1 _15508_ (.CLK(clknet_leaf_173_clk),
    .D(_01844_),
    .Q(net207));
 sky130_fd_sc_hd__dfxtp_1 _15509_ (.CLK(clknet_leaf_167_clk),
    .D(_01845_),
    .Q(net208));
 sky130_fd_sc_hd__dfxtp_1 _15510_ (.CLK(clknet_leaf_173_clk),
    .D(_01846_),
    .Q(net209));
 sky130_fd_sc_hd__dfxtp_1 _15511_ (.CLK(clknet_leaf_175_clk),
    .D(_01847_),
    .Q(net210));
 sky130_fd_sc_hd__dfxtp_1 _15512_ (.CLK(clknet_leaf_175_clk),
    .D(_01848_),
    .Q(net211));
 sky130_fd_sc_hd__dfxtp_1 _15513_ (.CLK(clknet_leaf_175_clk),
    .D(_01849_),
    .Q(net212));
 sky130_fd_sc_hd__dfxtp_1 _15514_ (.CLK(clknet_leaf_78_clk),
    .D(_01850_),
    .Q(net213));
 sky130_fd_sc_hd__dfxtp_1 _15515_ (.CLK(clknet_leaf_78_clk),
    .D(_01851_),
    .Q(net215));
 sky130_fd_sc_hd__dfxtp_1 _15516_ (.CLK(clknet_leaf_79_clk),
    .D(_01852_),
    .Q(net216));
 sky130_fd_sc_hd__dfxtp_1 _15517_ (.CLK(clknet_leaf_81_clk),
    .D(_01853_),
    .Q(net217));
 sky130_fd_sc_hd__dfxtp_1 _15518_ (.CLK(clknet_leaf_79_clk),
    .D(_01854_),
    .Q(net218));
 sky130_fd_sc_hd__dfxtp_1 _15519_ (.CLK(clknet_leaf_81_clk),
    .D(_01855_),
    .Q(net219));
 sky130_fd_sc_hd__dfxtp_1 _15520_ (.CLK(clknet_leaf_81_clk),
    .D(_01856_),
    .Q(net220));
 sky130_fd_sc_hd__dfxtp_1 _15521_ (.CLK(clknet_leaf_75_clk),
    .D(_01857_),
    .Q(net221));
 sky130_fd_sc_hd__dfxtp_1 _15522_ (.CLK(clknet_leaf_86_clk),
    .D(_01858_),
    .Q(net222));
 sky130_fd_sc_hd__dfxtp_1 _15523_ (.CLK(clknet_leaf_86_clk),
    .D(_01859_),
    .Q(net223));
 sky130_fd_sc_hd__dfxtp_1 _15524_ (.CLK(clknet_leaf_86_clk),
    .D(_01860_),
    .Q(net224));
 sky130_fd_sc_hd__dfxtp_1 _15525_ (.CLK(clknet_leaf_86_clk),
    .D(_01861_),
    .Q(net226));
 sky130_fd_sc_hd__dfxtp_1 _15526_ (.CLK(clknet_leaf_39_clk),
    .D(_01862_),
    .Q(\cpuregs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15527_ (.CLK(clknet_leaf_45_clk),
    .D(_01863_),
    .Q(\cpuregs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15528_ (.CLK(clknet_leaf_31_clk),
    .D(_01864_),
    .Q(\cpuregs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15529_ (.CLK(clknet_leaf_19_clk),
    .D(_01865_),
    .Q(\cpuregs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15530_ (.CLK(clknet_leaf_29_clk),
    .D(_01866_),
    .Q(\cpuregs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15531_ (.CLK(clknet_leaf_22_clk),
    .D(_01867_),
    .Q(\cpuregs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15532_ (.CLK(clknet_leaf_21_clk),
    .D(_01868_),
    .Q(\cpuregs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15533_ (.CLK(clknet_leaf_20_clk),
    .D(_01869_),
    .Q(\cpuregs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15534_ (.CLK(clknet_leaf_182_clk),
    .D(_01870_),
    .Q(\cpuregs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15535_ (.CLK(clknet_leaf_181_clk),
    .D(_01871_),
    .Q(\cpuregs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15536_ (.CLK(clknet_leaf_193_clk),
    .D(_01872_),
    .Q(\cpuregs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15537_ (.CLK(clknet_leaf_193_clk),
    .D(_01873_),
    .Q(\cpuregs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15538_ (.CLK(clknet_leaf_3_clk),
    .D(_01874_),
    .Q(\cpuregs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15539_ (.CLK(clknet_leaf_3_clk),
    .D(_01875_),
    .Q(\cpuregs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15540_ (.CLK(clknet_leaf_194_clk),
    .D(_01876_),
    .Q(\cpuregs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15541_ (.CLK(clknet_leaf_1_clk),
    .D(_01877_),
    .Q(\cpuregs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15542_ (.CLK(clknet_leaf_10_clk),
    .D(_01878_),
    .Q(\cpuregs[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15543_ (.CLK(clknet_leaf_9_clk),
    .D(_01879_),
    .Q(\cpuregs[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15544_ (.CLK(clknet_leaf_9_clk),
    .D(_01880_),
    .Q(\cpuregs[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15545_ (.CLK(clknet_leaf_42_clk),
    .D(_01881_),
    .Q(\cpuregs[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15546_ (.CLK(clknet_leaf_12_clk),
    .D(_01882_),
    .Q(\cpuregs[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15547_ (.CLK(clknet_leaf_15_clk),
    .D(_01883_),
    .Q(\cpuregs[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15548_ (.CLK(clknet_leaf_43_clk),
    .D(_01884_),
    .Q(\cpuregs[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15549_ (.CLK(clknet_leaf_17_clk),
    .D(_01885_),
    .Q(\cpuregs[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15550_ (.CLK(clknet_leaf_35_clk),
    .D(_01886_),
    .Q(\cpuregs[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15551_ (.CLK(clknet_leaf_58_clk),
    .D(_01887_),
    .Q(\cpuregs[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15552_ (.CLK(clknet_leaf_57_clk),
    .D(_01888_),
    .Q(\cpuregs[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15553_ (.CLK(clknet_leaf_50_clk),
    .D(_01889_),
    .Q(\cpuregs[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15554_ (.CLK(clknet_leaf_53_clk),
    .D(_01890_),
    .Q(\cpuregs[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15555_ (.CLK(clknet_leaf_59_clk),
    .D(_01891_),
    .Q(\cpuregs[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15556_ (.CLK(clknet_leaf_54_clk),
    .D(_01892_),
    .Q(\cpuregs[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15557_ (.CLK(clknet_leaf_56_clk),
    .D(_01893_),
    .Q(\cpuregs[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15558_ (.CLK(clknet_leaf_39_clk),
    .D(_01894_),
    .Q(\cpuregs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15559_ (.CLK(clknet_leaf_45_clk),
    .D(_01895_),
    .Q(\cpuregs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15560_ (.CLK(clknet_leaf_31_clk),
    .D(_01896_),
    .Q(\cpuregs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15561_ (.CLK(clknet_leaf_19_clk),
    .D(_01897_),
    .Q(\cpuregs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15562_ (.CLK(clknet_leaf_29_clk),
    .D(_01898_),
    .Q(\cpuregs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15563_ (.CLK(clknet_leaf_22_clk),
    .D(_01899_),
    .Q(\cpuregs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15564_ (.CLK(clknet_leaf_21_clk),
    .D(_01900_),
    .Q(\cpuregs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15565_ (.CLK(clknet_leaf_20_clk),
    .D(_01901_),
    .Q(\cpuregs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15566_ (.CLK(clknet_leaf_182_clk),
    .D(_01902_),
    .Q(\cpuregs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15567_ (.CLK(clknet_leaf_182_clk),
    .D(_01903_),
    .Q(\cpuregs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15568_ (.CLK(clknet_leaf_193_clk),
    .D(_01904_),
    .Q(\cpuregs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15569_ (.CLK(clknet_leaf_193_clk),
    .D(_01905_),
    .Q(\cpuregs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15570_ (.CLK(clknet_leaf_3_clk),
    .D(_01906_),
    .Q(\cpuregs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15571_ (.CLK(clknet_leaf_3_clk),
    .D(_01907_),
    .Q(\cpuregs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15572_ (.CLK(clknet_leaf_194_clk),
    .D(_01908_),
    .Q(\cpuregs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15573_ (.CLK(clknet_leaf_1_clk),
    .D(_01909_),
    .Q(\cpuregs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15574_ (.CLK(clknet_leaf_12_clk),
    .D(_01910_),
    .Q(\cpuregs[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15575_ (.CLK(clknet_leaf_9_clk),
    .D(_01911_),
    .Q(\cpuregs[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15576_ (.CLK(clknet_leaf_9_clk),
    .D(_01912_),
    .Q(\cpuregs[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15577_ (.CLK(clknet_leaf_42_clk),
    .D(_01913_),
    .Q(\cpuregs[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15578_ (.CLK(clknet_leaf_12_clk),
    .D(_01914_),
    .Q(\cpuregs[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15579_ (.CLK(clknet_leaf_15_clk),
    .D(_01915_),
    .Q(\cpuregs[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15580_ (.CLK(clknet_leaf_42_clk),
    .D(_01916_),
    .Q(\cpuregs[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15581_ (.CLK(clknet_leaf_17_clk),
    .D(_01917_),
    .Q(\cpuregs[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15582_ (.CLK(clknet_leaf_35_clk),
    .D(_01918_),
    .Q(\cpuregs[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15583_ (.CLK(clknet_leaf_58_clk),
    .D(_01919_),
    .Q(\cpuregs[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15584_ (.CLK(clknet_leaf_57_clk),
    .D(_01920_),
    .Q(\cpuregs[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15585_ (.CLK(clknet_leaf_50_clk),
    .D(_01921_),
    .Q(\cpuregs[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15586_ (.CLK(clknet_leaf_53_clk),
    .D(_01922_),
    .Q(\cpuregs[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15587_ (.CLK(clknet_leaf_59_clk),
    .D(_01923_),
    .Q(\cpuregs[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15588_ (.CLK(clknet_leaf_54_clk),
    .D(_01924_),
    .Q(\cpuregs[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15589_ (.CLK(clknet_leaf_57_clk),
    .D(_01925_),
    .Q(\cpuregs[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15590_ (.CLK(clknet_leaf_36_clk),
    .D(_01926_),
    .Q(\cpuregs[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15591_ (.CLK(clknet_leaf_45_clk),
    .D(_01927_),
    .Q(\cpuregs[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15592_ (.CLK(clknet_leaf_31_clk),
    .D(_01928_),
    .Q(\cpuregs[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15593_ (.CLK(clknet_leaf_22_clk),
    .D(_01929_),
    .Q(\cpuregs[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15594_ (.CLK(clknet_leaf_29_clk),
    .D(_01930_),
    .Q(\cpuregs[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15595_ (.CLK(clknet_leaf_21_clk),
    .D(_01931_),
    .Q(\cpuregs[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15596_ (.CLK(clknet_leaf_180_clk),
    .D(_01932_),
    .Q(\cpuregs[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15597_ (.CLK(clknet_leaf_192_clk),
    .D(_01933_),
    .Q(\cpuregs[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15598_ (.CLK(clknet_leaf_183_clk),
    .D(_01934_),
    .Q(\cpuregs[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15599_ (.CLK(clknet_leaf_182_clk),
    .D(_01935_),
    .Q(\cpuregs[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15600_ (.CLK(clknet_leaf_190_clk),
    .D(_01936_),
    .Q(\cpuregs[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15601_ (.CLK(clknet_leaf_191_clk),
    .D(_01937_),
    .Q(\cpuregs[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15602_ (.CLK(clknet_leaf_198_clk),
    .D(_01938_),
    .Q(\cpuregs[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15603_ (.CLK(clknet_leaf_196_clk),
    .D(_01939_),
    .Q(\cpuregs[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15604_ (.CLK(clknet_leaf_197_clk),
    .D(_01940_),
    .Q(\cpuregs[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15605_ (.CLK(clknet_leaf_199_clk),
    .D(_01941_),
    .Q(\cpuregs[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15606_ (.CLK(clknet_leaf_10_clk),
    .D(_01942_),
    .Q(\cpuregs[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15607_ (.CLK(clknet_leaf_0_clk),
    .D(_01943_),
    .Q(\cpuregs[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15608_ (.CLK(clknet_leaf_1_clk),
    .D(_01944_),
    .Q(\cpuregs[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15609_ (.CLK(clknet_leaf_42_clk),
    .D(_01945_),
    .Q(\cpuregs[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15610_ (.CLK(clknet_leaf_12_clk),
    .D(_01946_),
    .Q(\cpuregs[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15611_ (.CLK(clknet_leaf_13_clk),
    .D(_01947_),
    .Q(\cpuregs[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15612_ (.CLK(clknet_leaf_45_clk),
    .D(_01948_),
    .Q(\cpuregs[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15613_ (.CLK(clknet_leaf_16_clk),
    .D(_01949_),
    .Q(\cpuregs[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15614_ (.CLK(clknet_leaf_35_clk),
    .D(_01950_),
    .Q(\cpuregs[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15615_ (.CLK(clknet_leaf_71_clk),
    .D(_01951_),
    .Q(\cpuregs[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15616_ (.CLK(clknet_leaf_34_clk),
    .D(_01952_),
    .Q(\cpuregs[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15617_ (.CLK(clknet_leaf_48_clk),
    .D(_01953_),
    .Q(\cpuregs[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15618_ (.CLK(clknet_leaf_46_clk),
    .D(_01954_),
    .Q(\cpuregs[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15619_ (.CLK(clknet_4_11_0_clk),
    .D(_01955_),
    .Q(\cpuregs[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15620_ (.CLK(clknet_leaf_53_clk),
    .D(_01956_),
    .Q(\cpuregs[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15621_ (.CLK(clknet_leaf_49_clk),
    .D(_01957_),
    .Q(\cpuregs[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15622_ (.CLK(clknet_leaf_36_clk),
    .D(_01958_),
    .Q(\cpuregs[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15623_ (.CLK(clknet_leaf_45_clk),
    .D(_01959_),
    .Q(\cpuregs[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15624_ (.CLK(clknet_leaf_31_clk),
    .D(_01960_),
    .Q(\cpuregs[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15625_ (.CLK(clknet_leaf_22_clk),
    .D(_01961_),
    .Q(\cpuregs[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15626_ (.CLK(clknet_leaf_29_clk),
    .D(_01962_),
    .Q(\cpuregs[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15627_ (.CLK(clknet_leaf_21_clk),
    .D(_01963_),
    .Q(\cpuregs[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15628_ (.CLK(clknet_leaf_178_clk),
    .D(_01964_),
    .Q(\cpuregs[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15629_ (.CLK(clknet_leaf_192_clk),
    .D(_01965_),
    .Q(\cpuregs[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15630_ (.CLK(clknet_leaf_183_clk),
    .D(_01966_),
    .Q(\cpuregs[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15631_ (.CLK(clknet_leaf_182_clk),
    .D(_01967_),
    .Q(\cpuregs[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15632_ (.CLK(clknet_leaf_190_clk),
    .D(_01968_),
    .Q(\cpuregs[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15633_ (.CLK(clknet_leaf_191_clk),
    .D(_01969_),
    .Q(\cpuregs[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15634_ (.CLK(clknet_leaf_198_clk),
    .D(_01970_),
    .Q(\cpuregs[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15635_ (.CLK(clknet_leaf_196_clk),
    .D(_01971_),
    .Q(\cpuregs[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15636_ (.CLK(clknet_leaf_191_clk),
    .D(_01972_),
    .Q(\cpuregs[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15637_ (.CLK(clknet_leaf_199_clk),
    .D(_01973_),
    .Q(\cpuregs[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15638_ (.CLK(clknet_leaf_10_clk),
    .D(_01974_),
    .Q(\cpuregs[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15639_ (.CLK(clknet_leaf_0_clk),
    .D(_01975_),
    .Q(\cpuregs[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15640_ (.CLK(clknet_leaf_1_clk),
    .D(_01976_),
    .Q(\cpuregs[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15641_ (.CLK(clknet_leaf_41_clk),
    .D(_01977_),
    .Q(\cpuregs[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15642_ (.CLK(clknet_leaf_12_clk),
    .D(_01978_),
    .Q(\cpuregs[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15643_ (.CLK(clknet_leaf_13_clk),
    .D(_01979_),
    .Q(\cpuregs[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15644_ (.CLK(clknet_leaf_45_clk),
    .D(_01980_),
    .Q(\cpuregs[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15645_ (.CLK(clknet_leaf_16_clk),
    .D(_01981_),
    .Q(\cpuregs[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15646_ (.CLK(clknet_leaf_35_clk),
    .D(_01982_),
    .Q(\cpuregs[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15647_ (.CLK(clknet_leaf_71_clk),
    .D(_01983_),
    .Q(\cpuregs[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15648_ (.CLK(clknet_leaf_34_clk),
    .D(_01984_),
    .Q(\cpuregs[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15649_ (.CLK(clknet_leaf_49_clk),
    .D(_01985_),
    .Q(\cpuregs[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15650_ (.CLK(clknet_leaf_46_clk),
    .D(_01986_),
    .Q(\cpuregs[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15651_ (.CLK(clknet_leaf_70_clk),
    .D(_01987_),
    .Q(\cpuregs[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15652_ (.CLK(clknet_leaf_53_clk),
    .D(_01988_),
    .Q(\cpuregs[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15653_ (.CLK(clknet_leaf_49_clk),
    .D(_01989_),
    .Q(\cpuregs[17][31] ));
 sky130_fd_sc_hd__conb_1 picorv32_1243 (.LO(net1243));
 sky130_fd_sc_hd__conb_1 picorv32_1244 (.LO(net1244));
 sky130_fd_sc_hd__conb_1 picorv32_1245 (.LO(net1245));
 sky130_fd_sc_hd__conb_1 picorv32_1246 (.LO(net1246));
 sky130_fd_sc_hd__conb_1 picorv32_1247 (.LO(net1247));
 sky130_fd_sc_hd__conb_1 picorv32_1248 (.LO(net1248));
 sky130_fd_sc_hd__conb_1 picorv32_1249 (.LO(net1249));
 sky130_fd_sc_hd__conb_1 picorv32_1250 (.LO(net1250));
 sky130_fd_sc_hd__conb_1 picorv32_1251 (.LO(net1251));
 sky130_fd_sc_hd__conb_1 picorv32_1252 (.LO(net1252));
 sky130_fd_sc_hd__conb_1 picorv32_1253 (.LO(net1253));
 sky130_fd_sc_hd__conb_1 picorv32_1254 (.LO(net1254));
 sky130_fd_sc_hd__conb_1 picorv32_1255 (.LO(net1255));
 sky130_fd_sc_hd__conb_1 picorv32_1256 (.LO(net1256));
 sky130_fd_sc_hd__conb_1 picorv32_1257 (.LO(net1257));
 sky130_fd_sc_hd__conb_1 picorv32_1258 (.LO(net1258));
 sky130_fd_sc_hd__conb_1 picorv32_1259 (.LO(net1259));
 sky130_fd_sc_hd__conb_1 picorv32_1260 (.LO(net1260));
 sky130_fd_sc_hd__conb_1 picorv32_1261 (.LO(net1261));
 sky130_fd_sc_hd__conb_1 picorv32_1262 (.LO(net1262));
 sky130_fd_sc_hd__conb_1 picorv32_1263 (.LO(net1263));
 sky130_fd_sc_hd__conb_1 picorv32_1264 (.LO(net1264));
 sky130_fd_sc_hd__conb_1 picorv32_1265 (.LO(net1265));
 sky130_fd_sc_hd__conb_1 picorv32_1266 (.LO(net1266));
 sky130_fd_sc_hd__conb_1 picorv32_1267 (.LO(net1267));
 sky130_fd_sc_hd__conb_1 picorv32_1268 (.LO(net1268));
 sky130_fd_sc_hd__conb_1 picorv32_1269 (.LO(net1269));
 sky130_fd_sc_hd__conb_1 picorv32_1270 (.LO(net1270));
 sky130_fd_sc_hd__conb_1 picorv32_1271 (.LO(net1271));
 sky130_fd_sc_hd__conb_1 picorv32_1272 (.LO(net1272));
 sky130_fd_sc_hd__conb_1 picorv32_1273 (.LO(net1273));
 sky130_fd_sc_hd__conb_1 picorv32_1274 (.LO(net1274));
 sky130_fd_sc_hd__conb_1 picorv32_1275 (.LO(net1275));
 sky130_fd_sc_hd__conb_1 picorv32_1276 (.LO(net1276));
 sky130_fd_sc_hd__conb_1 picorv32_1277 (.LO(net1277));
 sky130_fd_sc_hd__conb_1 picorv32_1278 (.LO(net1278));
 sky130_fd_sc_hd__conb_1 picorv32_1279 (.LO(net1279));
 sky130_fd_sc_hd__conb_1 picorv32_1280 (.LO(net1280));
 sky130_fd_sc_hd__conb_1 picorv32_1281 (.LO(net1281));
 sky130_fd_sc_hd__conb_1 picorv32_1282 (.LO(net1282));
 sky130_fd_sc_hd__conb_1 picorv32_1283 (.LO(net1283));
 sky130_fd_sc_hd__conb_1 picorv32_1284 (.LO(net1284));
 sky130_fd_sc_hd__conb_1 picorv32_1285 (.LO(net1285));
 sky130_fd_sc_hd__conb_1 picorv32_1286 (.LO(net1286));
 sky130_fd_sc_hd__conb_1 picorv32_1287 (.LO(net1287));
 sky130_fd_sc_hd__conb_1 picorv32_1288 (.LO(net1288));
 sky130_fd_sc_hd__conb_1 picorv32_1289 (.LO(net1289));
 sky130_fd_sc_hd__conb_1 picorv32_1290 (.LO(net1290));
 sky130_fd_sc_hd__conb_1 picorv32_1291 (.LO(net1291));
 sky130_fd_sc_hd__conb_1 picorv32_1292 (.LO(net1292));
 sky130_fd_sc_hd__conb_1 picorv32_1293 (.LO(net1293));
 sky130_fd_sc_hd__conb_1 picorv32_1294 (.LO(net1294));
 sky130_fd_sc_hd__conb_1 picorv32_1295 (.LO(net1295));
 sky130_fd_sc_hd__conb_1 picorv32_1296 (.LO(net1296));
 sky130_fd_sc_hd__conb_1 picorv32_1297 (.LO(net1297));
 sky130_fd_sc_hd__conb_1 picorv32_1298 (.LO(net1298));
 sky130_fd_sc_hd__conb_1 picorv32_1299 (.LO(net1299));
 sky130_fd_sc_hd__conb_1 picorv32_1300 (.LO(net1300));
 sky130_fd_sc_hd__conb_1 picorv32_1301 (.LO(net1301));
 sky130_fd_sc_hd__conb_1 picorv32_1302 (.LO(net1302));
 sky130_fd_sc_hd__conb_1 picorv32_1303 (.LO(net1303));
 sky130_fd_sc_hd__conb_1 picorv32_1304 (.LO(net1304));
 sky130_fd_sc_hd__conb_1 picorv32_1305 (.LO(net1305));
 sky130_fd_sc_hd__conb_1 picorv32_1306 (.LO(net1306));
 sky130_fd_sc_hd__conb_1 picorv32_1307 (.LO(net1307));
 sky130_fd_sc_hd__conb_1 picorv32_1308 (.LO(net1308));
 sky130_fd_sc_hd__conb_1 picorv32_1309 (.LO(net1309));
 sky130_fd_sc_hd__conb_1 picorv32_1310 (.LO(net1310));
 sky130_fd_sc_hd__conb_1 picorv32_1311 (.LO(net1311));
 sky130_fd_sc_hd__conb_1 picorv32_1312 (.LO(net1312));
 sky130_fd_sc_hd__conb_1 picorv32_1313 (.LO(net1313));
 sky130_fd_sc_hd__conb_1 picorv32_1314 (.LO(net1314));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_1 _15727_ (.A(net1181),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 _15728_ (.A(net1179),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 _15729_ (.A(net119),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 _15730_ (.A(net122),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 _15731_ (.A(net1175),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 _15732_ (.A(net1173),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 _15733_ (.A(net125),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 _15734_ (.A(net1169),
    .X(net264));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3455 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(mem_rdata[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(mem_rdata[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(mem_rdata[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(mem_rdata[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(mem_rdata[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(mem_rdata[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(mem_rdata[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(mem_rdata[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(mem_rdata[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(mem_rdata[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(mem_rdata[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(mem_rdata[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(mem_rdata[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(mem_rdata[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(mem_rdata[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(mem_rdata[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(mem_rdata[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(mem_rdata[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(mem_rdata[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(mem_rdata[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(mem_rdata[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(mem_rdata[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(mem_rdata[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(mem_rdata[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(mem_rdata[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(mem_rdata[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(mem_rdata[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(mem_rdata[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(mem_rdata[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(mem_rdata[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(mem_rdata[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(mem_rdata[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(mem_ready),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(resetn),
    .X(net34));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(mem_instr));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(mem_la_read));
 sky130_fd_sc_hd__buf_2 output97 (.A(net1180),
    .X(mem_la_wdata[0]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net1179),
    .X(mem_la_wdata[1]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net1177),
    .X(mem_la_wdata[2]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net1176),
    .X(mem_la_wdata[3]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net1174),
    .X(mem_la_wdata[4]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net1173),
    .X(mem_la_wdata[5]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(mem_la_wdata[6]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net1170),
    .X(mem_la_wdata[7]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(mem_la_write));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(mem_la_wstrb[1]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(mem_valid));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(pcpi_insn[0]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(pcpi_insn[10]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(pcpi_insn[11]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(pcpi_insn[12]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(pcpi_insn[13]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(pcpi_insn[14]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(pcpi_insn[15]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(pcpi_insn[16]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(pcpi_insn[17]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(pcpi_insn[18]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(pcpi_insn[19]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(pcpi_insn[1]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(pcpi_insn[20]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(pcpi_insn[21]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(pcpi_insn[22]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(pcpi_insn[23]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(pcpi_insn[24]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(pcpi_insn[25]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(pcpi_insn[26]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(pcpi_insn[27]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(pcpi_insn[28]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(pcpi_insn[29]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(pcpi_insn[2]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(pcpi_insn[30]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(pcpi_insn[31]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(pcpi_insn[3]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(pcpi_insn[4]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(pcpi_insn[5]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(pcpi_insn[6]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(pcpi_insn[7]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(pcpi_insn[8]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(pcpi_insn[9]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(pcpi_rs1[0]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(pcpi_rs1[10]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(pcpi_rs1[11]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net1027),
    .X(pcpi_rs1[12]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net1025),
    .X(pcpi_rs1[13]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net1023),
    .X(pcpi_rs1[14]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net1021),
    .X(pcpi_rs1[15]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net1019),
    .X(pcpi_rs1[16]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net1016),
    .X(pcpi_rs1[17]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net1015),
    .X(pcpi_rs1[18]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net1013),
    .X(pcpi_rs1[19]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net1050),
    .X(pcpi_rs1[1]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net1011),
    .X(pcpi_rs1[20]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net1009),
    .X(pcpi_rs1[21]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net1008),
    .X(pcpi_rs1[22]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net1006),
    .X(pcpi_rs1[23]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net1005),
    .X(pcpi_rs1[24]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net1003),
    .X(pcpi_rs1[25]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net1001),
    .X(pcpi_rs1[26]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net999),
    .X(pcpi_rs1[27]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net997),
    .X(pcpi_rs1[28]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net995),
    .X(pcpi_rs1[29]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(pcpi_rs1[2]));
 sky130_fd_sc_hd__buf_2 output226 (.A(net993),
    .X(pcpi_rs1[30]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net1189),
    .X(pcpi_rs1[31]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(pcpi_rs1[3]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(pcpi_rs1[4]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net1041),
    .X(pcpi_rs1[5]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(pcpi_rs1[6]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net1037),
    .X(pcpi_rs1[7]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net1034),
    .X(pcpi_rs1[8]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(pcpi_rs1[9]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(pcpi_rs2[10]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(pcpi_rs2[11]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(pcpi_rs2[12]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net1163),
    .X(pcpi_rs2[13]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(pcpi_rs2[14]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net1162),
    .X(pcpi_rs2[15]));
 sky130_fd_sc_hd__buf_2 output242 (.A(net242),
    .X(pcpi_rs2[16]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(pcpi_rs2[17]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(pcpi_rs2[18]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(pcpi_rs2[19]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(pcpi_rs2[20]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(pcpi_rs2[21]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(pcpi_rs2[22]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(pcpi_rs2[23]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(pcpi_rs2[24]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(pcpi_rs2[25]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(pcpi_rs2[26]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(pcpi_rs2[27]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(pcpi_rs2[28]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(pcpi_rs2[29]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(pcpi_rs2[30]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(pcpi_rs2[31]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net1168),
    .X(pcpi_rs2[8]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net1167),
    .X(pcpi_rs2[9]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(pcpi_valid));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(trap));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net272),
    .X(net269));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout270 (.A(net272),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 fanout272 (.A(_06403_),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(net275),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(_06403_),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(_06403_),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 fanout278 (.A(_03873_),
    .X(net278));
 sky130_fd_sc_hd__buf_1 fanout279 (.A(_03873_),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 fanout280 (.A(_03873_),
    .X(net280));
 sky130_fd_sc_hd__buf_1 fanout281 (.A(_03873_),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(_03870_),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 fanout284 (.A(_03870_),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 fanout286 (.A(net288),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout288 (.A(_03865_),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 fanout289 (.A(_03860_),
    .X(net289));
 sky130_fd_sc_hd__buf_1 fanout290 (.A(_03860_),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 fanout291 (.A(_03860_),
    .X(net291));
 sky130_fd_sc_hd__buf_1 fanout292 (.A(_03860_),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(_03857_),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 fanout294 (.A(_03857_),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 fanout296 (.A(_03857_),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(_03852_),
    .X(net297));
 sky130_fd_sc_hd__buf_1 fanout298 (.A(_03852_),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 fanout299 (.A(_03852_),
    .X(net299));
 sky130_fd_sc_hd__buf_1 fanout300 (.A(_03852_),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 fanout301 (.A(_03849_),
    .X(net301));
 sky130_fd_sc_hd__buf_1 fanout302 (.A(_03849_),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 fanout304 (.A(_03849_),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 fanout305 (.A(_03844_),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_2 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 fanout307 (.A(_03844_),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 fanout308 (.A(net311),
    .X(net308));
 sky130_fd_sc_hd__buf_1 fanout309 (.A(net311),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 fanout311 (.A(_03839_),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 fanout312 (.A(net315),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 fanout313 (.A(net315),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout315 (.A(_03836_),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_2 fanout316 (.A(net319),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 fanout319 (.A(_03831_),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 fanout320 (.A(_03826_),
    .X(net320));
 sky130_fd_sc_hd__buf_1 fanout321 (.A(_03826_),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_2 fanout322 (.A(_03826_),
    .X(net322));
 sky130_fd_sc_hd__buf_1 fanout323 (.A(_03826_),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 fanout325 (.A(net327),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout327 (.A(_03823_),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 fanout328 (.A(_03818_),
    .X(net328));
 sky130_fd_sc_hd__buf_1 fanout329 (.A(_03818_),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 fanout330 (.A(_03818_),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 fanout331 (.A(_03818_),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout333 (.A(_03815_),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_2 fanout334 (.A(_03815_),
    .X(net334));
 sky130_fd_sc_hd__buf_1 fanout335 (.A(_03815_),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 fanout337 (.A(_03810_),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 fanout338 (.A(_03810_),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 fanout339 (.A(_03807_),
    .X(net339));
 sky130_fd_sc_hd__buf_1 fanout340 (.A(_03807_),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 fanout341 (.A(_03807_),
    .X(net341));
 sky130_fd_sc_hd__buf_1 fanout342 (.A(_03807_),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__buf_1 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 fanout345 (.A(_03802_),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 fanout346 (.A(_03802_),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_2 fanout348 (.A(_03799_),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_2 fanout349 (.A(_03799_),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 fanout351 (.A(net353),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout353 (.A(_03794_),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout355 (.A(net357),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 fanout356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 fanout357 (.A(_03791_),
    .X(net357));
 sky130_fd_sc_hd__buf_2 fanout358 (.A(_02914_),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 fanout359 (.A(_02914_),
    .X(net359));
 sky130_fd_sc_hd__buf_4 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_8 fanout361 (.A(net363),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_8 fanout362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__buf_4 fanout363 (.A(_06662_),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 fanout364 (.A(net370),
    .X(net364));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout365 (.A(net370),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_4 fanout366 (.A(net370),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 fanout367 (.A(net370),
    .X(net367));
 sky130_fd_sc_hd__buf_2 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_4 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout370 (.A(_06578_),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_4 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 fanout372 (.A(_06578_),
    .X(net372));
 sky130_fd_sc_hd__buf_4 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_8 fanout374 (.A(net376),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_8 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_4 fanout376 (.A(_06234_),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_4 fanout377 (.A(net384),
    .X(net377));
 sky130_fd_sc_hd__buf_2 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_2 fanout379 (.A(net384),
    .X(net379));
 sky130_fd_sc_hd__buf_2 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__buf_2 fanout381 (.A(net384),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_4 fanout382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_2 fanout384 (.A(net390),
    .X(net384));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(net388),
    .X(net385));
 sky130_fd_sc_hd__buf_2 fanout386 (.A(net388),
    .X(net386));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout388 (.A(net390),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_4 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_2 fanout390 (.A(_05097_),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_4 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(_04888_),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_4 fanout393 (.A(_04888_),
    .X(net393));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout394 (.A(_04888_),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_4 fanout395 (.A(net398),
    .X(net395));
 sky130_fd_sc_hd__buf_2 fanout396 (.A(net398),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_4 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_2 fanout398 (.A(_04887_),
    .X(net398));
 sky130_fd_sc_hd__buf_4 fanout399 (.A(_04293_),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_4 fanout400 (.A(_04293_),
    .X(net400));
 sky130_fd_sc_hd__buf_4 fanout401 (.A(_04293_),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_4 fanout402 (.A(_04293_),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 fanout404 (.A(_03785_),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(_03785_),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 fanout406 (.A(_03785_),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 fanout409 (.A(_03782_),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_2 max_cap410 (.A(_02455_),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_8 fanout411 (.A(_02358_),
    .X(net411));
 sky130_fd_sc_hd__buf_2 fanout412 (.A(_02358_),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(_02358_),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_4 fanout414 (.A(_02358_),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 fanout415 (.A(_02357_),
    .X(net415));
 sky130_fd_sc_hd__buf_2 fanout416 (.A(_02357_),
    .X(net416));
 sky130_fd_sc_hd__buf_4 fanout417 (.A(_02357_),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_4 fanout418 (.A(_02357_),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_8 fanout419 (.A(net422),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_4 fanout420 (.A(net422),
    .X(net420));
 sky130_fd_sc_hd__buf_4 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__buf_4 fanout422 (.A(_02356_),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_8 fanout423 (.A(net426),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_4 fanout424 (.A(net426),
    .X(net424));
 sky130_fd_sc_hd__buf_4 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_4 fanout426 (.A(_02355_),
    .X(net426));
 sky130_fd_sc_hd__buf_4 fanout427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_4 fanout428 (.A(net430),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_8 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_4 fanout430 (.A(_02129_),
    .X(net430));
 sky130_fd_sc_hd__buf_4 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_4 fanout432 (.A(net434),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_8 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_4 fanout434 (.A(_02128_),
    .X(net434));
 sky130_fd_sc_hd__buf_4 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_4 fanout436 (.A(net438),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_8 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_4 fanout438 (.A(_02126_),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_4 fanout440 (.A(net442),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_8 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_4 fanout442 (.A(_02125_),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_4 fanout444 (.A(net446),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_8 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 fanout446 (.A(_02124_),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_8 fanout448 (.A(net450),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_8 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_4 fanout450 (.A(_02123_),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_4 fanout452 (.A(net454),
    .X(net452));
 sky130_fd_sc_hd__buf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_2 fanout454 (.A(_02122_),
    .X(net454));
 sky130_fd_sc_hd__buf_4 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_4 fanout456 (.A(_02119_),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(_02119_),
    .X(net457));
 sky130_fd_sc_hd__buf_2 fanout458 (.A(_02119_),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_8 fanout459 (.A(_02118_),
    .X(net459));
 sky130_fd_sc_hd__buf_2 fanout460 (.A(_02118_),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_8 fanout461 (.A(_02118_),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 fanout462 (.A(_02118_),
    .X(net462));
 sky130_fd_sc_hd__buf_4 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(_02117_),
    .X(net464));
 sky130_fd_sc_hd__buf_4 fanout465 (.A(_02117_),
    .X(net465));
 sky130_fd_sc_hd__buf_2 fanout466 (.A(_02117_),
    .X(net466));
 sky130_fd_sc_hd__buf_4 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_4 fanout468 (.A(_02051_),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_2 fanout470 (.A(_02051_),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_4 fanout472 (.A(_06664_),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_2 fanout474 (.A(_06664_),
    .X(net474));
 sky130_fd_sc_hd__buf_4 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_4 fanout476 (.A(_04292_),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_8 fanout477 (.A(_04292_),
    .X(net477));
 sky130_fd_sc_hd__buf_2 fanout478 (.A(_04292_),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_8 fanout479 (.A(net483),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_4 fanout480 (.A(net483),
    .X(net480));
 sky130_fd_sc_hd__buf_4 fanout481 (.A(_04291_),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_4 fanout482 (.A(_04291_),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_2 max_cap483 (.A(_04291_),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_8 fanout484 (.A(_04288_),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_4 fanout485 (.A(_04288_),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_8 fanout486 (.A(_04288_),
    .X(net486));
 sky130_fd_sc_hd__buf_4 fanout487 (.A(_04288_),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_8 fanout488 (.A(_04287_),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_4 fanout489 (.A(_04287_),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_8 fanout490 (.A(_04287_),
    .X(net490));
 sky130_fd_sc_hd__buf_4 fanout491 (.A(_04287_),
    .X(net491));
 sky130_fd_sc_hd__buf_4 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_4 fanout493 (.A(_04286_),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_8 fanout494 (.A(_04286_),
    .X(net494));
 sky130_fd_sc_hd__buf_2 fanout495 (.A(_04286_),
    .X(net495));
 sky130_fd_sc_hd__buf_4 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(net499),
    .X(net497));
 sky130_fd_sc_hd__buf_4 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_2 fanout499 (.A(_04285_),
    .X(net499));
 sky130_fd_sc_hd__buf_4 fanout500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_8 fanout501 (.A(net503),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_8 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_4 fanout503 (.A(_04284_),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_8 fanout504 (.A(_04279_),
    .X(net504));
 sky130_fd_sc_hd__buf_2 fanout505 (.A(_04279_),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_8 fanout506 (.A(_04279_),
    .X(net506));
 sky130_fd_sc_hd__buf_4 fanout507 (.A(_04279_),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_8 fanout508 (.A(_04278_),
    .X(net508));
 sky130_fd_sc_hd__buf_2 fanout509 (.A(_04278_),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_8 fanout510 (.A(_04278_),
    .X(net510));
 sky130_fd_sc_hd__buf_4 fanout511 (.A(_04278_),
    .X(net511));
 sky130_fd_sc_hd__buf_4 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__buf_4 fanout513 (.A(net515),
    .X(net513));
 sky130_fd_sc_hd__buf_4 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_4 fanout515 (.A(_04276_),
    .X(net515));
 sky130_fd_sc_hd__buf_4 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_4 fanout517 (.A(net519),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_8 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_4 fanout519 (.A(_04274_),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_2 fanout520 (.A(net523),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_2 fanout521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_2 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_2 fanout523 (.A(_03777_),
    .X(net523));
 sky130_fd_sc_hd__buf_2 fanout524 (.A(_03774_),
    .X(net524));
 sky130_fd_sc_hd__buf_1 fanout525 (.A(_03774_),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_2 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_1 fanout527 (.A(_03774_),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_8 fanout528 (.A(_03746_),
    .X(net528));
 sky130_fd_sc_hd__buf_2 fanout529 (.A(_03746_),
    .X(net529));
 sky130_fd_sc_hd__buf_4 fanout530 (.A(_03746_),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_4 fanout531 (.A(_03746_),
    .X(net531));
 sky130_fd_sc_hd__buf_2 fanout532 (.A(_06620_),
    .X(net532));
 sky130_fd_sc_hd__buf_4 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__buf_8 fanout534 (.A(_06240_),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_8 fanout535 (.A(_06240_),
    .X(net535));
 sky130_fd_sc_hd__buf_4 fanout536 (.A(_06240_),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_2 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__buf_1 fanout538 (.A(net540),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_2 fanout539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__buf_2 fanout540 (.A(_03769_),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 fanout541 (.A(net544),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 fanout542 (.A(net544),
    .X(net542));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout543 (.A(net544),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_2 fanout544 (.A(_03766_),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_4 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 fanout546 (.A(_03741_),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_4 fanout548 (.A(_03741_),
    .X(net548));
 sky130_fd_sc_hd__buf_4 fanout549 (.A(net551),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_2 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__buf_4 fanout551 (.A(_03198_),
    .X(net551));
 sky130_fd_sc_hd__buf_4 fanout552 (.A(_03156_),
    .X(net552));
 sky130_fd_sc_hd__buf_2 fanout553 (.A(_03156_),
    .X(net553));
 sky130_fd_sc_hd__buf_4 fanout554 (.A(_03156_),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_4 fanout555 (.A(_03156_),
    .X(net555));
 sky130_fd_sc_hd__buf_2 fanout556 (.A(net557),
    .X(net556));
 sky130_fd_sc_hd__buf_2 fanout557 (.A(_02133_),
    .X(net557));
 sky130_fd_sc_hd__buf_2 fanout558 (.A(_02133_),
    .X(net558));
 sky130_fd_sc_hd__buf_2 fanout559 (.A(_06622_),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_1 max_cap560 (.A(_06229_),
    .X(net560));
 sky130_fd_sc_hd__buf_2 fanout561 (.A(net563),
    .X(net561));
 sky130_fd_sc_hd__buf_1 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__buf_2 fanout563 (.A(_06174_),
    .X(net563));
 sky130_fd_sc_hd__buf_2 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_4 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_2 fanout566 (.A(_05080_),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_4 fanout567 (.A(net570),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_2 fanout568 (.A(net570),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_2 fanout570 (.A(_05040_),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_2 fanout571 (.A(_03761_),
    .X(net571));
 sky130_fd_sc_hd__buf_1 fanout572 (.A(_03761_),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_2 fanout573 (.A(_03761_),
    .X(net573));
 sky130_fd_sc_hd__buf_1 fanout574 (.A(_03761_),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_2 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__buf_1 fanout576 (.A(_03756_),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_2 fanout577 (.A(_03756_),
    .X(net577));
 sky130_fd_sc_hd__buf_1 fanout578 (.A(_03756_),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_2 fanout579 (.A(_03753_),
    .X(net579));
 sky130_fd_sc_hd__buf_1 fanout580 (.A(_03753_),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 fanout581 (.A(_03753_),
    .X(net581));
 sky130_fd_sc_hd__buf_1 fanout582 (.A(_03753_),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_2 fanout583 (.A(_03751_),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_2 fanout584 (.A(_03751_),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_2 fanout585 (.A(_03751_),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_2 fanout587 (.A(_03749_),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_2 fanout588 (.A(_03749_),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_4 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__buf_2 fanout590 (.A(net592),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_4 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_2 fanout592 (.A(net596),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_4 fanout593 (.A(net596),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 fanout594 (.A(net596),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_4 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__buf_2 fanout596 (.A(_03153_),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_4 fanout597 (.A(net600),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_4 fanout598 (.A(net600),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_2 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_4 fanout600 (.A(_03153_),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_4 fanout601 (.A(_03153_),
    .X(net601));
 sky130_fd_sc_hd__buf_2 fanout602 (.A(_03153_),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_4 fanout603 (.A(net606),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_2 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_4 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_4 fanout606 (.A(_03148_),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_4 fanout607 (.A(net609),
    .X(net607));
 sky130_fd_sc_hd__buf_2 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_4 fanout609 (.A(_03148_),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 fanout610 (.A(net616),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_2 fanout611 (.A(net616),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_4 fanout612 (.A(net616),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_2 fanout613 (.A(net616),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_4 fanout614 (.A(net616),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_4 fanout615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_4 fanout616 (.A(_03148_),
    .X(net616));
 sky130_fd_sc_hd__buf_2 fanout617 (.A(net620),
    .X(net617));
 sky130_fd_sc_hd__buf_2 fanout618 (.A(net620),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_4 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_2 fanout620 (.A(net645),
    .X(net620));
 sky130_fd_sc_hd__buf_2 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__buf_2 fanout622 (.A(net624),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_4 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_2 fanout624 (.A(net645),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_4 fanout625 (.A(net628),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_4 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__buf_2 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_2 fanout628 (.A(net631),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(net631),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout630 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_2 fanout631 (.A(net645),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_4 fanout632 (.A(net635),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_2 fanout633 (.A(net635),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_4 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_2 fanout635 (.A(net645),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(net639),
    .X(net636));
 sky130_fd_sc_hd__buf_2 fanout637 (.A(net639),
    .X(net637));
 sky130_fd_sc_hd__buf_2 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__buf_2 fanout639 (.A(net645),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_4 fanout640 (.A(net641),
    .X(net640));
 sky130_fd_sc_hd__buf_2 fanout641 (.A(net645),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_4 fanout642 (.A(net644),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_2 fanout643 (.A(net644),
    .X(net643));
 sky130_fd_sc_hd__buf_2 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_4 fanout645 (.A(_03140_),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_4 fanout646 (.A(net649),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_4 fanout647 (.A(net649),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 fanout648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_2 fanout649 (.A(net654),
    .X(net649));
 sky130_fd_sc_hd__buf_2 fanout650 (.A(net654),
    .X(net650));
 sky130_fd_sc_hd__buf_2 fanout651 (.A(net654),
    .X(net651));
 sky130_fd_sc_hd__buf_2 fanout652 (.A(net654),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_2 fanout653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_2 fanout654 (.A(net679),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_4 fanout655 (.A(net663),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_2 fanout656 (.A(net663),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_4 fanout657 (.A(net663),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_2 fanout658 (.A(net663),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_4 fanout659 (.A(net663),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_2 fanout660 (.A(net663),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_4 fanout661 (.A(net663),
    .X(net661));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_2 fanout663 (.A(net679),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_4 fanout664 (.A(net672),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_2 fanout665 (.A(net672),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_4 fanout666 (.A(net672),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_2 fanout667 (.A(net672),
    .X(net667));
 sky130_fd_sc_hd__buf_2 fanout668 (.A(net672),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_2 fanout669 (.A(net672),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_4 fanout670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__buf_2 fanout671 (.A(net672),
    .X(net671));
 sky130_fd_sc_hd__buf_2 fanout672 (.A(net679),
    .X(net672));
 sky130_fd_sc_hd__buf_2 fanout673 (.A(net676),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_2 fanout674 (.A(net676),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_4 fanout675 (.A(net676),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_2 fanout676 (.A(net679),
    .X(net676));
 sky130_fd_sc_hd__buf_2 fanout677 (.A(net679),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_2 fanout678 (.A(net679),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_4 fanout679 (.A(_03139_),
    .X(net679));
 sky130_fd_sc_hd__buf_2 fanout680 (.A(net696),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_2 fanout681 (.A(net696),
    .X(net681));
 sky130_fd_sc_hd__buf_2 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_2 fanout683 (.A(net696),
    .X(net683));
 sky130_fd_sc_hd__buf_2 fanout684 (.A(net687),
    .X(net684));
 sky130_fd_sc_hd__buf_2 fanout685 (.A(net687),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_4 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_2 fanout687 (.A(net696),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 fanout688 (.A(net691),
    .X(net688));
 sky130_fd_sc_hd__buf_2 fanout689 (.A(net691),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_2 fanout690 (.A(net691),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_2 fanout691 (.A(net696),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_4 fanout692 (.A(net695),
    .X(net692));
 sky130_fd_sc_hd__buf_2 fanout693 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__buf_2 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__buf_2 fanout695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_2 fanout696 (.A(net707),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_4 fanout697 (.A(net701),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_2 fanout698 (.A(net701),
    .X(net698));
 sky130_fd_sc_hd__buf_2 fanout699 (.A(net701),
    .X(net699));
 sky130_fd_sc_hd__buf_2 fanout700 (.A(net701),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_4 fanout701 (.A(net707),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_4 fanout702 (.A(net705),
    .X(net702));
 sky130_fd_sc_hd__buf_2 fanout703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__buf_2 fanout704 (.A(net705),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_2 fanout705 (.A(net707),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_4 fanout706 (.A(net707),
    .X(net706));
 sky130_fd_sc_hd__buf_2 fanout707 (.A(_03139_),
    .X(net707));
 sky130_fd_sc_hd__buf_2 fanout708 (.A(net709),
    .X(net708));
 sky130_fd_sc_hd__buf_2 fanout709 (.A(_02501_),
    .X(net709));
 sky130_fd_sc_hd__buf_2 fanout710 (.A(_02501_),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_4 fanout711 (.A(_02083_),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 fanout712 (.A(_02083_),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_4 fanout713 (.A(_02083_),
    .X(net713));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout714 (.A(_02083_),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_2 fanout715 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_2 fanout716 (.A(_06674_),
    .X(net716));
 sky130_fd_sc_hd__buf_2 fanout717 (.A(net718),
    .X(net717));
 sky130_fd_sc_hd__buf_2 fanout718 (.A(net720),
    .X(net718));
 sky130_fd_sc_hd__buf_2 fanout719 (.A(net720),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_2 fanout720 (.A(_06673_),
    .X(net720));
 sky130_fd_sc_hd__buf_2 fanout721 (.A(net723),
    .X(net721));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout722 (.A(net723),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_4 fanout723 (.A(_06409_),
    .X(net723));
 sky130_fd_sc_hd__buf_2 fanout724 (.A(net725),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_2 fanout725 (.A(_06409_),
    .X(net725));
 sky130_fd_sc_hd__buf_2 fanout726 (.A(_06409_),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_4 fanout727 (.A(net728),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_2 fanout728 (.A(_06244_),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_4 fanout729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_8 fanout730 (.A(_06244_),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_1 wire731 (.A(_06219_),
    .X(net731));
 sky130_fd_sc_hd__buf_1 max_cap732 (.A(_06182_),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_2 fanout733 (.A(net735),
    .X(net733));
 sky130_fd_sc_hd__buf_1 fanout734 (.A(net735),
    .X(net734));
 sky130_fd_sc_hd__buf_2 fanout735 (.A(_06164_),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_4 fanout736 (.A(net738),
    .X(net736));
 sky130_fd_sc_hd__buf_2 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 fanout738 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout739 (.A(net742),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_4 fanout740 (.A(net742),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 fanout741 (.A(net742),
    .X(net741));
 sky130_fd_sc_hd__buf_6 fanout742 (.A(_06164_),
    .X(net742));
 sky130_fd_sc_hd__buf_2 fanout743 (.A(net744),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 fanout744 (.A(net745),
    .X(net744));
 sky130_fd_sc_hd__buf_2 fanout745 (.A(_06163_),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 fanout746 (.A(net747),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_2 fanout747 (.A(_06163_),
    .X(net747));
 sky130_fd_sc_hd__buf_2 fanout748 (.A(net749),
    .X(net748));
 sky130_fd_sc_hd__buf_2 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__buf_2 fanout750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__buf_2 fanout751 (.A(_05120_),
    .X(net751));
 sky130_fd_sc_hd__buf_2 fanout752 (.A(net754),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_2 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__buf_2 fanout754 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_4 fanout755 (.A(net757),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(net757),
    .X(net756));
 sky130_fd_sc_hd__buf_2 fanout757 (.A(_04885_),
    .X(net757));
 sky130_fd_sc_hd__buf_2 fanout758 (.A(_04884_),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_2 fanout759 (.A(_04884_),
    .X(net759));
 sky130_fd_sc_hd__buf_2 fanout760 (.A(_04884_),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_1 max_cap761 (.A(_03883_),
    .X(net761));
 sky130_fd_sc_hd__buf_2 fanout762 (.A(_03877_),
    .X(net762));
 sky130_fd_sc_hd__buf_1 fanout763 (.A(_03877_),
    .X(net763));
 sky130_fd_sc_hd__buf_2 fanout764 (.A(_03877_),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_2 fanout765 (.A(_03877_),
    .X(net765));
 sky130_fd_sc_hd__buf_4 fanout766 (.A(_03747_),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_4 fanout767 (.A(_03747_),
    .X(net767));
 sky130_fd_sc_hd__buf_4 fanout768 (.A(_03747_),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 fanout769 (.A(_03747_),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_4 fanout770 (.A(net771),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_4 fanout771 (.A(_03464_),
    .X(net771));
 sky130_fd_sc_hd__buf_4 fanout772 (.A(_03170_),
    .X(net772));
 sky130_fd_sc_hd__buf_4 fanout773 (.A(_03170_),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_8 fanout774 (.A(_03170_),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_4 fanout775 (.A(_03170_),
    .X(net775));
 sky130_fd_sc_hd__buf_4 fanout776 (.A(net778),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_2 fanout777 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(_03169_),
    .X(net778));
 sky130_fd_sc_hd__buf_4 fanout779 (.A(net782),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_4 fanout780 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_4 fanout781 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__buf_2 fanout782 (.A(_03152_),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_4 fanout783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_4 fanout784 (.A(_03152_),
    .X(net784));
 sky130_fd_sc_hd__buf_4 fanout785 (.A(_03152_),
    .X(net785));
 sky130_fd_sc_hd__buf_2 fanout786 (.A(_03152_),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 fanout787 (.A(net788),
    .X(net787));
 sky130_fd_sc_hd__buf_4 fanout788 (.A(net791),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_4 fanout789 (.A(net791),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_2 fanout790 (.A(net791),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 fanout791 (.A(net795),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_4 fanout792 (.A(net795),
    .X(net792));
 sky130_fd_sc_hd__buf_2 fanout793 (.A(net795),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_4 fanout794 (.A(net795),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_4 fanout795 (.A(_03151_),
    .X(net795));
 sky130_fd_sc_hd__buf_4 fanout796 (.A(net803),
    .X(net796));
 sky130_fd_sc_hd__buf_2 fanout797 (.A(net803),
    .X(net797));
 sky130_fd_sc_hd__buf_4 fanout798 (.A(net803),
    .X(net798));
 sky130_fd_sc_hd__buf_2 fanout799 (.A(net803),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 fanout800 (.A(net802),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 fanout801 (.A(net802),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_4 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_2 fanout803 (.A(_03143_),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_4 fanout804 (.A(net806),
    .X(net804));
 sky130_fd_sc_hd__buf_4 fanout805 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__buf_2 fanout806 (.A(_03143_),
    .X(net806));
 sky130_fd_sc_hd__buf_4 fanout807 (.A(_03143_),
    .X(net807));
 sky130_fd_sc_hd__buf_2 fanout808 (.A(_03143_),
    .X(net808));
 sky130_fd_sc_hd__buf_4 fanout809 (.A(net812),
    .X(net809));
 sky130_fd_sc_hd__buf_4 fanout810 (.A(net812),
    .X(net810));
 sky130_fd_sc_hd__buf_2 fanout811 (.A(net812),
    .X(net811));
 sky130_fd_sc_hd__buf_2 fanout812 (.A(net821),
    .X(net812));
 sky130_fd_sc_hd__buf_4 fanout813 (.A(net815),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_4 fanout814 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__buf_4 fanout815 (.A(net821),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_4 fanout816 (.A(net818),
    .X(net816));
 sky130_fd_sc_hd__buf_4 fanout817 (.A(net818),
    .X(net817));
 sky130_fd_sc_hd__buf_2 fanout818 (.A(net821),
    .X(net818));
 sky130_fd_sc_hd__buf_4 fanout819 (.A(net821),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_4 fanout820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__buf_2 fanout821 (.A(_03142_),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 fanout822 (.A(net823),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_4 fanout823 (.A(net826),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 fanout824 (.A(net825),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_4 fanout825 (.A(net826),
    .X(net825));
 sky130_fd_sc_hd__buf_2 fanout826 (.A(_03137_),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_4 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_4 fanout828 (.A(net830),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_4 fanout829 (.A(net830),
    .X(net829));
 sky130_fd_sc_hd__buf_2 fanout830 (.A(_03137_),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_4 fanout831 (.A(net834),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_4 fanout832 (.A(net833),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_4 fanout833 (.A(net834),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_2 fanout834 (.A(_03137_),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_4 fanout835 (.A(net837),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_4 fanout836 (.A(net837),
    .X(net836));
 sky130_fd_sc_hd__buf_2 fanout837 (.A(_03137_),
    .X(net837));
 sky130_fd_sc_hd__buf_4 fanout838 (.A(net839),
    .X(net838));
 sky130_fd_sc_hd__buf_4 fanout839 (.A(_03136_),
    .X(net839));
 sky130_fd_sc_hd__buf_2 fanout840 (.A(_03136_),
    .X(net840));
 sky130_fd_sc_hd__buf_2 fanout841 (.A(net842),
    .X(net841));
 sky130_fd_sc_hd__buf_2 fanout842 (.A(_02702_),
    .X(net842));
 sky130_fd_sc_hd__buf_2 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_2 fanout844 (.A(_02702_),
    .X(net844));
 sky130_fd_sc_hd__buf_2 fanout845 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__clkbuf_4 fanout846 (.A(net852),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_4 fanout847 (.A(net852),
    .X(net847));
 sky130_fd_sc_hd__buf_2 fanout848 (.A(net852),
    .X(net848));
 sky130_fd_sc_hd__buf_2 fanout849 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_4 fanout850 (.A(net851),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_4 fanout851 (.A(net852),
    .X(net851));
 sky130_fd_sc_hd__buf_2 fanout852 (.A(_02468_),
    .X(net852));
 sky130_fd_sc_hd__buf_2 fanout853 (.A(net854),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 fanout854 (.A(net855),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_4 fanout855 (.A(_05134_),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 fanout856 (.A(net859),
    .X(net856));
 sky130_fd_sc_hd__buf_2 fanout857 (.A(net858),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_2 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_2 fanout859 (.A(_05134_),
    .X(net859));
 sky130_fd_sc_hd__buf_4 fanout860 (.A(_05133_),
    .X(net860));
 sky130_fd_sc_hd__buf_2 fanout861 (.A(net862),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_4 fanout862 (.A(net865),
    .X(net862));
 sky130_fd_sc_hd__buf_2 fanout863 (.A(net865),
    .X(net863));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout864 (.A(net865),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_4 fanout865 (.A(net866),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_4 fanout866 (.A(_05083_),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_4 fanout867 (.A(net869),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_4 fanout868 (.A(net869),
    .X(net868));
 sky130_fd_sc_hd__buf_2 fanout869 (.A(_05082_),
    .X(net869));
 sky130_fd_sc_hd__buf_2 fanout870 (.A(net871),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_2 fanout871 (.A(net872),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_2 fanout872 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 fanout873 (.A(net874),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_4 fanout874 (.A(_05082_),
    .X(net874));
 sky130_fd_sc_hd__buf_2 fanout875 (.A(net876),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_4 fanout876 (.A(net882),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_4 fanout877 (.A(net882),
    .X(net877));
 sky130_fd_sc_hd__buf_2 fanout878 (.A(net882),
    .X(net878));
 sky130_fd_sc_hd__buf_2 fanout879 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_2 fanout880 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_4 fanout881 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__buf_2 fanout882 (.A(_04421_),
    .X(net882));
 sky130_fd_sc_hd__buf_2 fanout883 (.A(net898),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_2 fanout884 (.A(net898),
    .X(net884));
 sky130_fd_sc_hd__buf_2 fanout885 (.A(net891),
    .X(net885));
 sky130_fd_sc_hd__buf_2 fanout886 (.A(net891),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_2 fanout887 (.A(net891),
    .X(net887));
 sky130_fd_sc_hd__buf_2 fanout888 (.A(net890),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_2 fanout889 (.A(net890),
    .X(net889));
 sky130_fd_sc_hd__buf_2 fanout890 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout891 (.A(net898),
    .X(net891));
 sky130_fd_sc_hd__buf_2 fanout892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_2 fanout893 (.A(net898),
    .X(net893));
 sky130_fd_sc_hd__buf_2 fanout894 (.A(net896),
    .X(net894));
 sky130_fd_sc_hd__buf_2 fanout895 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_4 fanout897 (.A(net898),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_2 fanout898 (.A(_03879_),
    .X(net898));
 sky130_fd_sc_hd__buf_2 fanout899 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__buf_2 fanout900 (.A(net903),
    .X(net900));
 sky130_fd_sc_hd__buf_2 fanout901 (.A(net902),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_2 fanout902 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_2 fanout903 (.A(_03879_),
    .X(net903));
 sky130_fd_sc_hd__buf_2 fanout904 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_2 fanout905 (.A(_03879_),
    .X(net905));
 sky130_fd_sc_hd__buf_2 fanout906 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__buf_2 fanout907 (.A(net910),
    .X(net907));
 sky130_fd_sc_hd__buf_2 fanout908 (.A(net910),
    .X(net908));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout910 (.A(_03879_),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_4 fanout911 (.A(net913),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_2 fanout912 (.A(net913),
    .X(net912));
 sky130_fd_sc_hd__buf_2 fanout913 (.A(_03875_),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_4 fanout914 (.A(net919),
    .X(net914));
 sky130_fd_sc_hd__buf_2 fanout915 (.A(net919),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_4 fanout916 (.A(net919),
    .X(net916));
 sky130_fd_sc_hd__buf_2 fanout917 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__buf_2 fanout918 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__buf_2 fanout919 (.A(_03874_),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_4 fanout920 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_4 fanout921 (.A(net927),
    .X(net921));
 sky130_fd_sc_hd__buf_4 fanout922 (.A(net927),
    .X(net922));
 sky130_fd_sc_hd__buf_2 fanout923 (.A(net927),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_4 fanout924 (.A(net925),
    .X(net924));
 sky130_fd_sc_hd__buf_2 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_4 fanout926 (.A(net927),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_4 fanout927 (.A(_03708_),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout928 (.A(_03463_),
    .X(net928));
 sky130_fd_sc_hd__buf_2 fanout929 (.A(_03463_),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_4 fanout930 (.A(_03462_),
    .X(net930));
 sky130_fd_sc_hd__buf_2 fanout931 (.A(_03462_),
    .X(net931));
 sky130_fd_sc_hd__buf_2 fanout932 (.A(net933),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_2 fanout933 (.A(_03460_),
    .X(net933));
 sky130_fd_sc_hd__buf_2 fanout934 (.A(_03459_),
    .X(net934));
 sky130_fd_sc_hd__buf_2 fanout935 (.A(_03459_),
    .X(net935));
 sky130_fd_sc_hd__buf_2 fanout936 (.A(_02910_),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_2 fanout937 (.A(_02910_),
    .X(net937));
 sky130_fd_sc_hd__buf_2 fanout938 (.A(net939),
    .X(net938));
 sky130_fd_sc_hd__buf_2 fanout939 (.A(_02693_),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 fanout940 (.A(_02693_),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_2 fanout941 (.A(_02693_),
    .X(net941));
 sky130_fd_sc_hd__buf_4 fanout942 (.A(_02690_),
    .X(net942));
 sky130_fd_sc_hd__buf_4 fanout943 (.A(_00015_),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_4 fanout944 (.A(_00015_),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout945 (.A(_00015_),
    .X(net945));
 sky130_fd_sc_hd__clkbuf_2 fanout946 (.A(_00015_),
    .X(net946));
 sky130_fd_sc_hd__buf_2 fanout947 (.A(net948),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_4 fanout948 (.A(net949),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 fanout949 (.A(_02509_),
    .X(net949));
 sky130_fd_sc_hd__buf_2 fanout950 (.A(net952),
    .X(net950));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout951 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout952 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 fanout953 (.A(_02508_),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_4 fanout954 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_4 fanout955 (.A(net957),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_4 fanout956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout957 (.A(_02500_),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout958 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__buf_4 fanout959 (.A(_02463_),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 fanout960 (.A(_02462_),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_4 fanout961 (.A(_02462_),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout962 (.A(net965),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_2 fanout963 (.A(net965),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout964 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_2 fanout965 (.A(_02449_),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_4 fanout966 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__buf_4 fanout967 (.A(_02433_),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_4 fanout968 (.A(_02432_),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_2 fanout969 (.A(_02432_),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 fanout970 (.A(_02428_),
    .X(net970));
 sky130_fd_sc_hd__buf_2 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout972 (.A(net975),
    .X(net972));
 sky130_fd_sc_hd__buf_2 fanout973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_2 fanout974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__buf_2 fanout975 (.A(_02421_),
    .X(net975));
 sky130_fd_sc_hd__buf_2 fanout976 (.A(net979),
    .X(net976));
 sky130_fd_sc_hd__buf_2 fanout977 (.A(net979),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_4 fanout978 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_2 fanout979 (.A(_02420_),
    .X(net979));
 sky130_fd_sc_hd__buf_4 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__buf_4 fanout981 (.A(net983),
    .X(net981));
 sky130_fd_sc_hd__buf_4 fanout982 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout983 (.A(_02416_),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_4 fanout984 (.A(_02381_),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_4 fanout985 (.A(_02381_),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout986 (.A(_02379_),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_2 fanout987 (.A(_02379_),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_4 fanout988 (.A(net990),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_2 fanout989 (.A(net990),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_4 fanout990 (.A(_02364_),
    .X(net990));
 sky130_fd_sc_hd__buf_4 fanout991 (.A(_02363_),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_4 fanout992 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout993 (.A(net226),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_4 fanout994 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__buf_4 fanout995 (.A(net224),
    .X(net995));
 sky130_fd_sc_hd__buf_4 fanout996 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__buf_4 fanout997 (.A(net223),
    .X(net997));
 sky130_fd_sc_hd__buf_2 fanout998 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_4 fanout999 (.A(net222),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_4 fanout1000 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 fanout1001 (.A(net221),
    .X(net1001));
 sky130_fd_sc_hd__buf_2 fanout1002 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__buf_4 fanout1003 (.A(net220),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 fanout1004 (.A(net1005),
    .X(net1004));
 sky130_fd_sc_hd__buf_4 fanout1005 (.A(net219),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_8 fanout1006 (.A(net218),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_4 fanout1007 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout1008 (.A(net217),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_8 fanout1009 (.A(net216),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_4 fanout1010 (.A(net1011),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_4 fanout1011 (.A(net215),
    .X(net1011));
 sky130_fd_sc_hd__buf_4 fanout1012 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout1013 (.A(net213),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout1014 (.A(net1015),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout1015 (.A(net212),
    .X(net1015));
 sky130_fd_sc_hd__buf_4 fanout1016 (.A(net211),
    .X(net1016));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1017 (.A(net211),
    .X(net1017));
 sky130_fd_sc_hd__buf_4 fanout1018 (.A(net1019),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 fanout1019 (.A(net210),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_4 fanout1020 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout1021 (.A(net209),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_4 fanout1022 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout1023 (.A(net208),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_4 fanout1024 (.A(net1025),
    .X(net1024));
 sky130_fd_sc_hd__buf_2 fanout1025 (.A(net207),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout1026 (.A(net1027),
    .X(net1026));
 sky130_fd_sc_hd__buf_2 fanout1027 (.A(net206),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout1028 (.A(net205),
    .X(net1028));
 sky130_fd_sc_hd__buf_2 fanout1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_2 fanout1030 (.A(net204),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_4 fanout1031 (.A(net1032),
    .X(net1031));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1032 (.A(net234),
    .X(net1032));
 sky130_fd_sc_hd__buf_2 fanout1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__buf_2 fanout1034 (.A(net233),
    .X(net1034));
 sky130_fd_sc_hd__buf_2 fanout1035 (.A(net1037),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_2 fanout1036 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__buf_2 fanout1037 (.A(net232),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_4 fanout1038 (.A(net231),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_2 fanout1039 (.A(net231),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_4 fanout1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__buf_2 fanout1041 (.A(net230),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_4 fanout1042 (.A(net229),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_2 fanout1043 (.A(net229),
    .X(net1043));
 sky130_fd_sc_hd__buf_2 fanout1044 (.A(net228),
    .X(net1044));
 sky130_fd_sc_hd__buf_2 fanout1045 (.A(net225),
    .X(net1045));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1046 (.A(net225),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_4 fanout1047 (.A(net1049),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_4 fanout1048 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__buf_2 fanout1049 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_4 fanout1050 (.A(net214),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_4 fanout1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_4 fanout1052 (.A(net1053),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_4 fanout1053 (.A(net203),
    .X(net1053));
 sky130_fd_sc_hd__buf_4 fanout1054 (.A(\mem_wordsize[2] ),
    .X(net1054));
 sky130_fd_sc_hd__clkbuf_2 fanout1055 (.A(\mem_wordsize[2] ),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_4 fanout1056 (.A(net1058),
    .X(net1056));
 sky130_fd_sc_hd__buf_2 fanout1057 (.A(net1059),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_2 fanout1058 (.A(net1059),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 fanout1059 (.A(\mem_wordsize[1] ),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 fanout1060 (.A(net1062),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_2 fanout1061 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_4 fanout1062 (.A(\cpu_state[7] ),
    .X(net1062));
 sky130_fd_sc_hd__buf_2 fanout1063 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_2 fanout1064 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_4 fanout1065 (.A(net1070),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_4 fanout1066 (.A(net1070),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_2 fanout1067 (.A(net1070),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_4 fanout1068 (.A(net1070),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_2 fanout1069 (.A(net1070),
    .X(net1069));
 sky130_fd_sc_hd__clkbuf_4 fanout1070 (.A(\cpu_state[5] ),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_4 fanout1071 (.A(net1074),
    .X(net1071));
 sky130_fd_sc_hd__buf_2 fanout1072 (.A(net1073),
    .X(net1072));
 sky130_fd_sc_hd__clkbuf_4 fanout1073 (.A(net1074),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_4 fanout1074 (.A(\cpu_state[4] ),
    .X(net1074));
 sky130_fd_sc_hd__buf_2 fanout1075 (.A(\cpu_state[3] ),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sky130_fd_sc_hd__buf_2 fanout1077 (.A(net1079),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_4 fanout1078 (.A(net1079),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_4 fanout1079 (.A(\cpu_state[3] ),
    .X(net1079));
 sky130_fd_sc_hd__buf_2 fanout1080 (.A(net1081),
    .X(net1080));
 sky130_fd_sc_hd__buf_2 fanout1081 (.A(net1087),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_4 fanout1082 (.A(net1086),
    .X(net1082));
 sky130_fd_sc_hd__buf_2 fanout1083 (.A(net1084),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__buf_2 fanout1085 (.A(net1086),
    .X(net1085));
 sky130_fd_sc_hd__buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__clkbuf_2 fanout1087 (.A(\cpu_state[3] ),
    .X(net1087));
 sky130_fd_sc_hd__buf_2 fanout1088 (.A(\cpu_state[2] ),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_4 fanout1089 (.A(\cpu_state[1] ),
    .X(net1089));
 sky130_fd_sc_hd__buf_2 fanout1090 (.A(net1093),
    .X(net1090));
 sky130_fd_sc_hd__buf_2 fanout1091 (.A(net1093),
    .X(net1091));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1092 (.A(net1093),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_2 fanout1093 (.A(net1109),
    .X(net1093));
 sky130_fd_sc_hd__buf_2 fanout1094 (.A(net1109),
    .X(net1094));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1095 (.A(net1109),
    .X(net1095));
 sky130_fd_sc_hd__buf_2 fanout1096 (.A(net1100),
    .X(net1096));
 sky130_fd_sc_hd__buf_1 fanout1097 (.A(net1100),
    .X(net1097));
 sky130_fd_sc_hd__buf_2 fanout1098 (.A(net1100),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_2 fanout1100 (.A(net1109),
    .X(net1100));
 sky130_fd_sc_hd__buf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sky130_fd_sc_hd__buf_2 fanout1102 (.A(net1104),
    .X(net1102));
 sky130_fd_sc_hd__buf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_2 fanout1104 (.A(net1109),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 fanout1105 (.A(net1108),
    .X(net1105));
 sky130_fd_sc_hd__clkbuf_2 fanout1106 (.A(net1107),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sky130_fd_sc_hd__clkbuf_2 fanout1108 (.A(net1109),
    .X(net1108));
 sky130_fd_sc_hd__buf_2 fanout1109 (.A(\genblk1.genblk1.pcpi_mul.rs1[0] ),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_4 fanout1110 (.A(net1111),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_4 fanout1111 (.A(\genblk2.pcpi_div.pcpi_ready ),
    .X(net1111));
 sky130_fd_sc_hd__buf_4 fanout1112 (.A(\genblk2.pcpi_div.pcpi_ready ),
    .X(net1112));
 sky130_fd_sc_hd__buf_2 fanout1113 (.A(\genblk2.pcpi_div.pcpi_ready ),
    .X(net1113));
 sky130_fd_sc_hd__buf_2 fanout1114 (.A(net1116),
    .X(net1114));
 sky130_fd_sc_hd__buf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sky130_fd_sc_hd__buf_1 fanout1116 (.A(net1117),
    .X(net1116));
 sky130_fd_sc_hd__buf_2 fanout1117 (.A(net1124),
    .X(net1117));
 sky130_fd_sc_hd__buf_2 fanout1118 (.A(net1120),
    .X(net1118));
 sky130_fd_sc_hd__clkbuf_2 fanout1119 (.A(net1120),
    .X(net1119));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1120 (.A(net1124),
    .X(net1120));
 sky130_fd_sc_hd__buf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sky130_fd_sc_hd__buf_2 fanout1122 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__buf_2 fanout1123 (.A(net1124),
    .X(net1123));
 sky130_fd_sc_hd__clkbuf_2 fanout1124 (.A(net1125),
    .X(net1124));
 sky130_fd_sc_hd__clkbuf_4 fanout1125 (.A(net1126),
    .X(net1125));
 sky130_fd_sc_hd__buf_2 fanout1126 (.A(\genblk2.pcpi_div.outsign ),
    .X(net1126));
 sky130_fd_sc_hd__buf_2 fanout1127 (.A(net1128),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_2 fanout1128 (.A(\decoded_imm_j[20] ),
    .X(net1128));
 sky130_fd_sc_hd__clkbuf_4 fanout1129 (.A(\decoded_imm_j[20] ),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_4 fanout1130 (.A(net1132),
    .X(net1130));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1131 (.A(net1132),
    .X(net1131));
 sky130_fd_sc_hd__clkbuf_2 fanout1132 (.A(instr_rdinstrh),
    .X(net1132));
 sky130_fd_sc_hd__buf_2 fanout1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__buf_2 fanout1134 (.A(instr_rdinstrh),
    .X(net1134));
 sky130_fd_sc_hd__buf_2 fanout1135 (.A(net1136),
    .X(net1135));
 sky130_fd_sc_hd__buf_2 fanout1136 (.A(instr_rdinstr),
    .X(net1136));
 sky130_fd_sc_hd__buf_2 fanout1137 (.A(net1138),
    .X(net1137));
 sky130_fd_sc_hd__clkbuf_2 fanout1138 (.A(instr_rdinstr),
    .X(net1138));
 sky130_fd_sc_hd__buf_2 fanout1139 (.A(net1140),
    .X(net1139));
 sky130_fd_sc_hd__buf_2 fanout1140 (.A(instr_rdcycleh),
    .X(net1140));
 sky130_fd_sc_hd__buf_2 fanout1141 (.A(net1142),
    .X(net1141));
 sky130_fd_sc_hd__clkbuf_2 fanout1142 (.A(instr_rdcycleh),
    .X(net1142));
 sky130_fd_sc_hd__clkbuf_4 fanout1143 (.A(net1145),
    .X(net1143));
 sky130_fd_sc_hd__clkbuf_2 fanout1144 (.A(net1145),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_4 fanout1145 (.A(instr_sub),
    .X(net1145));
 sky130_fd_sc_hd__buf_2 fanout1146 (.A(net1147),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_2 fanout1147 (.A(net1148),
    .X(net1147));
 sky130_fd_sc_hd__clkbuf_2 fanout1148 (.A(net1149),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_4 fanout1149 (.A(instr_jal),
    .X(net1149));
 sky130_fd_sc_hd__buf_2 fanout1150 (.A(net1152),
    .X(net1150));
 sky130_fd_sc_hd__buf_1 fanout1151 (.A(net1152),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_4 fanout1152 (.A(instr_jal),
    .X(net1152));
 sky130_fd_sc_hd__buf_4 fanout1153 (.A(net1156),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_4 fanout1154 (.A(net1156),
    .X(net1154));
 sky130_fd_sc_hd__buf_4 fanout1155 (.A(net1156),
    .X(net1155));
 sky130_fd_sc_hd__clkbuf_4 fanout1156 (.A(latched_stalu),
    .X(net1156));
 sky130_fd_sc_hd__clkbuf_4 fanout1157 (.A(net259),
    .X(net1157));
 sky130_fd_sc_hd__buf_4 fanout1158 (.A(net249),
    .X(net1158));
 sky130_fd_sc_hd__buf_4 fanout1159 (.A(net245),
    .X(net1159));
 sky130_fd_sc_hd__clkbuf_4 fanout1160 (.A(net243),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_4 fanout1161 (.A(net242),
    .X(net1161));
 sky130_fd_sc_hd__buf_4 fanout1162 (.A(net241),
    .X(net1162));
 sky130_fd_sc_hd__buf_4 fanout1163 (.A(net239),
    .X(net1163));
 sky130_fd_sc_hd__buf_4 fanout1164 (.A(net238),
    .X(net1164));
 sky130_fd_sc_hd__clkbuf_4 fanout1165 (.A(net237),
    .X(net1165));
 sky130_fd_sc_hd__clkbuf_4 fanout1166 (.A(net236),
    .X(net1166));
 sky130_fd_sc_hd__clkbuf_4 fanout1167 (.A(net266),
    .X(net1167));
 sky130_fd_sc_hd__buf_4 fanout1168 (.A(net265),
    .X(net1168));
 sky130_fd_sc_hd__buf_4 fanout1169 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_4 fanout1170 (.A(net126),
    .X(net1170));
 sky130_fd_sc_hd__buf_4 fanout1171 (.A(net125),
    .X(net1171));
 sky130_fd_sc_hd__clkbuf_4 fanout1172 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__buf_4 fanout1173 (.A(net124),
    .X(net1173));
 sky130_fd_sc_hd__buf_4 fanout1174 (.A(net1175),
    .X(net1174));
 sky130_fd_sc_hd__buf_4 fanout1175 (.A(net123),
    .X(net1175));
 sky130_fd_sc_hd__clkbuf_8 fanout1176 (.A(net122),
    .X(net1176));
 sky130_fd_sc_hd__buf_4 fanout1177 (.A(net119),
    .X(net1177));
 sky130_fd_sc_hd__buf_4 fanout1178 (.A(net1179),
    .X(net1178));
 sky130_fd_sc_hd__buf_4 fanout1179 (.A(net108),
    .X(net1179));
 sky130_fd_sc_hd__buf_4 fanout1180 (.A(net97),
    .X(net1180));
 sky130_fd_sc_hd__buf_4 fanout1181 (.A(net97),
    .X(net1181));
 sky130_fd_sc_hd__clkbuf_4 fanout1182 (.A(net1187),
    .X(net1182));
 sky130_fd_sc_hd__clkbuf_4 fanout1183 (.A(net1187),
    .X(net1183));
 sky130_fd_sc_hd__buf_4 fanout1184 (.A(net1186),
    .X(net1184));
 sky130_fd_sc_hd__clkbuf_4 fanout1185 (.A(net1186),
    .X(net1185));
 sky130_fd_sc_hd__buf_2 fanout1186 (.A(net1187),
    .X(net1186));
 sky130_fd_sc_hd__clkbuf_4 fanout1187 (.A(decoder_trigger),
    .X(net1187));
 sky130_fd_sc_hd__clkbuf_4 fanout1188 (.A(net1189),
    .X(net1188));
 sky130_fd_sc_hd__buf_4 fanout1189 (.A(net227),
    .X(net1189));
 sky130_fd_sc_hd__buf_2 fanout1190 (.A(net1191),
    .X(net1190));
 sky130_fd_sc_hd__buf_2 fanout1191 (.A(net1205),
    .X(net1191));
 sky130_fd_sc_hd__buf_2 fanout1192 (.A(net1198),
    .X(net1192));
 sky130_fd_sc_hd__buf_2 fanout1193 (.A(net1197),
    .X(net1193));
 sky130_fd_sc_hd__buf_2 fanout1194 (.A(net1197),
    .X(net1194));
 sky130_fd_sc_hd__buf_2 fanout1195 (.A(net1196),
    .X(net1195));
 sky130_fd_sc_hd__buf_2 fanout1196 (.A(net1197),
    .X(net1196));
 sky130_fd_sc_hd__buf_2 fanout1197 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_2 fanout1198 (.A(net1205),
    .X(net1198));
 sky130_fd_sc_hd__buf_2 fanout1199 (.A(net1204),
    .X(net1199));
 sky130_fd_sc_hd__buf_2 fanout1200 (.A(net1204),
    .X(net1200));
 sky130_fd_sc_hd__clkbuf_2 fanout1201 (.A(net1204),
    .X(net1201));
 sky130_fd_sc_hd__buf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sky130_fd_sc_hd__buf_2 fanout1203 (.A(net1204),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_2 fanout1204 (.A(net1205),
    .X(net1204));
 sky130_fd_sc_hd__buf_2 fanout1205 (.A(_02378_),
    .X(net1205));
 sky130_fd_sc_hd__clkbuf_4 fanout1206 (.A(net1207),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_2 fanout1207 (.A(_02378_),
    .X(net1207));
 sky130_fd_sc_hd__clkbuf_4 fanout1208 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__buf_2 fanout1209 (.A(_02378_),
    .X(net1209));
 sky130_fd_sc_hd__buf_2 fanout1210 (.A(net1222),
    .X(net1210));
 sky130_fd_sc_hd__clkbuf_2 fanout1211 (.A(net1222),
    .X(net1211));
 sky130_fd_sc_hd__buf_2 fanout1212 (.A(net1214),
    .X(net1212));
 sky130_fd_sc_hd__clkbuf_2 fanout1213 (.A(net1222),
    .X(net1213));
 sky130_fd_sc_hd__clkbuf_4 fanout1214 (.A(net1222),
    .X(net1214));
 sky130_fd_sc_hd__buf_2 fanout1215 (.A(net1216),
    .X(net1215));
 sky130_fd_sc_hd__buf_2 fanout1216 (.A(net1222),
    .X(net1216));
 sky130_fd_sc_hd__buf_2 fanout1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__clkbuf_2 fanout1218 (.A(net1222),
    .X(net1218));
 sky130_fd_sc_hd__buf_2 fanout1219 (.A(net1221),
    .X(net1219));
 sky130_fd_sc_hd__buf_2 fanout1220 (.A(net1221),
    .X(net1220));
 sky130_fd_sc_hd__clkbuf_2 fanout1221 (.A(net1222),
    .X(net1221));
 sky130_fd_sc_hd__buf_2 fanout1222 (.A(_02378_),
    .X(net1222));
 sky130_fd_sc_hd__clkbuf_4 fanout1223 (.A(net34),
    .X(net1223));
 sky130_fd_sc_hd__clkbuf_2 fanout1224 (.A(net34),
    .X(net1224));
 sky130_fd_sc_hd__clkbuf_2 fanout1225 (.A(net1227),
    .X(net1225));
 sky130_fd_sc_hd__clkbuf_2 fanout1226 (.A(net1227),
    .X(net1226));
 sky130_fd_sc_hd__buf_2 fanout1227 (.A(net1241),
    .X(net1227));
 sky130_fd_sc_hd__clkbuf_2 fanout1228 (.A(net1230),
    .X(net1228));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1229 (.A(net1230),
    .X(net1229));
 sky130_fd_sc_hd__clkbuf_2 fanout1230 (.A(net1241),
    .X(net1230));
 sky130_fd_sc_hd__buf_2 fanout1231 (.A(net1241),
    .X(net1231));
 sky130_fd_sc_hd__buf_2 fanout1232 (.A(net1233),
    .X(net1232));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1233 (.A(net1234),
    .X(net1233));
 sky130_fd_sc_hd__clkbuf_2 fanout1234 (.A(net1241),
    .X(net1234));
 sky130_fd_sc_hd__buf_2 fanout1235 (.A(net1237),
    .X(net1235));
 sky130_fd_sc_hd__buf_1 fanout1236 (.A(net1237),
    .X(net1236));
 sky130_fd_sc_hd__buf_2 fanout1237 (.A(net1241),
    .X(net1237));
 sky130_fd_sc_hd__clkbuf_2 fanout1238 (.A(net1239),
    .X(net1238));
 sky130_fd_sc_hd__clkbuf_2 fanout1239 (.A(net1240),
    .X(net1239));
 sky130_fd_sc_hd__buf_1 fanout1240 (.A(net1241),
    .X(net1240));
 sky130_fd_sc_hd__buf_2 fanout1241 (.A(net34),
    .X(net1241));
 sky130_fd_sc_hd__conb_1 picorv32_1242 (.LO(net1242));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_66_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_67_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_75_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_76_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_77_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_78_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_79_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_80_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_81_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_82_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_83_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_84_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_85_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_86_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_87_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_88_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_89_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_90_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_91_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_92_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_93_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_94_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_95_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_96_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_97_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_98_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_99_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_100_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_101_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_102_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_103_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_104_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_105_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_106_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_107_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_108_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_109_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_110_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_111_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_112_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_113_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_114_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_115_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_116_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_117_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_118_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_119_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_120_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_121_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_122_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_123_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_124_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_125_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_126_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_127_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_128_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_129_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_130_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_131_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_132_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_133_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_134_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_135_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_136_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_137_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_138_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_139_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_140_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_141_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_142_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_143_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_144_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_145_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_146_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_147_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_148_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_149_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_150_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_151_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_152_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_153_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_154_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_155_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_156_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_157_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_158_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_159_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_160_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_161_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_162_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_163_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_164_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_165_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_166_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_167_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_169_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_170_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_171_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_172_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_173_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_174_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_175_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_176_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_177_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_178_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_179_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_180_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_181_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_182_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_183_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_184_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_185_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_186_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_187_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_188_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_189_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_190_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_191_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_192_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_193_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_194_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_195_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_196_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_197_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_198_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_199_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__inv_8 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_8 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__inv_16 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__inv_16 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_8 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__inv_12 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__inv_16 clkload10 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload11 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload12 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload15 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload16 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload17 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload18 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_4 clkload19 (.A(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkinv_4 clkload20 (.A(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload21 (.A(clknet_leaf_195_clk));
 sky130_fd_sc_hd__bufinv_16 clkload22 (.A(clknet_leaf_196_clk));
 sky130_fd_sc_hd__inv_6 clkload23 (.A(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkinv_2 clkload24 (.A(clknet_leaf_198_clk));
 sky130_fd_sc_hd__bufinv_16 clkload25 (.A(clknet_leaf_199_clk));
 sky130_fd_sc_hd__bufinv_16 clkload26 (.A(clknet_leaf_178_clk));
 sky130_fd_sc_hd__inv_6 clkload27 (.A(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload28 (.A(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload29 (.A(clknet_leaf_182_clk));
 sky130_fd_sc_hd__inv_8 clkload30 (.A(clknet_leaf_183_clk));
 sky130_fd_sc_hd__inv_6 clkload31 (.A(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_185_clk));
 sky130_fd_sc_hd__inv_8 clkload33 (.A(clknet_leaf_186_clk));
 sky130_fd_sc_hd__inv_6 clkload34 (.A(clknet_leaf_187_clk));
 sky130_fd_sc_hd__inv_8 clkload35 (.A(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkinv_8 clkload36 (.A(clknet_leaf_189_clk));
 sky130_fd_sc_hd__bufinv_16 clkload37 (.A(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkinv_2 clkload38 (.A(clknet_leaf_192_clk));
 sky130_fd_sc_hd__inv_6 clkload39 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload40 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkinv_2 clkload41 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__inv_8 clkload42 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_2 clkload43 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_2 clkload44 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__bufinv_16 clkload45 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkinv_4 clkload46 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload47 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_4 clkload48 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload49 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_2 clkload50 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload51 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload52 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload53 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload54 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload55 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__inv_6 clkload56 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__inv_8 clkload57 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__inv_6 clkload58 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinv_4 clkload59 (.A(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload60 (.A(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload61 (.A(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload62 (.A(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload63 (.A(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkinv_4 clkload64 (.A(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload65 (.A(clknet_leaf_166_clk));
 sky130_fd_sc_hd__bufinv_16 clkload66 (.A(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkinv_4 clkload67 (.A(clknet_leaf_169_clk));
 sky130_fd_sc_hd__inv_6 clkload68 (.A(clknet_leaf_172_clk));
 sky130_fd_sc_hd__inv_8 clkload69 (.A(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkinv_4 clkload70 (.A(clknet_leaf_152_clk));
 sky130_fd_sc_hd__inv_12 clkload71 (.A(clknet_leaf_154_clk));
 sky130_fd_sc_hd__inv_8 clkload72 (.A(clknet_leaf_155_clk));
 sky130_fd_sc_hd__inv_8 clkload73 (.A(clknet_leaf_156_clk));
 sky130_fd_sc_hd__inv_12 clkload74 (.A(clknet_leaf_157_clk));
 sky130_fd_sc_hd__inv_12 clkload75 (.A(clknet_leaf_158_clk));
 sky130_fd_sc_hd__inv_12 clkload76 (.A(clknet_leaf_159_clk));
 sky130_fd_sc_hd__inv_12 clkload77 (.A(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkinv_8 clkload78 (.A(clknet_leaf_161_clk));
 sky130_fd_sc_hd__bufinv_16 clkload79 (.A(clknet_leaf_162_clk));
 sky130_fd_sc_hd__bufinv_16 clkload80 (.A(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload81 (.A(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload82 (.A(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload83 (.A(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload84 (.A(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload85 (.A(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload86 (.A(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkinv_4 clkload87 (.A(clknet_leaf_138_clk));
 sky130_fd_sc_hd__inv_6 clkload88 (.A(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload89 (.A(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkinv_2 clkload90 (.A(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkinv_4 clkload91 (.A(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload92 (.A(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload93 (.A(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkinv_4 clkload94 (.A(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload95 (.A(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload96 (.A(clknet_leaf_147_clk));
 sky130_fd_sc_hd__bufinv_16 clkload97 (.A(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload98 (.A(clknet_leaf_150_clk));
 sky130_fd_sc_hd__inv_8 clkload99 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_4 clkload100 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_2 clkload101 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__inv_8 clkload102 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkinv_4 clkload103 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__inv_6 clkload104 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkinv_8 clkload105 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload106 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__bufinv_16 clkload107 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__inv_6 clkload108 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__inv_8 clkload109 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload110 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__inv_6 clkload111 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__inv_8 clkload112 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_4 clkload113 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__bufinv_16 clkload114 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload115 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__bufinv_16 clkload116 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload117 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkinv_4 clkload118 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload119 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload120 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload121 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__inv_8 clkload122 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkinv_4 clkload123 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__bufinv_16 clkload124 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__inv_6 clkload125 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinv_8 clkload126 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload127 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__inv_12 clkload128 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__inv_6 clkload129 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__inv_8 clkload130 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__inv_12 clkload131 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkinv_2 clkload132 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinv_4 clkload133 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload134 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__inv_6 clkload135 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__bufinv_16 clkload136 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__inv_12 clkload137 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload138 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__bufinv_16 clkload139 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload140 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__bufinv_16 clkload141 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinv_2 clkload142 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__bufinv_16 clkload143 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload144 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload145 (.A(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkinv_2 clkload146 (.A(clknet_leaf_129_clk));
 sky130_fd_sc_hd__inv_6 clkload147 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload148 (.A(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload149 (.A(clknet_leaf_132_clk));
 sky130_fd_sc_hd__inv_6 clkload150 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__inv_6 clkload151 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkinv_2 clkload152 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__inv_6 clkload153 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__inv_8 clkload154 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkinv_4 clkload155 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload156 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__inv_6 clkload157 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__bufinv_16 clkload158 (.A(clknet_leaf_118_clk));
 sky130_fd_sc_hd__inv_6 clkload159 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__inv_6 clkload160 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__inv_8 clkload161 (.A(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload162 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__inv_8 clkload163 (.A(clknet_leaf_123_clk));
 sky130_fd_sc_hd__inv_8 clkload164 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__inv_6 clkload165 (.A(clknet_leaf_125_clk));
 sky130_fd_sc_hd__inv_6 clkload166 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__bufinv_16 clkload167 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_4 clkload168 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__bufinv_16 clkload169 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkinv_4 clkload170 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload171 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload172 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__inv_8 clkload173 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload174 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload175 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkinv_4 clkload176 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__bufinv_16 clkload177 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkinv_2 clkload178 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkinv_8 clkload179 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload180 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__inv_6 clkload181 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkinv_4 clkload182 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload183 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__inv_6 clkload184 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkinv_4 clkload185 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload186 (.A(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload187 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\genblk1.genblk1.pcpi_mul.pcpi_wait ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\genblk1.genblk1.pcpi_mul.instr_mul ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\cpuregs[0][25] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\cpuregs[0][30] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\cpuregs[0][2] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\cpuregs[0][16] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\cpuregs[0][17] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\cpuregs[0][31] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\cpuregs[0][7] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\cpuregs[0][19] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\cpuregs[0][0] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[15] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_01385_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[22] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_01392_),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\reg_next_pc[1] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[14] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_01384_),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net62),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net64),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[10] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_01380_),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[18] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_01388_),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[4] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\cpuregs[26][12] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\cpuregs[26][25] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\cpuregs[26][20] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\cpuregs[14][29] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\cpuregs[30][12] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net63),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\cpuregs[30][18] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net36),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net61),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\cpuregs[24][7] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\cpuregs[24][13] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\cpuregs[24][11] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net38),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(instr_ecall_ebreak),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[7] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_01377_),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\cpuregs[28][25] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\cpuregs[24][9] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\cpuregs[28][24] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\cpuregs[28][4] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\cpuregs[22][2] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\cpuregs[20][5] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\cpuregs[26][9] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net39),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[6] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_01376_),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net59),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\cpuregs[12][10] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\cpuregs[24][17] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\cpuregs[24][10] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\genblk2.pcpi_div.instr_remu ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_00048_),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\cpuregs[26][5] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net50),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[9] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\cpuregs[12][27] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\cpuregs[26][3] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\cpuregs[26][4] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\cpuregs[28][23] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\cpuregs[24][14] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\cpuregs[24][2] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\cpuregs[30][24] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[27] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\cpuregs[26][15] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\cpuregs[28][29] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\cpuregs[22][20] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\cpuregs[20][4] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\cpuregs[26][2] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\cpuregs[26][17] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[24] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\cpuregs[24][20] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\cpuregs[26][18] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\cpuregs[22][14] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[0] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\cpuregs[28][5] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\cpuregs[20][22] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\cpuregs[12][29] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\cpuregs[30][0] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net145),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\cpuregs[14][2] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\cpuregs[24][22] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\cpuregs[24][21] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\cpuregs[28][1] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\cpuregs[26][29] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\cpuregs[20][2] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\decoded_rd[4] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\decoded_rd[2] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\cpuregs[14][28] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\cpuregs[30][28] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\cpuregs[12][11] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\cpuregs[24][25] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\cpuregs[26][6] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\cpuregs[12][25] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\cpuregs[14][4] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(instr_auipc),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\cpuregs[14][10] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\cpuregs[20][25] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\cpuregs[28][28] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\cpuregs[26][31] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net35),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\cpuregs[14][22] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\cpuregs[22][26] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\cpuregs[31][13] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\cpuregs[26][24] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[25] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\cpuregs[30][20] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net135),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\cpuregs[29][12] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\cpuregs[30][30] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\cpuregs[14][13] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\cpuregs[29][10] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\cpuregs[14][3] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\cpuregs[26][23] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\cpuregs[16][14] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\cpuregs[20][3] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\cpuregs[24][16] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[2] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net148),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\cpuregs[28][21] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net56),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\cpuregs[22][19] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\cpuregs[26][14] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\cpuregs[30][23] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\cpuregs[16][8] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\cpuregs[12][2] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\cpuregs[14][21] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\cpuregs[26][13] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net136),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\cpuregs[12][16] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\cpuregs[24][4] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[29] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\cpuregs[28][2] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\cpuregs[26][16] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\cpuregs[29][13] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\cpuregs[23][15] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\cpuregs[24][5] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\cpuregs[20][27] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\cpuregs[26][27] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\cpuregs[12][30] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net55),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[23] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net46),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net163),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\cpuregs[12][7] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net60),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\decoded_rd[1] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_00966_),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[1] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net146),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\cpuregs[22][9] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\cpuregs[13][3] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\cpuregs[20][18] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\cpuregs[12][8] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\cpuregs[14][27] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\cpuregs[31][2] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\cpuregs[21][15] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\cpuregs[12][14] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net37),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\cpuregs[24][6] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net159),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\cpuregs[30][13] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\cpuregs[22][22] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net139),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\cpuregs[15][11] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\cpuregs[12][1] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\cpuregs[15][4] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\cpuregs[28][14] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\cpuregs[26][28] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\cpuregs[8][13] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\cpuregs[12][3] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\cpuregs[22][1] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[2] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_01372_),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\cpuregs[12][18] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net42),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net165),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[30] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\cpuregs[30][6] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\cpuregs[20][30] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\cpuregs[12][13] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\cpuregs[23][21] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\cpuregs[21][7] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\cpuregs[21][20] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\cpuregs[24][3] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[29] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\cpuregs[24][12] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\cpuregs[12][23] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\cpuregs[20][7] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net141),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\cpuregs[31][21] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\cpuregs[30][25] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\cpuregs[29][21] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net144),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\cpuregs[22][29] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\cpuregs[20][17] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\cpuregs[13][18] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\cpuregs[4][26] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\cpuregs[23][4] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\cpuregs[30][15] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\cpuregs[15][13] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net150),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\cpuregs[14][15] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\cpuregs[26][7] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\cpuregs[31][24] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\cpuregs[12][5] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\cpuregs[23][16] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\cpuregs[13][2] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\cpuregs[30][31] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\cpuregs[22][16] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\cpuregs[22][8] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\cpuregs[24][8] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\cpuregs[8][18] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\cpuregs[30][3] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\cpuregs[15][10] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\cpuregs[20][10] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\cpuregs[12][0] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\cpuregs[29][5] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\cpuregs[28][0] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\cpuregs[20][23] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\cpuregs[29][0] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\cpuregs[13][8] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\cpuregs[30][21] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[9] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_01379_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\cpuregs[14][9] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\cpuregs[20][29] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net147),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\cpuregs[26][8] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\cpuregs[22][11] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\cpuregs[13][6] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[25] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\cpuregs[14][23] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\cpuregs[20][12] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\cpuregs[24][28] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\cpuregs[14][26] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\cpuregs[22][0] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(net53),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\cpuregs[28][12] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\cpuregs[16][2] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\cpuregs[14][31] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\cpuregs[14][25] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\cpuregs[10][18] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\cpuregs[28][26] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\cpuregs[30][11] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\cpuregs[31][10] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\cpuregs[28][13] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\cpuregs[13][11] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\cpuregs[30][19] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\cpuregs[21][10] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\cpuregs[24][26] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\cpuregs[2][24] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\cpuregs[26][26] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\cpuregs[20][0] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\cpuregs[23][18] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\cpuregs[13][15] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net162),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\cpuregs[14][18] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\cpuregs[23][14] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[27] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_01397_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\cpuregs[28][15] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\cpuregs[14][0] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[62] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\cpuregs[14][6] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\cpuregs[28][27] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net43),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\cpuregs[15][29] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\cpuregs[29][6] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\cpuregs[12][9] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net187),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\cpuregs[4][29] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\cpuregs[22][21] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\cpuregs[29][22] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net58),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\cpuregs[12][31] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\cpuregs[14][17] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net48),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\cpuregs[26][30] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\cpuregs[20][20] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\cpuregs[20][15] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\cpuregs[31][8] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\cpuregs[12][4] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\cpuregs[22][23] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\cpuregs[31][7] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\cpuregs[13][23] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\cpuregs[24][30] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\cpuregs[29][20] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\cpuregs[20][8] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\cpuregs[20][28] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\cpuregs[29][3] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\cpuregs[14][30] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\cpuregs[23][13] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\cpuregs[23][23] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\decoded_rd[3] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(net52),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\cpuregs[12][15] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\cpuregs[31][6] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\cpuregs[28][6] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\cpuregs[31][23] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\cpuregs[22][25] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\cpuregs[31][3] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\cpuregs[15][30] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\cpuregs[30][10] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net41),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\cpuregs[24][24] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\cpuregs[12][19] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[28] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\cpuregs[26][10] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\cpuregs[10][15] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[26] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\cpuregs[28][20] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\cpuregs[10][9] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\cpuregs[30][14] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[3] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\cpuregs[14][8] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(net166),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\cpuregs[26][1] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\cpuregs[22][6] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\cpuregs[30][29] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\cpuregs[10][10] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\cpuregs[13][4] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[26] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(net137),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\cpuregs[23][6] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(net149),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\cpuregs[26][21] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(net51),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\cpuregs[12][20] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\cpuregs[29][11] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(instr_bltu),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\cpuregs[21][5] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\cpuregs[23][3] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\cpuregs[31][11] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\cpuregs[21][21] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\cpuregs[29][27] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\cpuregs[28][18] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\cpuregs[31][15] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\cpuregs[15][7] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\cpuregs[22][4] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\cpuregs[24][31] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\cpuregs[22][24] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\cpuregs[16][3] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\cpuregs[8][28] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\cpuregs[27][14] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\cpuregs[12][17] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\cpuregs[8][21] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\cpuregs[20][24] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\cpuregs[22][15] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\cpuregs[21][8] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net152),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\cpuregs[12][6] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\cpuregs[13][17] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\cpuregs[30][27] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(net156),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\cpuregs[29][30] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\cpuregs[28][22] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[19] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\cpuregs[14][1] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\cpuregs[15][23] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\cpuregs[22][27] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\cpuregs[12][22] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(net40),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\cpuregs[10][14] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\cpuregs[31][12] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\cpuregs[25][12] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\cpuregs[8][8] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\cpuregs[16][26] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\cpuregs[31][18] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[5] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\cpuregs[22][12] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\cpuregs[15][21] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\cpuregs[23][12] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\cpuregs[28][11] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\cpuregs[14][20] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\cpuregs[14][16] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\cpuregs[30][9] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\cpuregs[27][2] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\cpuregs[29][15] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\cpuregs[10][21] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\cpuregs[8][2] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(net164),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\cpuregs[22][17] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\cpuregs[21][24] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\cpuregs[23][9] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\cpuregs[20][21] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\cpuregs[8][14] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\cpuregs[28][3] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\cpuregs[15][14] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\cpuregs[14][14] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\cpuregs[16][17] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\cpuregs[14][7] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\cpuregs[13][21] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\cpuregs[30][8] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\cpuregs[29][18] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\cpuregs[29][17] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\cpuregs[22][5] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\cpuregs[10][7] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\cpuregs[4][6] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(net142),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\cpuregs[20][26] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\cpuregs[13][20] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\cpuregs[23][25] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\cpuregs[16][7] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net45),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\cpuregs[6][29] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\cpuregs[21][17] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\cpuregs[15][26] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\cpuregs[4][13] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\cpuregs[20][11] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\cpuregs[2][18] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\cpuregs[8][3] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[22] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[11] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\cpuregs[10][13] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\cpuregs[29][16] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net161),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(net157),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\cpuregs[25][2] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\cpuregs[4][20] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\cpuregs[30][7] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\decoded_rd[0] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\cpuregs[8][17] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\cpuregs[14][24] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\cpuregs[24][29] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\cpuregs[21][12] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\cpuregs[20][13] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\cpuregs[24][1] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\cpuregs[27][10] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[31] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\cpuregs[22][10] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\cpuregs[31][5] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\cpuregs[29][31] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\cpuregs[16][16] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\cpuregs[13][5] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\cpuregs[24][15] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\cpuregs[13][10] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\cpuregs[4][16] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\cpuregs[16][21] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\cpuregs[31][14] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\cpuregs[12][21] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\cpuregs[8][11] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(net155),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\cpuregs[25][13] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\cpuregs[31][17] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\cpuregs[31][16] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\cpuregs[2][25] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\cpuregs[29][9] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\cpuregs[8][10] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\cpuregs[22][31] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\cpuregs[27][15] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\cpuregs[10][6] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\cpuregs[15][3] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\cpuregs[29][28] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\cpuregs[21][9] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\cpuregs[2][2] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\cpuregs[15][2] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\cpuregs[15][15] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\cpuregs[13][16] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\cpuregs[25][5] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\cpuregs[14][19] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\cpuregs[22][28] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\cpuregs[6][12] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(net173),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\cpuregs[2][19] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\cpuregs[28][16] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\cpuregs[30][1] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\cpuregs[28][30] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\cpuregs[15][28] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\cpuregs[24][27] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\cpuregs[16][18] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\cpuregs[28][10] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(net158),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\cpuregs[21][6] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\cpuregs[7][26] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\cpuregs[15][20] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\cpuregs[16][4] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\cpuregs[27][7] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\cpuregs[28][19] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\cpuregs[28][9] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\cpuregs[23][29] ),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\cpuregs[16][6] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\cpuregs[21][25] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\cpuregs[8][12] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\cpuregs[25][20] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\cpuregs[23][10] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\cpuregs[28][8] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\cpuregs[13][12] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(net153),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\cpuregs[2][16] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\cpuregs[26][19] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\cpuregs[22][18] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\cpuregs[25][18] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\cpuregs[30][17] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\cpuregs[25][15] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\cpuregs[10][23] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\cpuregs[10][17] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\cpuregs[16][12] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\cpuregs[16][15] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\cpuregs[23][27] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\cpuregs[2][8] ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\cpuregs[29][25] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\cpuregs[30][4] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\cpuregs[23][19] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\cpuregs[25][7] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\cpuregs[13][9] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\cpuregs[31][4] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\cpuregs[30][22] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(net44),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\cpuregs[4][2] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\cpuregs[29][29] ),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\cpuregs[23][2] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[8] ),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\cpuregs[12][26] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\cpuregs[10][12] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net65),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\cpuregs[21][18] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[30] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\cpuregs[25][21] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\cpuregs[8][29] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\cpuregs[15][17] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\cpuregs[21][11] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\cpuregs[29][14] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\cpuregs[6][26] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\cpuregs[25][14] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\cpuregs[16][1] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\cpuregs[22][3] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\cpuregs[6][6] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\cpuregs[28][7] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\cpuregs[3][6] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\cpuregs[26][11] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\cpuregs[20][14] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\cpuregs[29][8] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\cpuregs[20][16] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\cpuregs[27][3] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\cpuregs[27][5] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\cpuregs[15][22] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\cpuregs[15][5] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\cpuregs[13][14] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\cpuregs[27][8] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\cpuregs[27][9] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\cpuregs[13][22] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[7] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(instr_srai),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(net202),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\cpuregs[24][18] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\cpuregs[21][31] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\cpuregs[4][7] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\cpuregs[31][9] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\cpuregs[16][25] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\cpuregs[23][17] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\cpuregs[16][9] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\cpuregs[30][5] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\cpuregs[6][18] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\cpuregs[26][0] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\cpuregs[30][2] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\cpuregs[31][20] ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(net160),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_00973_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\cpuregs[16][22] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\cpuregs[4][12] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\cpuregs[23][11] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\cpuregs[6][4] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\cpuregs[21][22] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\cpuregs[13][13] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\cpuregs[6][2] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\cpuregs[15][16] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\cpuregs[25][16] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\cpuregs[21][13] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\cpuregs[27][20] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\cpuregs[21][3] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(net140),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\cpuregs[4][19] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\cpuregs[22][13] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\cpuregs[10][11] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\cpuregs[24][0] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\cpuregs[10][8] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(net184),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\cpuregs[29][7] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\cpuregs[25][3] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\cpuregs[25][11] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\cpuregs[2][0] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\cpuregs[8][24] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\cpuregs[10][25] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\cpuregs[28][31] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\cpuregs[16][19] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\cpuregs[8][1] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\cpuregs[27][21] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\cpuregs[7][3] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\cpuregs[31][28] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\cpuregs[27][18] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\cpuregs[5][0] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\cpuregs[5][8] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\cpuregs[21][16] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\cpuregs[5][18] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\cpuregs[6][11] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\cpuregs[13][1] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\cpuregs[29][4] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\cpuregs[10][30] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\cpuregs[21][4] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\cpuregs[4][21] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\cpuregs[25][10] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\cpuregs[2][9] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\cpuregs[5][7] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\cpuregs[6][28] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(net201),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\cpuregs[27][24] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\cpuregs[7][11] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\cpuregs[8][4] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\cpuregs[25][8] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\cpuregs[14][5] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\cpuregs[20][9] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\cpuregs[24][23] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\cpuregs[29][26] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\cpuregs[21][14] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\cpuregs[31][30] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\cpuregs[31][25] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\cpuregs[13][29] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\cpuregs[27][0] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\cpuregs[6][0] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\cpuregs[4][25] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\count_instr[63] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\cpuregs[25][4] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\cpuregs[4][5] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\cpuregs[15][8] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\cpuregs[3][15] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\cpuregs[2][26] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\cpuregs[12][12] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\cpuregs[15][24] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\cpuregs[23][7] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\cpuregs[2][28] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\cpuregs[20][1] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\cpuregs[3][18] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\cpuregs[15][19] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\cpuregs[10][2] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\cpuregs[4][15] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\cpuregs[28][17] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\cpuregs[7][25] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\cpuregs[8][7] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\cpuregs[22][7] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\cpuregs[21][27] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\cpuregs[7][13] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[61] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_01431_),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\cpuregs[25][27] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\cpuregs[8][6] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(net138),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\cpuregs[4][28] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\cpuregs[7][4] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\cpuregs[27][27] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\cpuregs[8][23] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\cpuregs[23][24] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\cpuregs[6][17] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\cpuregs[6][15] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(net178),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\cpuregs[8][0] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\cpuregs[15][12] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\cpuregs[2][13] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\cpuregs[4][17] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\cpuregs[27][13] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\cpuregs[6][27] ),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\cpuregs[15][18] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\cpuregs[13][30] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\cpuregs[27][6] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\cpuregs[16][11] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\cpuregs[9][11] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\cpuregs[10][26] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\cpuregs[4][23] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\cpuregs[2][22] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\cpuregs[27][17] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\cpuregs[25][28] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\cpuregs[4][0] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\cpuregs[27][16] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\cpuregs[21][29] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\cpuregs[29][23] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\cpuregs[14][12] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\cpuregs[20][31] ),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\cpuregs[6][13] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\cpuregs[29][24] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(instr_beq),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\cpuregs[4][30] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\cpuregs[4][14] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net47),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\cpuregs[22][30] ),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\cpuregs[10][20] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\cpuregs[25][17] ),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\cpuregs[7][10] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\cpuregs[7][12] ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\cpuregs[29][2] ),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\cpuregs[10][3] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\cpuregs[8][16] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\cpuregs[4][31] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\cpuregs[27][26] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\cpuregs[23][8] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\cpuregs[15][25] ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\cpuregs[2][20] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\cpuregs[4][9] ),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\cpuregs[6][22] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\cpuregs[25][23] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\cpuregs[25][24] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\cpuregs[16][10] ),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\cpuregs[31][22] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\cpuregs[2][10] ),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\cpuregs[15][31] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\cpuregs[5][10] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\cpuregs[3][13] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\cpuregs[10][19] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\cpuregs[6][9] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\cpuregs[5][23] ),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\cpuregs[3][20] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\cpuregs[27][12] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\cpuregs[5][12] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\cpuregs[5][17] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\cpuregs[4][4] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\cpuregs[27][11] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\cpuregs[7][20] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\cpuregs[3][26] ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\cpuregs[3][4] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\cpuregs[2][15] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\cpuregs[7][6] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\cpuregs[4][27] ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\cpuregs[27][28] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\cpuregs[8][22] ),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(net172),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\cpuregs[4][10] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\cpuregs[16][20] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\cpuregs[16][30] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\cpuregs[4][3] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\cpuregs[21][2] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\cpuregs[13][31] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\cpuregs[19][10] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\cpuregs[2][3] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\cpuregs[2][27] ),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\cpuregs[27][22] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(net186),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\cpuregs[2][30] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(net200),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\cpuregs[8][15] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\cpuregs[19][21] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\cpuregs[6][24] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\cpuregs[13][0] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\cpuregs[10][16] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\cpuregs[31][31] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\cpuregs[10][22] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\cpuregs[4][1] ),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\cpuregs[6][5] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\cpuregs[3][21] ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\cpuregs[27][23] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\cpuregs[8][5] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\cpuregs[6][20] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\cpuregs[6][21] ),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\cpuregs[16][13] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\cpuregs[31][0] ),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\cpuregs[16][24] ),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\cpuregs[31][19] ),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\cpuregs[6][1] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\cpuregs[16][5] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\cpuregs[8][30] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\cpuregs[23][31] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\cpuregs[8][26] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\cpuregs[27][1] ),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\cpuregs[14][11] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\cpuregs[8][9] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\cpuregs[23][26] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\cpuregs[6][8] ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\cpuregs[8][31] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\cpuregs[25][22] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\cpuregs[6][25] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\cpuregs[23][5] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\cpuregs[16][27] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[19] ),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\cpuregs[8][27] ),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[17] ),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\cpuregs[25][6] ),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\cpuregs[31][26] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\cpuregs[21][23] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\cpuregs[1][24] ),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\cpuregs[27][30] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\cpuregs[11][11] ),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\cpuregs[31][27] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\cpuregs[7][2] ),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\cpuregs[15][27] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(net181),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\cpuregs[7][8] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\cpuregs[20][19] ),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\cpuregs[19][29] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[21] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_01391_),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[44] ),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_01414_),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(net179),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\cpuregs[19][8] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\cpuregs[16][23] ),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\cpuregs[2][21] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\cpuregs[15][1] ),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\cpuregs[3][3] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\cpuregs[25][9] ),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\cpuregs[13][7] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\cpuregs[7][9] ),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\cpuregs[27][31] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\cpuregs[6][31] ),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\cpuregs[8][20] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\cpuregs[11][10] ),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\cpuregs[26][22] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\cpuregs[4][11] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\cpuregs[31][29] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\cpuregs[2][29] ),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\cpuregs[11][14] ),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\cpuregs[30][16] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\cpuregs[6][30] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\cpuregs[20][6] ),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\cpuregs[10][28] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\cpuregs[18][17] ),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\mem_wordsize[0] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[12] ),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\cpuregs[9][10] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\cpuregs[4][8] ),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\cpuregs[25][26] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\cpuregs[1][20] ),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\cpuregs[11][13] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\cpuregs[7][15] ),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\cpuregs[2][11] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\cpuregs[5][16] ),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\cpuregs[3][10] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\cpuregs[1][8] ),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\cpuregs[17][12] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\cpuregs[25][29] ),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\cpuregs[18][21] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\cpuregs[19][18] ),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\cpuregs[6][10] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\cpuregs[27][19] ),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\cpuregs[25][0] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\cpuregs[2][17] ),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\cpuregs[9][15] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\cpuregs[7][18] ),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\cpuregs[13][25] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\cpuregs[3][16] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\cpuregs[18][10] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\cpuregs[19][11] ),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\cpuregs[13][27] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\cpuregs[5][13] ),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\cpuregs[10][4] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\cpuregs[10][0] ),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\cpuregs[9][14] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\cpuregs[27][29] ),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\cpuregs[3][23] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\cpuregs[15][9] ),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\cpuregs[4][22] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\cpuregs[1][25] ),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\cpuregs[17][29] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\cpuregs[5][29] ),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\reg_sh[1] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\cpuregs[17][15] ),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\cpuregs[3][25] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\genblk2.pcpi_div.divisor[31] ),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_01136_),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\cpuregs[10][31] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\cpuregs[19][15] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\cpuregs[23][22] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\cpuregs[3][17] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\cpuregs[5][25] ),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\cpuregs[17][13] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\cpuregs[5][11] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\cpuregs[18][9] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\cpuregs[11][4] ),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\cpuregs[3][2] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\cpuregs[3][9] ),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\cpuregs[16][31] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\cpuregs[2][12] ),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\cpuregs[15][6] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\cpuregs[6][16] ),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\cpuregs[29][19] ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\cpuregs[23][0] ),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\cpuregs[17][10] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\cpuregs[27][4] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\cpuregs[9][20] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\cpuregs[8][25] ),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\cpuregs[3][14] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[16] ),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\cpuregs[9][13] ),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\cpuregs[29][1] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\cpuregs[6][14] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\cpuregs[23][20] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\cpuregs[3][8] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\cpuregs[19][2] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\cpuregs[18][15] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\cpuregs[10][5] ),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\cpuregs[18][2] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\cpuregs[11][9] ),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\cpuregs[2][6] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\cpuregs[3][24] ),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\cpuregs[18][13] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\cpuregs[5][5] ),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\cpuregs[17][2] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\cpuregs[11][16] ),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\cpuregs[17][16] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\cpuregs[5][20] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\cpuregs[18][0] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\cpuregs[18][26] ),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\cpuregs[4][18] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\cpuregs[21][26] ),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\cpuregs[9][4] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\cpuregs[1][7] ),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\cpuregs[18][22] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\cpuregs[5][15] ),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\cpuregs[2][5] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\cpuregs[31][1] ),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\cpuregs[25][19] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\cpuregs[3][27] ),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\cpuregs[17][17] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\cpuregs[1][16] ),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\cpuregs[17][23] ),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\cpuregs[3][12] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\cpuregs[17][8] ),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[47] ),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_01417_),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\cpuregs[9][17] ),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[55] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(_01425_),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(net177),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\cpuregs[11][12] ),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\cpuregs[19][9] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\cpuregs[2][23] ),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\cpuregs[6][7] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\cpuregs[9][5] ),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\cpuregs[21][30] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\cpuregs[19][13] ),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\cpuregs[13][28] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\cpuregs[18][25] ),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\cpuregs[11][7] ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\cpuregs[7][7] ),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\cpuregs[21][0] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\cpuregs[17][26] ),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\cpuregs[19][26] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\cpuregs[7][30] ),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\cpuregs[1][4] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\cpuregs[15][0] ),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\reg_next_pc[8] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\cpuregs[6][23] ),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(net57),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\cpuregs[11][21] ),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\cpuregs[19][20] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\cpuregs[3][7] ),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\cpuregs[25][1] ),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\cpuregs[25][30] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[50] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(_01420_),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\cpuregs[1][10] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\cpuregs[1][17] ),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\cpuregs[5][4] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\cpuregs[9][12] ),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\cpuregs[11][15] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\cpuregs[24][19] ),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\cpuregs[17][25] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\cpuregs[9][28] ),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\cpuregs[19][3] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\cpuregs[8][19] ),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\cpuregs[11][20] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\cpuregs[10][1] ),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\cpuregs[7][19] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\cpuregs[18][6] ),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\cpuregs[9][1] ),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(instr_addi),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\cpuregs[17][9] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\cpuregs[5][3] ),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\cpuregs[9][19] ),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\cpuregs[2][31] ),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[56] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\cpuregs[19][25] ),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\cpuregs[17][3] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[40] ),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_01410_),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\cpuregs[21][19] ),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\cpuregs[19][4] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[24] ),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\cpuregs[11][27] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\cpuregs[19][30] ),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\reg_next_pc[20] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\cpuregs[1][6] ),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\cpuregs[1][12] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\cpuregs[9][7] ),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[21] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\cpuregs[17][11] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\cpuregs[11][24] ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\cpuregs[13][26] ),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\cpuregs[5][6] ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\cpuregs[18][30] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\cpuregs[19][16] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\cpuregs[6][19] ),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\cpuregs[19][0] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\cpuregs[18][7] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\cpuregs[11][5] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\cpuregs[6][3] ),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\cpuregs[1][11] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\cpuregs[9][29] ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\cpuregs[7][29] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\cpuregs[18][16] ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\cpuregs[3][5] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\cpuregs[9][9] ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\cpuregs[10][24] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\cpuregs[5][2] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\cpuregs[2][1] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\cpuregs[16][28] ),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\cpuregs[23][1] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\cpuregs[7][5] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\cpuregs[12][24] ),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\cpuregs[17][18] ),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\cpuregs[1][0] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\cpuregs[1][1] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\cpuregs[9][0] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\cpuregs[1][22] ),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\cpuregs[9][25] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\cpuregs[18][24] ),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\cpuregs[25][25] ),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\cpuregs[9][3] ),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\cpuregs[9][27] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\cpuregs[10][27] ),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\cpuregs[7][21] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[32] ),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_01402_),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\cpuregs[19][12] ),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\cpuregs[7][0] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\cpuregs[2][4] ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\cpuregs[9][30] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\cpuregs[11][22] ),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\cpuregs[9][2] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\cpuregs[19][7] ),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\cpuregs[1][21] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\cpuregs[7][14] ),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\cpuregs[1][29] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(net183),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\cpuregs[5][1] ),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\cpuregs[1][13] ),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\cpuregs[5][31] ),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\cpuregs[5][27] ),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\cpuregs[11][17] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\cpuregs[23][28] ),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\cpuregs[5][21] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\cpuregs[19][19] ),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\cpuregs[17][14] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\cpuregs[17][24] ),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\cpuregs[11][23] ),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\cpuregs[25][31] ),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(instr_slli),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\cpuregs[4][24] ),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[17] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\cpuregs[7][16] ),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\cpuregs[18][8] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[58] ),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_01428_),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\cpuregs[13][24] ),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\cpuregs[18][12] ),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\cpuregs[9][22] ),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\cpuregs[17][27] ),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\cpuregs[21][28] ),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\cpuregs[17][21] ),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[53] ),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_01423_),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\cpuregs[9][24] ),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\cpuregs[11][31] ),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\cpuregs[18][18] ),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\cpuregs[19][14] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\cpuregs[5][24] ),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\cpuregs[5][22] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\cpuregs[19][28] ),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\cpuregs[7][24] ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\cpuregs[2][14] ),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\cpuregs[10][29] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\cpuregs[2][7] ),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\cpuregs[18][14] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\cpuregs[12][28] ),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\cpuregs[19][6] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\cpuregs[9][21] ),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[23] ),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[51] ),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\cpuregs[9][6] ),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\cpuregs[19][24] ),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\cpuregs[17][7] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\cpuregs[5][26] ),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(instr_fence),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\cpuregs[11][29] ),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(instr_add),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\cpuregs[5][14] ),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\cpuregs[5][9] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\cpuregs[1][15] ),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\cpuregs[7][31] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\cpuregs[11][3] ),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\cpuregs[18][23] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\cpuregs[17][22] ),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\cpuregs[11][8] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[1] ),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_01371_),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\cpuregs[1][19] ),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(\cpuregs[17][20] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\cpuregs[1][28] ),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\cpuregs[3][22] ),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\cpuregs[3][1] ),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\cpuregs[17][1] ),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\cpuregs[17][5] ),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\cpuregs[1][27] ),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\cpuregs[1][31] ),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\reg_next_pc[18] ),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[13] ),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\cpuregs[1][23] ),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(net185),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\cpuregs[11][19] ),
    .X(net2424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\cpuregs[5][19] ),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\cpuregs[1][18] ),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\cpuregs[3][19] ),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\cpuregs[13][19] ),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\cpuregs[19][22] ),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[13] ),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\cpuregs[17][31] ),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[37] ),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(_01407_),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\cpuregs[3][11] ),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[10] ),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\cpuregs[17][4] ),
    .X(net2436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\cpuregs[7][22] ),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\cpuregs[7][27] ),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\cpuregs[17][6] ),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\cpuregs[18][4] ),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\cpuregs[17][30] ),
    .X(net2441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\cpuregs[27][25] ),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[54] ),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\cpuregs[7][1] ),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\cpuregs[1][14] ),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\reg_next_pc[11] ),
    .X(net2446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\cpuregs[9][8] ),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(\cpuregs[19][5] ),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\cpuregs[7][17] ),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\cpuregs[18][19] ),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\cpuregs[11][6] ),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\cpuregs[18][11] ),
    .X(net2452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\cpuregs[3][29] ),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\cpuregs[19][23] ),
    .X(net2454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\genblk2.pcpi_div.divisor[62] ),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(\cpuregs[3][30] ),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\cpuregs[1][26] ),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\cpuregs[18][27] ),
    .X(net2458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\cpuregs[16][0] ),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\cpuregs[19][1] ),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\cpuregs[11][2] ),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\cpuregs[9][18] ),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\cpuregs[7][28] ),
    .X(net2463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\cpuregs[11][18] ),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\cpuregs[9][23] ),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\cpuregs[19][31] ),
    .X(net2466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(net49),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\cpuregs[5][30] ),
    .X(net2468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[49] ),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_01419_),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\cpuregs[7][23] ),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[36] ),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(_01406_),
    .X(net2473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\cpuregs[18][3] ),
    .X(net2474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\cpuregs[18][20] ),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[59] ),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[31] ),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[35] ),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(_01405_),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[39] ),
    .X(net2480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(_01409_),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(\cpuregs[1][5] ),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[18] ),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(\cpuregs[17][28] ),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\cpuregs[1][3] ),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(\cpuregs[11][30] ),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\reg_next_pc[23] ),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(\cpuregs[9][16] ),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[48] ),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\cpuregs[9][31] ),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[57] ),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\cpuregs[19][27] ),
    .X(net2492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\cpuregs[18][29] ),
    .X(net2493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\cpuregs[17][19] ),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\cpuregs[3][28] ),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(\cpuregs[11][25] ),
    .X(net2496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\cpuregs[11][0] ),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(net54),
    .X(net2498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\cpuregs[23][30] ),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(\cpuregs[11][26] ),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[34] ),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_01404_),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\cpuregs[5][28] ),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[43] ),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(_01413_),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(\cpuregs[18][31] ),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\cpuregs[11][1] ),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[60] ),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\cpuregs[11][28] ),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\cpuregs[9][26] ),
    .X(net2510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[20] ),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(\reg_next_pc[31] ),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\cpuregs[1][9] ),
    .X(net2513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(\cpuregs[1][30] ),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\genblk1.genblk1.pcpi_mul.mul_counter[6] ),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_00195_),
    .X(net2516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[46] ),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_01416_),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[52] ),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[8] ),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[33] ),
    .X(net2521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\cpuregs[19][17] ),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\cpuregs[18][1] ),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\cpuregs[1][2] ),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\cpuregs[3][31] ),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\cpuregs[17][0] ),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\genblk1.genblk1.pcpi_mul.rs2[63] ),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_01369_),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\genblk2.pcpi_div.quotient_msk[5] ),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_01046_),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\cpuregs[18][28] ),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\cpuregs[3][0] ),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\genblk2.pcpi_div.divisor[41] ),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\genblk2.pcpi_div.divisor[53] ),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\genblk2.pcpi_div.divisor[57] ),
    .X(net2535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\genblk2.pcpi_div.divisor[44] ),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\cpuregs[18][5] ),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\cpuregs[21][1] ),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[5] ),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[41] ),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[45] ),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\pcpi_timeout_counter[3] ),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\genblk2.pcpi_div.divisor[47] ),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[3] ),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\genblk2.pcpi_div.divisor[35] ),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(\genblk2.pcpi_div.divisor[37] ),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\cpuregs[30][26] ),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(net151),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[12] ),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(instr_sltiu),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\genblk2.pcpi_div.divisor[36] ),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\genblk2.pcpi_div.divisor[33] ),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\genblk2.pcpi_div.divisor[58] ),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(net171),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(_00822_),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(net216),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(instr_lui),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\count_instr[1] ),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\genblk1.genblk1.pcpi_mul.rd[20] ),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\reg_next_pc[7] ),
    .X(net2560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\count_instr[17] ),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_00600_),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\genblk2.pcpi_div.divisor[48] ),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\reg_next_pc[22] ),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\reg_next_pc[21] ),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\genblk2.pcpi_div.divisor[39] ),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\genblk1.genblk1.pcpi_mul.rd[16] ),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[15] ),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\reg_next_pc[16] ),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\genblk2.pcpi_div.divisor[34] ),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\genblk2.pcpi_div.divisor[38] ),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(instr_sltu),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[42] ),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(\genblk1.genblk1.pcpi_mul.rd[12] ),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[28] ),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(\genblk1.genblk1.pcpi_mul.rd[48] ),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\genblk1.genblk1.pcpi_mul.rd[28] ),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(\reg_next_pc[19] ),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\genblk2.pcpi_div.divisor[0] ),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_01106_),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\genblk2.pcpi_div.divisor[54] ),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\count_instr[34] ),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(_00617_),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\count_instr[49] ),
    .X(net2584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(_00632_),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(\reg_next_pc[29] ),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\genblk1.genblk1.pcpi_mul.rd[24] ),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(net195),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\genblk2.pcpi_div.divisor[61] ),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\count_instr[53] ),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(_00636_),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\genblk1.genblk1.pcpi_mul.rd[8] ),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\reg_next_pc[6] ),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[38] ),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\genblk2.pcpi_div.quotient[26] ),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_06605_),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\reg_next_pc[27] ),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\genblk1.genblk1.pcpi_mul.rd[40] ),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\genblk2.pcpi_div.divisor[40] ),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\genblk2.pcpi_div.divisor[50] ),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[14] ),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\genblk2.pcpi_div.quotient_msk[0] ),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(_01042_),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\genblk1.genblk1.pcpi_mul.rd[4] ),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\count_cycle[0] ),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\pcpi_timeout_counter[2] ),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\reg_next_pc[30] ),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(instr_sra),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(instr_blt),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\genblk1.genblk1.pcpi_mul.rd[52] ),
    .X(net2610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(net180),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(net196),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(_00825_),
    .X(net2613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\genblk1.genblk1.pcpi_mul.rd[1] ),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\count_instr[23] ),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_00606_),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\reg_next_pc[15] ),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\genblk2.pcpi_div.quotient[31] ),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(_06610_),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\cpuregs[16][29] ),
    .X(net2620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\genblk1.genblk1.pcpi_mul.rdx[20] ),
    .X(net2621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\genblk1.genblk1.pcpi_mul.rd[32] ),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\genblk2.pcpi_div.divisor[45] ),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\genblk1.genblk1.pcpi_mul.rd[2] ),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\genblk1.genblk1.pcpi_mul.rdx[28] ),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\genblk1.genblk1.pcpi_mul.rd[14] ),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\genblk2.pcpi_div.divisor[59] ),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\genblk1.genblk1.pcpi_mul.rd[10] ),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[11] ),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\reg_next_pc[2] ),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\genblk2.pcpi_div.divisor[56] ),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\genblk1.genblk1.pcpi_mul.rd[18] ),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[17] ),
    .X(net2633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\genblk2.pcpi_div.divisor[60] ),
    .X(net2634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[4] ),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(net197),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(_00826_),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\reg_next_pc[9] ),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\reg_next_pc[28] ),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\genblk1.genblk1.pcpi_mul.rdx[48] ),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\genblk1.genblk1.pcpi_mul.rd[56] ),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\reg_next_pc[14] ),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(net192),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\reg_next_pc[26] ),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\mem_rdata_q[1] ),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\genblk1.genblk1.pcpi_mul.rdx[8] ),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(net143),
    .X(net2647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(net182),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\genblk1.genblk1.pcpi_mul.rdx[12] ),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\genblk1.genblk1.pcpi_mul.rd[36] ),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\reg_next_pc[3] ),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\genblk1.genblk1.pcpi_mul.rd[50] ),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\genblk2.pcpi_div.divisor[51] ),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(instr_slt),
    .X(net2654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(_00002_),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[20] ),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\genblk2.pcpi_div.divisor[15] ),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\genblk1.genblk1.pcpi_mul.rd[6] ),
    .X(net2659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\genblk1.genblk1.pcpi_mul.rd[22] ),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\genblk2.pcpi_div.divisor[9] ),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\genblk1.genblk1.pcpi_mul.rdx[36] ),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\genblk2.pcpi_div.running ),
    .X(net2663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\genblk2.pcpi_div.divisor[49] ),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\genblk1.genblk1.pcpi_mul.rdx[60] ),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\genblk2.pcpi_div.divisor[46] ),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\reg_next_pc[17] ),
    .X(net2667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[8] ),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\genblk2.pcpi_div.divisor[43] ),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\genblk1.genblk1.pcpi_mul.rdx[56] ),
    .X(net2670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(is_slli_srli_srai),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(_00924_),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\cpu_state[0] ),
    .X(net2673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\genblk1.genblk1.pcpi_mul.rdx[4] ),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\reg_next_pc[12] ),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(\genblk1.genblk1.pcpi_mul.rd[44] ),
    .X(net2676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\genblk2.pcpi_div.divisor[13] ),
    .X(net2677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_01118_),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\genblk1.genblk1.pcpi_mul.rdx[44] ),
    .X(net2679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(net188),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\genblk1.genblk1.pcpi_mul.rd[0] ),
    .X(net2681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(\genblk1.genblk1.pcpi_mul.rd[42] ),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\genblk1.genblk1.pcpi_mul.rd[26] ),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(net189),
    .X(net2684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\genblk2.pcpi_div.quotient[6] ),
    .X(net2685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_06585_),
    .X(net2686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\genblk2.pcpi_div.divisor[42] ),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(is_sll_srl_sra),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\reg_next_pc[10] ),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(\genblk2.pcpi_div.divisor[52] ),
    .X(net2690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\genblk1.genblk1.pcpi_mul.rd[38] ),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\genblk2.pcpi_div.divisor[24] ),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(_01129_),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\genblk2.pcpi_div.quotient[3] ),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(_06582_),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\genblk1.genblk1.pcpi_mul.rd[30] ),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\genblk1.genblk1.pcpi_mul.rd[46] ),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(net154),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\mem_rdata_q[0] ),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[2] ),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\count_cycle[48] ),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\genblk2.pcpi_div.divisor[17] ),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\genblk1.genblk1.pcpi_mul.rd[34] ),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\genblk2.pcpi_div.divisor[12] ),
    .X(net2704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(_01117_),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\genblk1.genblk1.pcpi_mul.rdx[24] ),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\genblk1.genblk1.pcpi_mul.rd[58] ),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\genblk1.genblk1.pcpi_mul.rdx[52] ),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\genblk1.genblk1.pcpi_mul.mul_counter[2] ),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(is_alu_reg_reg),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\genblk1.genblk1.pcpi_mul.rdx[40] ),
    .X(net2711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\genblk1.genblk1.pcpi_mul.rdx[16] ),
    .X(net2712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\genblk2.pcpi_div.quotient[11] ),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(_06590_),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\genblk2.pcpi_div.divisor[7] ),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(_01112_),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\genblk2.pcpi_div.divisor[4] ),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_01109_),
    .X(net2718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\genblk2.pcpi_div.divisor[16] ),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\count_cycle[15] ),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\genblk1.genblk1.pcpi_mul.rd[61] ),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\genblk2.pcpi_div.divisor[55] ),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[9] ),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[25] ),
    .X(net2724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\genblk2.pcpi_div.quotient[24] ),
    .X(net2725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_06603_),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(instr_or),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(\genblk2.pcpi_div.divisor[14] ),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(net191),
    .X(net2729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[28] ),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\genblk2.pcpi_div.divisor[21] ),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\genblk2.pcpi_div.quotient_msk[29] ),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(_01070_),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\genblk2.pcpi_div.divisor[5] ),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\genblk2.pcpi_div.quotient[17] ),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(_06596_),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(net199),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(_00828_),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[11] ),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\reg_next_pc[4] ),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\reg_next_pc[13] ),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\genblk2.pcpi_div.divisor[10] ),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\genblk2.pcpi_div.divisor[27] ),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_01132_),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\count_cycle[37] ),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\genblk2.pcpi_div.quotient[0] ),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\count_cycle[28] ),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(\genblk1.genblk1.pcpi_mul.rd[21] ),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\genblk1.genblk1.pcpi_mul.rd[9] ),
    .X(net2749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(\genblk2.pcpi_div.quotient_msk[2] ),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(_01043_),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[19] ),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\genblk2.pcpi_div.quotient[30] ),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(_06609_),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\genblk1.genblk1.pcpi_mul.rd[54] ),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\genblk2.pcpi_div.quotient_msk[9] ),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(_01050_),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\count_cycle[56] ),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[1] ),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\mem_state[0] ),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\genblk2.pcpi_div.quotient[20] ),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_06599_),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[20] ),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(net218),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\genblk1.genblk1.pcpi_mul.rd[13] ),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(\genblk2.pcpi_div.quotient[23] ),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(_06602_),
    .X(net2767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(\reg_sh[2] ),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\genblk2.pcpi_div.divisor[18] ),
    .X(net2769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(_01123_),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\genblk2.pcpi_div.divisor[32] ),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[0] ),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\genblk1.genblk1.pcpi_mul.rd[5] ),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(\count_instr[18] ),
    .X(net2774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\genblk2.pcpi_div.divisor[25] ),
    .X(net2775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\genblk2.pcpi_div.quotient_msk[16] ),
    .X(net2776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(_01057_),
    .X(net2777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(instr_bge),
    .X(net2778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\count_instr[14] ),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(\genblk1.genblk1.pcpi_mul.rdx[32] ),
    .X(net2780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\genblk1.genblk1.pcpi_mul.rd[25] ),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(\genblk2.pcpi_div.divisor[26] ),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(\count_cycle[50] ),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(\count_cycle[12] ),
    .X(net2784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\genblk2.pcpi_div.quotient_msk[15] ),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(_01056_),
    .X(net2786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\count_cycle[17] ),
    .X(net2787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(\count_cycle[31] ),
    .X(net2788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\genblk1.genblk1.pcpi_mul.rd[29] ),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(\count_cycle[9] ),
    .X(net2790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\genblk2.pcpi_div.quotient_msk[25] ),
    .X(net2791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(_01066_),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\mem_rdata_q[3] ),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\genblk2.pcpi_div.quotient_msk[20] ),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(_01061_),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\count_instr[39] ),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\count_cycle[60] ),
    .X(net2797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\genblk2.pcpi_div.quotient_msk[10] ),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\count_instr[36] ),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(instr_sll),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\genblk2.pcpi_div.quotient[10] ),
    .X(net2801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(instr_slti),
    .X(net2802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\genblk2.pcpi_div.quotient_msk[12] ),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_01053_),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\count_instr[31] ),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\genblk2.pcpi_div.quotient[28] ),
    .X(net2806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(_06607_),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\genblk2.pcpi_div.quotient[22] ),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(_06601_),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\genblk2.pcpi_div.quotient_msk[21] ),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\genblk1.genblk1.pcpi_mul.mul_counter[4] ),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\genblk2.pcpi_div.quotient[19] ),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(_06598_),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[15] ),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\genblk1.genblk1.pcpi_mul.rd[60] ),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\genblk2.pcpi_div.divisor[22] ),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(net134),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\genblk2.pcpi_div.divisor[19] ),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\genblk2.pcpi_div.quotient[16] ),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\genblk2.pcpi_div.quotient[25] ),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(\reg_next_pc[5] ),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[16] ),
    .X(net2822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[21] ),
    .X(net2823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(\count_cycle[46] ),
    .X(net2824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\count_instr[21] ),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[44] ),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(_01350_),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\genblk2.pcpi_div.quotient_msk[22] ),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\genblk2.pcpi_div.quotient[15] ),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[12] ),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\count_instr[8] ),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\count_instr[45] ),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\genblk2.pcpi_div.quotient_msk[6] ),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\genblk2.pcpi_div.quotient[13] ),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(_06592_),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\count_instr[42] ),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\genblk1.genblk1.pcpi_mul.pcpi_rd[6] ),
    .X(net2837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\genblk1.genblk1.pcpi_mul.rd[17] ),
    .X(net2838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\genblk2.pcpi_div.quotient_msk[19] ),
    .X(net2839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(_01060_),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\count_cycle[40] ),
    .X(net2841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\genblk1.genblk1.pcpi_mul.rd[41] ),
    .X(net2842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\genblk2.pcpi_div.quotient_msk[28] ),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(_01069_),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[51] ),
    .X(net2845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(_01357_),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\genblk2.pcpi_div.quotient_msk[30] ),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(\count_cycle[6] ),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(instr_lhu),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(\pcpi_timeout_counter[0] ),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\count_cycle[22] ),
    .X(net2851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(instr_jalr),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(\genblk2.pcpi_div.divisor[11] ),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\genblk2.pcpi_div.quotient[27] ),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(\count_instr[59] ),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(\genblk2.pcpi_div.quotient_msk[17] ),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\count_cycle[3] ),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(\genblk2.pcpi_div.quotient_msk[3] ),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\genblk2.pcpi_div.quotient_msk[13] ),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(\count_cycle[43] ),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\pcpi_timeout_counter[1] ),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(\count_cycle[53] ),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(\genblk2.pcpi_div.quotient_msk[14] ),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(instr_ori),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\count_instr[62] ),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(\genblk2.pcpi_div.quotient_msk[11] ),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\genblk2.pcpi_div.quotient_msk[24] ),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_01065_),
    .X(net2868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\genblk1.genblk1.pcpi_mul.rd[37] ),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(\genblk1.genblk1.pcpi_mul.rd[49] ),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\genblk1.genblk1.pcpi_mul.rd[45] ),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\genblk1.genblk1.pcpi_mul.rd[3] ),
    .X(net2872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\genblk2.pcpi_div.divisor[29] ),
    .X(net2873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_01134_),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(net190),
    .X(net2875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\genblk2.pcpi_div.divisor[23] ),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\genblk2.pcpi_div.quotient[9] ),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(\genblk1.genblk1.pcpi_mul.rd[57] ),
    .X(net2878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\genblk2.pcpi_div.quotient_msk[31] ),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(\genblk1.genblk1.pcpi_mul.rd[15] ),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\genblk2.pcpi_div.quotient[21] ),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(\genblk2.pcpi_div.quotient_msk[26] ),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\genblk1.genblk1.pcpi_mul.rd[7] ),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\genblk1.genblk1.pcpi_mul.rd[53] ),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\count_cycle[19] ),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(\genblk2.pcpi_div.quotient_msk[23] ),
    .X(net2886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\genblk2.pcpi_div.divisor[6] ),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(\genblk1.genblk1.pcpi_mul.rd[19] ),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\count_instr[56] ),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[16] ),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\genblk2.pcpi_div.divisor[30] ),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(\count_instr[28] ),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\genblk2.pcpi_div.quotient_msk[18] ),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[37] ),
    .X(net2894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(_01343_),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(instr_sw),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\genblk1.genblk1.pcpi_mul.rd[23] ),
    .X(net2897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\genblk2.pcpi_div.divisor[3] ),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(_01108_),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[57] ),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(_01363_),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[6] ),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\genblk2.pcpi_div.divisor[28] ),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(instr_lw),
    .X(net2904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[53] ),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(\count_cycle[1] ),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(_00710_),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\genblk2.pcpi_div.quotient[2] ),
    .X(net2908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\genblk2.pcpi_div.quotient_msk[7] ),
    .X(net2909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(\reg_next_pc[24] ),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\genblk1.genblk1.pcpi_mul.rd[11] ),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(instr_sb),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\genblk1.genblk1.pcpi_mul.rd[47] ),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[5] ),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[47] ),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(_01353_),
    .X(net2916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\genblk1.genblk1.pcpi_mul.rd[59] ),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(\genblk1.genblk1.pcpi_mul.rd[33] ),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\genblk1.genblk1.pcpi_mul.rd[31] ),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(\genblk2.pcpi_div.quotient_msk[8] ),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(\genblk1.genblk1.pcpi_mul.rd[27] ),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(instr_andi),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[22] ),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(\genblk1.genblk1.pcpi_mul.rd[39] ),
    .X(net2924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\genblk2.pcpi_div.quotient[5] ),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(\genblk2.pcpi_div.quotient[18] ),
    .X(net2926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\genblk1.genblk1.pcpi_mul.rd[55] ),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[49] ),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(_01355_),
    .X(net2929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(instr_lbu),
    .X(net2930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\genblk1.genblk1.pcpi_mul.rd[35] ),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(instr_sh),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\genblk2.pcpi_div.quotient[8] ),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_06587_),
    .X(net2934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\count_instr[25] ),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\mem_rdata_q[4] ),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\genblk2.pcpi_div.quotient[7] ),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[43] ),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[33] ),
    .X(net2939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\count_cycle[34] ),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(\genblk1.genblk1.pcpi_mul.rd[63] ),
    .X(net2941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[41] ),
    .X(net2942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(_01347_),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(\genblk2.pcpi_div.quotient[14] ),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[61] ),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_01367_),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\mem_rdata_q[6] ),
    .X(net2947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[48] ),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\genblk1.genblk1.pcpi_mul.rd[62] ),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[4] ),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(_01310_),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[56] ),
    .X(net2952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[36] ),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(\count_instr[51] ),
    .X(net2954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[55] ),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[62] ),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(_01368_),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[59] ),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(_01365_),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\mem_state[1] ),
    .X(net2960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\genblk2.pcpi_div.quotient[12] ),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_06591_),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[60] ),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\genblk2.pcpi_div.divisor[2] ),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(_01107_),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\genblk2.pcpi_div.quotient_msk[4] ),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\genblk1.genblk1.pcpi_mul.rd[43] ),
    .X(net2967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\count_cycle[59] ),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[58] ),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[18] ),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[24] ),
    .X(net2971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(\count_cycle[21] ),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\count_instr[7] ),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\count_instr[13] ),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[42] ),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\count_instr[27] ),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[52] ),
    .X(net2977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[46] ),
    .X(net2978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[35] ),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(net198),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(_00827_),
    .X(net2981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(\count_instr[3] ),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[7] ),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(\decoded_imm_j[8] ),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\genblk2.pcpi_div.quotient[29] ),
    .X(net2985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\genblk2.pcpi_div.quotient_msk[27] ),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\count_cycle[27] ),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(\count_cycle[16] ),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\genblk2.pcpi_div.dividend[31] ),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\genblk1.genblk1.pcpi_mul.mul_counter[0] ),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\count_cycle[62] ),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\count_instr[35] ),
    .X(net2992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[13] ),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(instr_bgeu),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\genblk1.genblk1.pcpi_mul.rd[51] ),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(\count_cycle[24] ),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\count_instr[20] ),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(\count_instr[24] ),
    .X(net2998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(\genblk2.pcpi_div.quotient[1] ),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(_06580_),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\count_cycle[52] ),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[23] ),
    .X(net3002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[29] ),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[10] ),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(instr_and),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[40] ),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[34] ),
    .X(net3007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(mem_do_rdata),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[27] ),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(\genblk2.pcpi_div.dividend[5] ),
    .X(net3010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\genblk2.pcpi_div.quotient[4] ),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(\genblk1.genblk1.pcpi_mul.mul_counter[1] ),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\count_instr[55] ),
    .X(net3013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[26] ),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\mem_rdata_q[5] ),
    .X(net3015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\reg_sh[0] ),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\reg_next_pc[25] ),
    .X(net3017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(instr_bne),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\decoded_imm[2] ),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(\genblk2.pcpi_div.dividend[13] ),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\genblk2.pcpi_div.dividend[18] ),
    .X(net3021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[3] ),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[31] ),
    .X(net3023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(instr_xori),
    .X(net3024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\genblk2.pcpi_div.dividend[12] ),
    .X(net3025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(latched_is_lh),
    .X(net3026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[30] ),
    .X(net3027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\count_instr[2] ),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(instr_rdinstr),
    .X(net3029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(\count_cycle[35] ),
    .X(net3030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\genblk2.pcpi_div.pcpi_wait ),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(instr_xor),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\genblk2.pcpi_div.dividend[28] ),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(\count_instr[54] ),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[38] ),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(instr_lb),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\reg_pc[19] ),
    .X(net3037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\count_cycle[23] ),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\count_cycle[4] ),
    .X(net3039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\count_instr[19] ),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\count_cycle[13] ),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\count_instr[15] ),
    .X(net3042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\genblk2.pcpi_div.dividend[14] ),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\decoded_imm_j[19] ),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\count_cycle[54] ),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[50] ),
    .X(net3046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\count_instr[29] ),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\mem_rdata_q[2] ),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(net176),
    .X(net3049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\genblk2.pcpi_div.dividend[23] ),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\count_instr[50] ),
    .X(net3051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(is_compare),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\count_instr[6] ),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\count_cycle[10] ),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(\decoded_imm[16] ),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\decoded_imm[19] ),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(instr_rdcycle),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(\genblk2.pcpi_div.dividend[4] ),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(\reg_pc[23] ),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(\count_instr[37] ),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(\reg_pc[16] ),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\count_cycle[32] ),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\decoded_imm[15] ),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(\decoded_imm_j[5] ),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\count_instr[12] ),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(\count_instr[26] ),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\count_cycle[41] ),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(\genblk1.genblk1.pcpi_mul.next_rs1[24] ),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\genblk2.pcpi_div.divisor[16] ),
    .X(net3069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[46] ),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\genblk1.genblk1.pcpi_mul.next_rs2[34] ),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\genblk2.pcpi_div.quotient_msk[27] ),
    .X(net3072));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02829_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_02832_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_02950_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_03097_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_03124_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_03743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_03747_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_03839_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_04256_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_04888_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_05637_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_05637_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_06718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\alu_out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\alu_out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\alu_out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\alu_out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\alu_out[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\cpu_state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\cpu_state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\cpu_state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\genblk2.pcpi_div.pcpi_rd[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\genblk2.pcpi_div.pcpi_rd[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\genblk2.pcpi_div.pcpi_rd[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\genblk2.pcpi_div.pcpi_rd[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\genblk2.pcpi_div.pcpi_rd[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\genblk2.pcpi_div.pcpi_rd[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\genblk2.pcpi_div.pcpi_rd[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\genblk2.pcpi_div.pcpi_rd[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\genblk2.pcpi_div.pcpi_rd[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\genblk2.pcpi_div.pcpi_rd[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\genblk2.pcpi_div.pcpi_rd[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\genblk2.pcpi_div.pcpi_rd[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\genblk2.pcpi_div.pcpi_rd[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\genblk2.pcpi_div.pcpi_rd[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\genblk2.pcpi_div.pcpi_rd[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\genblk2.pcpi_div.pcpi_rd[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\genblk2.pcpi_div.pcpi_rd[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\genblk2.pcpi_div.pcpi_rd[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\genblk2.pcpi_div.pcpi_rd[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\genblk2.pcpi_div.pcpi_rd[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\genblk2.pcpi_div.pcpi_rd[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\genblk2.pcpi_div.pcpi_rd[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\genblk2.pcpi_div.pcpi_rd[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\genblk2.pcpi_div.pcpi_rd[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\genblk2.pcpi_div.pcpi_rd[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\genblk2.pcpi_div.pcpi_rd[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\genblk2.pcpi_div.pcpi_rd[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\genblk2.pcpi_div.pcpi_rd[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\genblk2.pcpi_div.pcpi_rd[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\genblk2.pcpi_div.pcpi_rd[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\genblk2.pcpi_div.pcpi_rd[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\genblk2.pcpi_div.pcpi_rd[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\genblk2.pcpi_div.pcpi_rd[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\genblk2.pcpi_div.pcpi_rd[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\mem_rdata_q[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\mem_rdata_q[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_02756_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\alu_out_q[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\genblk2.pcpi_div.pcpi_rd[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\genblk2.pcpi_div.pcpi_rd[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\genblk2.pcpi_div.pcpi_rd[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\genblk2.pcpi_div.pcpi_rd[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\genblk2.pcpi_div.pcpi_rd[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\genblk2.pcpi_div.pcpi_rd[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(instr_rdcycleh));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\mem_rdata_q[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(\mem_rdata_q[16] ));
 sky130_ef_sc_hd__decap_12 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1009 ();
 assign eoi[0] = net1242;
 assign eoi[10] = net1252;
 assign eoi[11] = net1253;
 assign eoi[12] = net1254;
 assign eoi[13] = net1255;
 assign eoi[14] = net1256;
 assign eoi[15] = net1257;
 assign eoi[16] = net1258;
 assign eoi[17] = net1259;
 assign eoi[18] = net1260;
 assign eoi[19] = net1261;
 assign eoi[1] = net1243;
 assign eoi[20] = net1262;
 assign eoi[21] = net1263;
 assign eoi[22] = net1264;
 assign eoi[23] = net1265;
 assign eoi[24] = net1266;
 assign eoi[25] = net1267;
 assign eoi[26] = net1268;
 assign eoi[27] = net1269;
 assign eoi[28] = net1270;
 assign eoi[29] = net1271;
 assign eoi[2] = net1244;
 assign eoi[30] = net1272;
 assign eoi[31] = net1273;
 assign eoi[3] = net1245;
 assign eoi[4] = net1246;
 assign eoi[5] = net1247;
 assign eoi[6] = net1248;
 assign eoi[7] = net1249;
 assign eoi[8] = net1250;
 assign eoi[9] = net1251;
 assign mem_addr[0] = net1274;
 assign mem_addr[1] = net1275;
 assign mem_la_addr[0] = net1276;
 assign mem_la_addr[1] = net1277;
 assign trace_data[0] = net1278;
 assign trace_data[10] = net1288;
 assign trace_data[11] = net1289;
 assign trace_data[12] = net1290;
 assign trace_data[13] = net1291;
 assign trace_data[14] = net1292;
 assign trace_data[15] = net1293;
 assign trace_data[16] = net1294;
 assign trace_data[17] = net1295;
 assign trace_data[18] = net1296;
 assign trace_data[19] = net1297;
 assign trace_data[1] = net1279;
 assign trace_data[20] = net1298;
 assign trace_data[21] = net1299;
 assign trace_data[22] = net1300;
 assign trace_data[23] = net1301;
 assign trace_data[24] = net1302;
 assign trace_data[25] = net1303;
 assign trace_data[26] = net1304;
 assign trace_data[27] = net1305;
 assign trace_data[28] = net1306;
 assign trace_data[29] = net1307;
 assign trace_data[2] = net1280;
 assign trace_data[30] = net1308;
 assign trace_data[31] = net1309;
 assign trace_data[32] = net1310;
 assign trace_data[33] = net1311;
 assign trace_data[34] = net1312;
 assign trace_data[35] = net1313;
 assign trace_data[3] = net1281;
 assign trace_data[4] = net1282;
 assign trace_data[5] = net1283;
 assign trace_data[6] = net1284;
 assign trace_data[7] = net1285;
 assign trace_data[8] = net1286;
 assign trace_data[9] = net1287;
 assign trace_valid = net1314;
endmodule
